`timescale 1ns / 1ps
`default_nettype none


//Created by script createsinelookup.py
module sinetable(input wire [11:0] phase, output reg [9:0] result);

always @(*)
  case(phase)
   0: result <= 10'b0000000000;
   1: result <= 10'b0000000001;
   2: result <= 10'b0000000010;
   3: result <= 10'b0000000010;
   4: result <= 10'b0000000011;
   5: result <= 10'b0000000100;
   6: result <= 10'b0000000101;
   7: result <= 10'b0000000101;
   8: result <= 10'b0000000110;
   9: result <= 10'b0000000111;
   10: result <= 10'b0000001000;
   11: result <= 10'b0000001001;
   12: result <= 10'b0000001001;
   13: result <= 10'b0000001010;
   14: result <= 10'b0000001011;
   15: result <= 10'b0000001100;
   16: result <= 10'b0000001101;
   17: result <= 10'b0000001101;
   18: result <= 10'b0000001110;
   19: result <= 10'b0000001111;
   20: result <= 10'b0000010000;
   21: result <= 10'b0000010000;
   22: result <= 10'b0000010001;
   23: result <= 10'b0000010010;
   24: result <= 10'b0000010011;
   25: result <= 10'b0000010100;
   26: result <= 10'b0000010100;
   27: result <= 10'b0000010101;
   28: result <= 10'b0000010110;
   29: result <= 10'b0000010111;
   30: result <= 10'b0000011000;
   31: result <= 10'b0000011000;
   32: result <= 10'b0000011001;
   33: result <= 10'b0000011010;
   34: result <= 10'b0000011011;
   35: result <= 10'b0000011011;
   36: result <= 10'b0000011100;
   37: result <= 10'b0000011101;
   38: result <= 10'b0000011110;
   39: result <= 10'b0000011111;
   40: result <= 10'b0000011111;
   41: result <= 10'b0000100000;
   42: result <= 10'b0000100001;
   43: result <= 10'b0000100010;
   44: result <= 10'b0000100011;
   45: result <= 10'b0000100011;
   46: result <= 10'b0000100100;
   47: result <= 10'b0000100101;
   48: result <= 10'b0000100110;
   49: result <= 10'b0000100110;
   50: result <= 10'b0000100111;
   51: result <= 10'b0000101000;
   52: result <= 10'b0000101001;
   53: result <= 10'b0000101010;
   54: result <= 10'b0000101010;
   55: result <= 10'b0000101011;
   56: result <= 10'b0000101100;
   57: result <= 10'b0000101101;
   58: result <= 10'b0000101101;
   59: result <= 10'b0000101110;
   60: result <= 10'b0000101111;
   61: result <= 10'b0000110000;
   62: result <= 10'b0000110001;
   63: result <= 10'b0000110001;
   64: result <= 10'b0000110010;
   65: result <= 10'b0000110011;
   66: result <= 10'b0000110100;
   67: result <= 10'b0000110101;
   68: result <= 10'b0000110101;
   69: result <= 10'b0000110110;
   70: result <= 10'b0000110111;
   71: result <= 10'b0000111000;
   72: result <= 10'b0000111000;
   73: result <= 10'b0000111001;
   74: result <= 10'b0000111010;
   75: result <= 10'b0000111011;
   76: result <= 10'b0000111100;
   77: result <= 10'b0000111100;
   78: result <= 10'b0000111101;
   79: result <= 10'b0000111110;
   80: result <= 10'b0000111111;
   81: result <= 10'b0000111111;
   82: result <= 10'b0001000000;
   83: result <= 10'b0001000001;
   84: result <= 10'b0001000010;
   85: result <= 10'b0001000011;
   86: result <= 10'b0001000011;
   87: result <= 10'b0001000100;
   88: result <= 10'b0001000101;
   89: result <= 10'b0001000110;
   90: result <= 10'b0001000110;
   91: result <= 10'b0001000111;
   92: result <= 10'b0001001000;
   93: result <= 10'b0001001001;
   94: result <= 10'b0001001010;
   95: result <= 10'b0001001010;
   96: result <= 10'b0001001011;
   97: result <= 10'b0001001100;
   98: result <= 10'b0001001101;
   99: result <= 10'b0001001101;
   100: result <= 10'b0001001110;
   101: result <= 10'b0001001111;
   102: result <= 10'b0001010000;
   103: result <= 10'b0001010001;
   104: result <= 10'b0001010001;
   105: result <= 10'b0001010010;
   106: result <= 10'b0001010011;
   107: result <= 10'b0001010100;
   108: result <= 10'b0001010100;
   109: result <= 10'b0001010101;
   110: result <= 10'b0001010110;
   111: result <= 10'b0001010111;
   112: result <= 10'b0001011000;
   113: result <= 10'b0001011000;
   114: result <= 10'b0001011001;
   115: result <= 10'b0001011010;
   116: result <= 10'b0001011011;
   117: result <= 10'b0001011011;
   118: result <= 10'b0001011100;
   119: result <= 10'b0001011101;
   120: result <= 10'b0001011110;
   121: result <= 10'b0001011110;
   122: result <= 10'b0001011111;
   123: result <= 10'b0001100000;
   124: result <= 10'b0001100001;
   125: result <= 10'b0001100010;
   126: result <= 10'b0001100010;
   127: result <= 10'b0001100011;
   128: result <= 10'b0001100100;
   129: result <= 10'b0001100101;
   130: result <= 10'b0001100101;
   131: result <= 10'b0001100110;
   132: result <= 10'b0001100111;
   133: result <= 10'b0001101000;
   134: result <= 10'b0001101001;
   135: result <= 10'b0001101001;
   136: result <= 10'b0001101010;
   137: result <= 10'b0001101011;
   138: result <= 10'b0001101100;
   139: result <= 10'b0001101100;
   140: result <= 10'b0001101101;
   141: result <= 10'b0001101110;
   142: result <= 10'b0001101111;
   143: result <= 10'b0001101111;
   144: result <= 10'b0001110000;
   145: result <= 10'b0001110001;
   146: result <= 10'b0001110010;
   147: result <= 10'b0001110010;
   148: result <= 10'b0001110011;
   149: result <= 10'b0001110100;
   150: result <= 10'b0001110101;
   151: result <= 10'b0001110110;
   152: result <= 10'b0001110110;
   153: result <= 10'b0001110111;
   154: result <= 10'b0001111000;
   155: result <= 10'b0001111001;
   156: result <= 10'b0001111001;
   157: result <= 10'b0001111010;
   158: result <= 10'b0001111011;
   159: result <= 10'b0001111100;
   160: result <= 10'b0001111100;
   161: result <= 10'b0001111101;
   162: result <= 10'b0001111110;
   163: result <= 10'b0001111111;
   164: result <= 10'b0001111111;
   165: result <= 10'b0010000000;
   166: result <= 10'b0010000001;
   167: result <= 10'b0010000010;
   168: result <= 10'b0010000010;
   169: result <= 10'b0010000011;
   170: result <= 10'b0010000100;
   171: result <= 10'b0010000101;
   172: result <= 10'b0010000110;
   173: result <= 10'b0010000110;
   174: result <= 10'b0010000111;
   175: result <= 10'b0010001000;
   176: result <= 10'b0010001001;
   177: result <= 10'b0010001001;
   178: result <= 10'b0010001010;
   179: result <= 10'b0010001011;
   180: result <= 10'b0010001100;
   181: result <= 10'b0010001100;
   182: result <= 10'b0010001101;
   183: result <= 10'b0010001110;
   184: result <= 10'b0010001111;
   185: result <= 10'b0010001111;
   186: result <= 10'b0010010000;
   187: result <= 10'b0010010001;
   188: result <= 10'b0010010010;
   189: result <= 10'b0010010010;
   190: result <= 10'b0010010011;
   191: result <= 10'b0010010100;
   192: result <= 10'b0010010101;
   193: result <= 10'b0010010101;
   194: result <= 10'b0010010110;
   195: result <= 10'b0010010111;
   196: result <= 10'b0010011000;
   197: result <= 10'b0010011000;
   198: result <= 10'b0010011001;
   199: result <= 10'b0010011010;
   200: result <= 10'b0010011011;
   201: result <= 10'b0010011011;
   202: result <= 10'b0010011100;
   203: result <= 10'b0010011101;
   204: result <= 10'b0010011110;
   205: result <= 10'b0010011110;
   206: result <= 10'b0010011111;
   207: result <= 10'b0010100000;
   208: result <= 10'b0010100001;
   209: result <= 10'b0010100001;
   210: result <= 10'b0010100010;
   211: result <= 10'b0010100011;
   212: result <= 10'b0010100100;
   213: result <= 10'b0010100100;
   214: result <= 10'b0010100101;
   215: result <= 10'b0010100110;
   216: result <= 10'b0010100111;
   217: result <= 10'b0010100111;
   218: result <= 10'b0010101000;
   219: result <= 10'b0010101001;
   220: result <= 10'b0010101010;
   221: result <= 10'b0010101010;
   222: result <= 10'b0010101011;
   223: result <= 10'b0010101100;
   224: result <= 10'b0010101100;
   225: result <= 10'b0010101101;
   226: result <= 10'b0010101110;
   227: result <= 10'b0010101111;
   228: result <= 10'b0010101111;
   229: result <= 10'b0010110000;
   230: result <= 10'b0010110001;
   231: result <= 10'b0010110010;
   232: result <= 10'b0010110010;
   233: result <= 10'b0010110011;
   234: result <= 10'b0010110100;
   235: result <= 10'b0010110101;
   236: result <= 10'b0010110101;
   237: result <= 10'b0010110110;
   238: result <= 10'b0010110111;
   239: result <= 10'b0010111000;
   240: result <= 10'b0010111000;
   241: result <= 10'b0010111001;
   242: result <= 10'b0010111010;
   243: result <= 10'b0010111010;
   244: result <= 10'b0010111011;
   245: result <= 10'b0010111100;
   246: result <= 10'b0010111101;
   247: result <= 10'b0010111101;
   248: result <= 10'b0010111110;
   249: result <= 10'b0010111111;
   250: result <= 10'b0011000000;
   251: result <= 10'b0011000000;
   252: result <= 10'b0011000001;
   253: result <= 10'b0011000010;
   254: result <= 10'b0011000010;
   255: result <= 10'b0011000011;
   256: result <= 10'b0011000100;
   257: result <= 10'b0011000101;
   258: result <= 10'b0011000101;
   259: result <= 10'b0011000110;
   260: result <= 10'b0011000111;
   261: result <= 10'b0011001000;
   262: result <= 10'b0011001000;
   263: result <= 10'b0011001001;
   264: result <= 10'b0011001010;
   265: result <= 10'b0011001010;
   266: result <= 10'b0011001011;
   267: result <= 10'b0011001100;
   268: result <= 10'b0011001101;
   269: result <= 10'b0011001101;
   270: result <= 10'b0011001110;
   271: result <= 10'b0011001111;
   272: result <= 10'b0011001111;
   273: result <= 10'b0011010000;
   274: result <= 10'b0011010001;
   275: result <= 10'b0011010010;
   276: result <= 10'b0011010010;
   277: result <= 10'b0011010011;
   278: result <= 10'b0011010100;
   279: result <= 10'b0011010100;
   280: result <= 10'b0011010101;
   281: result <= 10'b0011010110;
   282: result <= 10'b0011010111;
   283: result <= 10'b0011010111;
   284: result <= 10'b0011011000;
   285: result <= 10'b0011011001;
   286: result <= 10'b0011011001;
   287: result <= 10'b0011011010;
   288: result <= 10'b0011011011;
   289: result <= 10'b0011011100;
   290: result <= 10'b0011011100;
   291: result <= 10'b0011011101;
   292: result <= 10'b0011011110;
   293: result <= 10'b0011011110;
   294: result <= 10'b0011011111;
   295: result <= 10'b0011100000;
   296: result <= 10'b0011100001;
   297: result <= 10'b0011100001;
   298: result <= 10'b0011100010;
   299: result <= 10'b0011100011;
   300: result <= 10'b0011100011;
   301: result <= 10'b0011100100;
   302: result <= 10'b0011100101;
   303: result <= 10'b0011100101;
   304: result <= 10'b0011100110;
   305: result <= 10'b0011100111;
   306: result <= 10'b0011101000;
   307: result <= 10'b0011101000;
   308: result <= 10'b0011101001;
   309: result <= 10'b0011101010;
   310: result <= 10'b0011101010;
   311: result <= 10'b0011101011;
   312: result <= 10'b0011101100;
   313: result <= 10'b0011101100;
   314: result <= 10'b0011101101;
   315: result <= 10'b0011101110;
   316: result <= 10'b0011101111;
   317: result <= 10'b0011101111;
   318: result <= 10'b0011110000;
   319: result <= 10'b0011110001;
   320: result <= 10'b0011110001;
   321: result <= 10'b0011110010;
   322: result <= 10'b0011110011;
   323: result <= 10'b0011110011;
   324: result <= 10'b0011110100;
   325: result <= 10'b0011110101;
   326: result <= 10'b0011110110;
   327: result <= 10'b0011110110;
   328: result <= 10'b0011110111;
   329: result <= 10'b0011111000;
   330: result <= 10'b0011111000;
   331: result <= 10'b0011111001;
   332: result <= 10'b0011111010;
   333: result <= 10'b0011111010;
   334: result <= 10'b0011111011;
   335: result <= 10'b0011111100;
   336: result <= 10'b0011111100;
   337: result <= 10'b0011111101;
   338: result <= 10'b0011111110;
   339: result <= 10'b0011111110;
   340: result <= 10'b0011111111;
   341: result <= 10'b0100000000;
   342: result <= 10'b0100000000;
   343: result <= 10'b0100000001;
   344: result <= 10'b0100000010;
   345: result <= 10'b0100000010;
   346: result <= 10'b0100000011;
   347: result <= 10'b0100000100;
   348: result <= 10'b0100000101;
   349: result <= 10'b0100000101;
   350: result <= 10'b0100000110;
   351: result <= 10'b0100000111;
   352: result <= 10'b0100000111;
   353: result <= 10'b0100001000;
   354: result <= 10'b0100001001;
   355: result <= 10'b0100001001;
   356: result <= 10'b0100001010;
   357: result <= 10'b0100001011;
   358: result <= 10'b0100001011;
   359: result <= 10'b0100001100;
   360: result <= 10'b0100001101;
   361: result <= 10'b0100001101;
   362: result <= 10'b0100001110;
   363: result <= 10'b0100001111;
   364: result <= 10'b0100001111;
   365: result <= 10'b0100010000;
   366: result <= 10'b0100010001;
   367: result <= 10'b0100010001;
   368: result <= 10'b0100010010;
   369: result <= 10'b0100010011;
   370: result <= 10'b0100010011;
   371: result <= 10'b0100010100;
   372: result <= 10'b0100010101;
   373: result <= 10'b0100010101;
   374: result <= 10'b0100010110;
   375: result <= 10'b0100010111;
   376: result <= 10'b0100010111;
   377: result <= 10'b0100011000;
   378: result <= 10'b0100011001;
   379: result <= 10'b0100011001;
   380: result <= 10'b0100011010;
   381: result <= 10'b0100011010;
   382: result <= 10'b0100011011;
   383: result <= 10'b0100011100;
   384: result <= 10'b0100011100;
   385: result <= 10'b0100011101;
   386: result <= 10'b0100011110;
   387: result <= 10'b0100011110;
   388: result <= 10'b0100011111;
   389: result <= 10'b0100100000;
   390: result <= 10'b0100100000;
   391: result <= 10'b0100100001;
   392: result <= 10'b0100100010;
   393: result <= 10'b0100100010;
   394: result <= 10'b0100100011;
   395: result <= 10'b0100100100;
   396: result <= 10'b0100100100;
   397: result <= 10'b0100100101;
   398: result <= 10'b0100100110;
   399: result <= 10'b0100100110;
   400: result <= 10'b0100100111;
   401: result <= 10'b0100100111;
   402: result <= 10'b0100101000;
   403: result <= 10'b0100101001;
   404: result <= 10'b0100101001;
   405: result <= 10'b0100101010;
   406: result <= 10'b0100101011;
   407: result <= 10'b0100101011;
   408: result <= 10'b0100101100;
   409: result <= 10'b0100101101;
   410: result <= 10'b0100101101;
   411: result <= 10'b0100101110;
   412: result <= 10'b0100101110;
   413: result <= 10'b0100101111;
   414: result <= 10'b0100110000;
   415: result <= 10'b0100110000;
   416: result <= 10'b0100110001;
   417: result <= 10'b0100110010;
   418: result <= 10'b0100110010;
   419: result <= 10'b0100110011;
   420: result <= 10'b0100110100;
   421: result <= 10'b0100110100;
   422: result <= 10'b0100110101;
   423: result <= 10'b0100110101;
   424: result <= 10'b0100110110;
   425: result <= 10'b0100110111;
   426: result <= 10'b0100110111;
   427: result <= 10'b0100111000;
   428: result <= 10'b0100111001;
   429: result <= 10'b0100111001;
   430: result <= 10'b0100111010;
   431: result <= 10'b0100111010;
   432: result <= 10'b0100111011;
   433: result <= 10'b0100111100;
   434: result <= 10'b0100111100;
   435: result <= 10'b0100111101;
   436: result <= 10'b0100111101;
   437: result <= 10'b0100111110;
   438: result <= 10'b0100111111;
   439: result <= 10'b0100111111;
   440: result <= 10'b0101000000;
   441: result <= 10'b0101000001;
   442: result <= 10'b0101000001;
   443: result <= 10'b0101000010;
   444: result <= 10'b0101000010;
   445: result <= 10'b0101000011;
   446: result <= 10'b0101000100;
   447: result <= 10'b0101000100;
   448: result <= 10'b0101000101;
   449: result <= 10'b0101000101;
   450: result <= 10'b0101000110;
   451: result <= 10'b0101000111;
   452: result <= 10'b0101000111;
   453: result <= 10'b0101001000;
   454: result <= 10'b0101001000;
   455: result <= 10'b0101001001;
   456: result <= 10'b0101001010;
   457: result <= 10'b0101001010;
   458: result <= 10'b0101001011;
   459: result <= 10'b0101001011;
   460: result <= 10'b0101001100;
   461: result <= 10'b0101001101;
   462: result <= 10'b0101001101;
   463: result <= 10'b0101001110;
   464: result <= 10'b0101001110;
   465: result <= 10'b0101001111;
   466: result <= 10'b0101010000;
   467: result <= 10'b0101010000;
   468: result <= 10'b0101010001;
   469: result <= 10'b0101010001;
   470: result <= 10'b0101010010;
   471: result <= 10'b0101010011;
   472: result <= 10'b0101010011;
   473: result <= 10'b0101010100;
   474: result <= 10'b0101010100;
   475: result <= 10'b0101010101;
   476: result <= 10'b0101010110;
   477: result <= 10'b0101010110;
   478: result <= 10'b0101010111;
   479: result <= 10'b0101010111;
   480: result <= 10'b0101011000;
   481: result <= 10'b0101011000;
   482: result <= 10'b0101011001;
   483: result <= 10'b0101011010;
   484: result <= 10'b0101011010;
   485: result <= 10'b0101011011;
   486: result <= 10'b0101011011;
   487: result <= 10'b0101011100;
   488: result <= 10'b0101011100;
   489: result <= 10'b0101011101;
   490: result <= 10'b0101011110;
   491: result <= 10'b0101011110;
   492: result <= 10'b0101011111;
   493: result <= 10'b0101011111;
   494: result <= 10'b0101100000;
   495: result <= 10'b0101100000;
   496: result <= 10'b0101100001;
   497: result <= 10'b0101100010;
   498: result <= 10'b0101100010;
   499: result <= 10'b0101100011;
   500: result <= 10'b0101100011;
   501: result <= 10'b0101100100;
   502: result <= 10'b0101100100;
   503: result <= 10'b0101100101;
   504: result <= 10'b0101100110;
   505: result <= 10'b0101100110;
   506: result <= 10'b0101100111;
   507: result <= 10'b0101100111;
   508: result <= 10'b0101101000;
   509: result <= 10'b0101101000;
   510: result <= 10'b0101101001;
   511: result <= 10'b0101101001;
   512: result <= 10'b0101101010;
   513: result <= 10'b0101101011;
   514: result <= 10'b0101101011;
   515: result <= 10'b0101101100;
   516: result <= 10'b0101101100;
   517: result <= 10'b0101101101;
   518: result <= 10'b0101101101;
   519: result <= 10'b0101101110;
   520: result <= 10'b0101101110;
   521: result <= 10'b0101101111;
   522: result <= 10'b0101110000;
   523: result <= 10'b0101110000;
   524: result <= 10'b0101110001;
   525: result <= 10'b0101110001;
   526: result <= 10'b0101110010;
   527: result <= 10'b0101110010;
   528: result <= 10'b0101110011;
   529: result <= 10'b0101110011;
   530: result <= 10'b0101110100;
   531: result <= 10'b0101110100;
   532: result <= 10'b0101110101;
   533: result <= 10'b0101110110;
   534: result <= 10'b0101110110;
   535: result <= 10'b0101110111;
   536: result <= 10'b0101110111;
   537: result <= 10'b0101111000;
   538: result <= 10'b0101111000;
   539: result <= 10'b0101111001;
   540: result <= 10'b0101111001;
   541: result <= 10'b0101111010;
   542: result <= 10'b0101111010;
   543: result <= 10'b0101111011;
   544: result <= 10'b0101111011;
   545: result <= 10'b0101111100;
   546: result <= 10'b0101111100;
   547: result <= 10'b0101111101;
   548: result <= 10'b0101111101;
   549: result <= 10'b0101111110;
   550: result <= 10'b0101111111;
   551: result <= 10'b0101111111;
   552: result <= 10'b0110000000;
   553: result <= 10'b0110000000;
   554: result <= 10'b0110000001;
   555: result <= 10'b0110000001;
   556: result <= 10'b0110000010;
   557: result <= 10'b0110000010;
   558: result <= 10'b0110000011;
   559: result <= 10'b0110000011;
   560: result <= 10'b0110000100;
   561: result <= 10'b0110000100;
   562: result <= 10'b0110000101;
   563: result <= 10'b0110000101;
   564: result <= 10'b0110000110;
   565: result <= 10'b0110000110;
   566: result <= 10'b0110000111;
   567: result <= 10'b0110000111;
   568: result <= 10'b0110001000;
   569: result <= 10'b0110001000;
   570: result <= 10'b0110001001;
   571: result <= 10'b0110001001;
   572: result <= 10'b0110001010;
   573: result <= 10'b0110001010;
   574: result <= 10'b0110001011;
   575: result <= 10'b0110001011;
   576: result <= 10'b0110001100;
   577: result <= 10'b0110001100;
   578: result <= 10'b0110001101;
   579: result <= 10'b0110001101;
   580: result <= 10'b0110001110;
   581: result <= 10'b0110001110;
   582: result <= 10'b0110001111;
   583: result <= 10'b0110001111;
   584: result <= 10'b0110010000;
   585: result <= 10'b0110010000;
   586: result <= 10'b0110010001;
   587: result <= 10'b0110010001;
   588: result <= 10'b0110010010;
   589: result <= 10'b0110010010;
   590: result <= 10'b0110010011;
   591: result <= 10'b0110010011;
   592: result <= 10'b0110010100;
   593: result <= 10'b0110010100;
   594: result <= 10'b0110010101;
   595: result <= 10'b0110010101;
   596: result <= 10'b0110010110;
   597: result <= 10'b0110010110;
   598: result <= 10'b0110010111;
   599: result <= 10'b0110010111;
   600: result <= 10'b0110010111;
   601: result <= 10'b0110011000;
   602: result <= 10'b0110011000;
   603: result <= 10'b0110011001;
   604: result <= 10'b0110011001;
   605: result <= 10'b0110011010;
   606: result <= 10'b0110011010;
   607: result <= 10'b0110011011;
   608: result <= 10'b0110011011;
   609: result <= 10'b0110011100;
   610: result <= 10'b0110011100;
   611: result <= 10'b0110011101;
   612: result <= 10'b0110011101;
   613: result <= 10'b0110011110;
   614: result <= 10'b0110011110;
   615: result <= 10'b0110011110;
   616: result <= 10'b0110011111;
   617: result <= 10'b0110011111;
   618: result <= 10'b0110100000;
   619: result <= 10'b0110100000;
   620: result <= 10'b0110100001;
   621: result <= 10'b0110100001;
   622: result <= 10'b0110100010;
   623: result <= 10'b0110100010;
   624: result <= 10'b0110100011;
   625: result <= 10'b0110100011;
   626: result <= 10'b0110100100;
   627: result <= 10'b0110100100;
   628: result <= 10'b0110100100;
   629: result <= 10'b0110100101;
   630: result <= 10'b0110100101;
   631: result <= 10'b0110100110;
   632: result <= 10'b0110100110;
   633: result <= 10'b0110100111;
   634: result <= 10'b0110100111;
   635: result <= 10'b0110101000;
   636: result <= 10'b0110101000;
   637: result <= 10'b0110101000;
   638: result <= 10'b0110101001;
   639: result <= 10'b0110101001;
   640: result <= 10'b0110101010;
   641: result <= 10'b0110101010;
   642: result <= 10'b0110101011;
   643: result <= 10'b0110101011;
   644: result <= 10'b0110101011;
   645: result <= 10'b0110101100;
   646: result <= 10'b0110101100;
   647: result <= 10'b0110101101;
   648: result <= 10'b0110101101;
   649: result <= 10'b0110101110;
   650: result <= 10'b0110101110;
   651: result <= 10'b0110101110;
   652: result <= 10'b0110101111;
   653: result <= 10'b0110101111;
   654: result <= 10'b0110110000;
   655: result <= 10'b0110110000;
   656: result <= 10'b0110110001;
   657: result <= 10'b0110110001;
   658: result <= 10'b0110110001;
   659: result <= 10'b0110110010;
   660: result <= 10'b0110110010;
   661: result <= 10'b0110110011;
   662: result <= 10'b0110110011;
   663: result <= 10'b0110110011;
   664: result <= 10'b0110110100;
   665: result <= 10'b0110110100;
   666: result <= 10'b0110110101;
   667: result <= 10'b0110110101;
   668: result <= 10'b0110110110;
   669: result <= 10'b0110110110;
   670: result <= 10'b0110110110;
   671: result <= 10'b0110110111;
   672: result <= 10'b0110110111;
   673: result <= 10'b0110111000;
   674: result <= 10'b0110111000;
   675: result <= 10'b0110111000;
   676: result <= 10'b0110111001;
   677: result <= 10'b0110111001;
   678: result <= 10'b0110111010;
   679: result <= 10'b0110111010;
   680: result <= 10'b0110111010;
   681: result <= 10'b0110111011;
   682: result <= 10'b0110111011;
   683: result <= 10'b0110111100;
   684: result <= 10'b0110111100;
   685: result <= 10'b0110111100;
   686: result <= 10'b0110111101;
   687: result <= 10'b0110111101;
   688: result <= 10'b0110111101;
   689: result <= 10'b0110111110;
   690: result <= 10'b0110111110;
   691: result <= 10'b0110111111;
   692: result <= 10'b0110111111;
   693: result <= 10'b0110111111;
   694: result <= 10'b0111000000;
   695: result <= 10'b0111000000;
   696: result <= 10'b0111000001;
   697: result <= 10'b0111000001;
   698: result <= 10'b0111000001;
   699: result <= 10'b0111000010;
   700: result <= 10'b0111000010;
   701: result <= 10'b0111000010;
   702: result <= 10'b0111000011;
   703: result <= 10'b0111000011;
   704: result <= 10'b0111000100;
   705: result <= 10'b0111000100;
   706: result <= 10'b0111000100;
   707: result <= 10'b0111000101;
   708: result <= 10'b0111000101;
   709: result <= 10'b0111000101;
   710: result <= 10'b0111000110;
   711: result <= 10'b0111000110;
   712: result <= 10'b0111000110;
   713: result <= 10'b0111000111;
   714: result <= 10'b0111000111;
   715: result <= 10'b0111001000;
   716: result <= 10'b0111001000;
   717: result <= 10'b0111001000;
   718: result <= 10'b0111001001;
   719: result <= 10'b0111001001;
   720: result <= 10'b0111001001;
   721: result <= 10'b0111001010;
   722: result <= 10'b0111001010;
   723: result <= 10'b0111001010;
   724: result <= 10'b0111001011;
   725: result <= 10'b0111001011;
   726: result <= 10'b0111001011;
   727: result <= 10'b0111001100;
   728: result <= 10'b0111001100;
   729: result <= 10'b0111001100;
   730: result <= 10'b0111001101;
   731: result <= 10'b0111001101;
   732: result <= 10'b0111001101;
   733: result <= 10'b0111001110;
   734: result <= 10'b0111001110;
   735: result <= 10'b0111001111;
   736: result <= 10'b0111001111;
   737: result <= 10'b0111001111;
   738: result <= 10'b0111010000;
   739: result <= 10'b0111010000;
   740: result <= 10'b0111010000;
   741: result <= 10'b0111010001;
   742: result <= 10'b0111010001;
   743: result <= 10'b0111010001;
   744: result <= 10'b0111010001;
   745: result <= 10'b0111010010;
   746: result <= 10'b0111010010;
   747: result <= 10'b0111010010;
   748: result <= 10'b0111010011;
   749: result <= 10'b0111010011;
   750: result <= 10'b0111010011;
   751: result <= 10'b0111010100;
   752: result <= 10'b0111010100;
   753: result <= 10'b0111010100;
   754: result <= 10'b0111010101;
   755: result <= 10'b0111010101;
   756: result <= 10'b0111010101;
   757: result <= 10'b0111010110;
   758: result <= 10'b0111010110;
   759: result <= 10'b0111010110;
   760: result <= 10'b0111010111;
   761: result <= 10'b0111010111;
   762: result <= 10'b0111010111;
   763: result <= 10'b0111011000;
   764: result <= 10'b0111011000;
   765: result <= 10'b0111011000;
   766: result <= 10'b0111011000;
   767: result <= 10'b0111011001;
   768: result <= 10'b0111011001;
   769: result <= 10'b0111011001;
   770: result <= 10'b0111011010;
   771: result <= 10'b0111011010;
   772: result <= 10'b0111011010;
   773: result <= 10'b0111011011;
   774: result <= 10'b0111011011;
   775: result <= 10'b0111011011;
   776: result <= 10'b0111011011;
   777: result <= 10'b0111011100;
   778: result <= 10'b0111011100;
   779: result <= 10'b0111011100;
   780: result <= 10'b0111011101;
   781: result <= 10'b0111011101;
   782: result <= 10'b0111011101;
   783: result <= 10'b0111011101;
   784: result <= 10'b0111011110;
   785: result <= 10'b0111011110;
   786: result <= 10'b0111011110;
   787: result <= 10'b0111011111;
   788: result <= 10'b0111011111;
   789: result <= 10'b0111011111;
   790: result <= 10'b0111011111;
   791: result <= 10'b0111100000;
   792: result <= 10'b0111100000;
   793: result <= 10'b0111100000;
   794: result <= 10'b0111100000;
   795: result <= 10'b0111100001;
   796: result <= 10'b0111100001;
   797: result <= 10'b0111100001;
   798: result <= 10'b0111100010;
   799: result <= 10'b0111100010;
   800: result <= 10'b0111100010;
   801: result <= 10'b0111100010;
   802: result <= 10'b0111100011;
   803: result <= 10'b0111100011;
   804: result <= 10'b0111100011;
   805: result <= 10'b0111100011;
   806: result <= 10'b0111100100;
   807: result <= 10'b0111100100;
   808: result <= 10'b0111100100;
   809: result <= 10'b0111100100;
   810: result <= 10'b0111100101;
   811: result <= 10'b0111100101;
   812: result <= 10'b0111100101;
   813: result <= 10'b0111100101;
   814: result <= 10'b0111100110;
   815: result <= 10'b0111100110;
   816: result <= 10'b0111100110;
   817: result <= 10'b0111100110;
   818: result <= 10'b0111100111;
   819: result <= 10'b0111100111;
   820: result <= 10'b0111100111;
   821: result <= 10'b0111100111;
   822: result <= 10'b0111101000;
   823: result <= 10'b0111101000;
   824: result <= 10'b0111101000;
   825: result <= 10'b0111101000;
   826: result <= 10'b0111101001;
   827: result <= 10'b0111101001;
   828: result <= 10'b0111101001;
   829: result <= 10'b0111101001;
   830: result <= 10'b0111101001;
   831: result <= 10'b0111101010;
   832: result <= 10'b0111101010;
   833: result <= 10'b0111101010;
   834: result <= 10'b0111101010;
   835: result <= 10'b0111101011;
   836: result <= 10'b0111101011;
   837: result <= 10'b0111101011;
   838: result <= 10'b0111101011;
   839: result <= 10'b0111101100;
   840: result <= 10'b0111101100;
   841: result <= 10'b0111101100;
   842: result <= 10'b0111101100;
   843: result <= 10'b0111101100;
   844: result <= 10'b0111101101;
   845: result <= 10'b0111101101;
   846: result <= 10'b0111101101;
   847: result <= 10'b0111101101;
   848: result <= 10'b0111101101;
   849: result <= 10'b0111101110;
   850: result <= 10'b0111101110;
   851: result <= 10'b0111101110;
   852: result <= 10'b0111101110;
   853: result <= 10'b0111101110;
   854: result <= 10'b0111101111;
   855: result <= 10'b0111101111;
   856: result <= 10'b0111101111;
   857: result <= 10'b0111101111;
   858: result <= 10'b0111101111;
   859: result <= 10'b0111110000;
   860: result <= 10'b0111110000;
   861: result <= 10'b0111110000;
   862: result <= 10'b0111110000;
   863: result <= 10'b0111110000;
   864: result <= 10'b0111110001;
   865: result <= 10'b0111110001;
   866: result <= 10'b0111110001;
   867: result <= 10'b0111110001;
   868: result <= 10'b0111110001;
   869: result <= 10'b0111110010;
   870: result <= 10'b0111110010;
   871: result <= 10'b0111110010;
   872: result <= 10'b0111110010;
   873: result <= 10'b0111110010;
   874: result <= 10'b0111110011;
   875: result <= 10'b0111110011;
   876: result <= 10'b0111110011;
   877: result <= 10'b0111110011;
   878: result <= 10'b0111110011;
   879: result <= 10'b0111110011;
   880: result <= 10'b0111110100;
   881: result <= 10'b0111110100;
   882: result <= 10'b0111110100;
   883: result <= 10'b0111110100;
   884: result <= 10'b0111110100;
   885: result <= 10'b0111110100;
   886: result <= 10'b0111110101;
   887: result <= 10'b0111110101;
   888: result <= 10'b0111110101;
   889: result <= 10'b0111110101;
   890: result <= 10'b0111110101;
   891: result <= 10'b0111110101;
   892: result <= 10'b0111110110;
   893: result <= 10'b0111110110;
   894: result <= 10'b0111110110;
   895: result <= 10'b0111110110;
   896: result <= 10'b0111110110;
   897: result <= 10'b0111110110;
   898: result <= 10'b0111110110;
   899: result <= 10'b0111110111;
   900: result <= 10'b0111110111;
   901: result <= 10'b0111110111;
   902: result <= 10'b0111110111;
   903: result <= 10'b0111110111;
   904: result <= 10'b0111110111;
   905: result <= 10'b0111110111;
   906: result <= 10'b0111111000;
   907: result <= 10'b0111111000;
   908: result <= 10'b0111111000;
   909: result <= 10'b0111111000;
   910: result <= 10'b0111111000;
   911: result <= 10'b0111111000;
   912: result <= 10'b0111111000;
   913: result <= 10'b0111111001;
   914: result <= 10'b0111111001;
   915: result <= 10'b0111111001;
   916: result <= 10'b0111111001;
   917: result <= 10'b0111111001;
   918: result <= 10'b0111111001;
   919: result <= 10'b0111111001;
   920: result <= 10'b0111111001;
   921: result <= 10'b0111111010;
   922: result <= 10'b0111111010;
   923: result <= 10'b0111111010;
   924: result <= 10'b0111111010;
   925: result <= 10'b0111111010;
   926: result <= 10'b0111111010;
   927: result <= 10'b0111111010;
   928: result <= 10'b0111111010;
   929: result <= 10'b0111111011;
   930: result <= 10'b0111111011;
   931: result <= 10'b0111111011;
   932: result <= 10'b0111111011;
   933: result <= 10'b0111111011;
   934: result <= 10'b0111111011;
   935: result <= 10'b0111111011;
   936: result <= 10'b0111111011;
   937: result <= 10'b0111111011;
   938: result <= 10'b0111111100;
   939: result <= 10'b0111111100;
   940: result <= 10'b0111111100;
   941: result <= 10'b0111111100;
   942: result <= 10'b0111111100;
   943: result <= 10'b0111111100;
   944: result <= 10'b0111111100;
   945: result <= 10'b0111111100;
   946: result <= 10'b0111111100;
   947: result <= 10'b0111111100;
   948: result <= 10'b0111111101;
   949: result <= 10'b0111111101;
   950: result <= 10'b0111111101;
   951: result <= 10'b0111111101;
   952: result <= 10'b0111111101;
   953: result <= 10'b0111111101;
   954: result <= 10'b0111111101;
   955: result <= 10'b0111111101;
   956: result <= 10'b0111111101;
   957: result <= 10'b0111111101;
   958: result <= 10'b0111111101;
   959: result <= 10'b0111111101;
   960: result <= 10'b0111111110;
   961: result <= 10'b0111111110;
   962: result <= 10'b0111111110;
   963: result <= 10'b0111111110;
   964: result <= 10'b0111111110;
   965: result <= 10'b0111111110;
   966: result <= 10'b0111111110;
   967: result <= 10'b0111111110;
   968: result <= 10'b0111111110;
   969: result <= 10'b0111111110;
   970: result <= 10'b0111111110;
   971: result <= 10'b0111111110;
   972: result <= 10'b0111111110;
   973: result <= 10'b0111111110;
   974: result <= 10'b0111111110;
   975: result <= 10'b0111111111;
   976: result <= 10'b0111111111;
   977: result <= 10'b0111111111;
   978: result <= 10'b0111111111;
   979: result <= 10'b0111111111;
   980: result <= 10'b0111111111;
   981: result <= 10'b0111111111;
   982: result <= 10'b0111111111;
   983: result <= 10'b0111111111;
   984: result <= 10'b0111111111;
   985: result <= 10'b0111111111;
   986: result <= 10'b0111111111;
   987: result <= 10'b0111111111;
   988: result <= 10'b0111111111;
   989: result <= 10'b0111111111;
   990: result <= 10'b0111111111;
   991: result <= 10'b0111111111;
   992: result <= 10'b0111111111;
   993: result <= 10'b0111111111;
   994: result <= 10'b0111111111;
   995: result <= 10'b0111111111;
   996: result <= 10'b0111111111;
   997: result <= 10'b0111111111;
   998: result <= 10'b0111111111;
   999: result <= 10'b0111111111;
   1000: result <= 10'b0111111111;
   1001: result <= 10'b0111111111;
   1002: result <= 10'b0111111111;
   1003: result <= 10'b0111111111;
   1004: result <= 10'b0111111111;
   1005: result <= 10'b0111111111;
   1006: result <= 10'b0111111111;
   1007: result <= 10'b0111111111;
   1008: result <= 10'b0111111111;
   1009: result <= 10'b0111111111;
   1010: result <= 10'b0111111111;
   1011: result <= 10'b0111111111;
   1012: result <= 10'b0111111111;
   1013: result <= 10'b0111111111;
   1014: result <= 10'b0111111111;
   1015: result <= 10'b0111111111;
   1016: result <= 10'b0111111111;
   1017: result <= 10'b0111111111;
   1018: result <= 10'b0111111111;
   1019: result <= 10'b0111111111;
   1020: result <= 10'b0111111111;
   1021: result <= 10'b0111111111;
   1022: result <= 10'b0111111111;
   1023: result <= 10'b0111111111;
   1024: result <= 10'b0111111111;
   1025: result <= 10'b0111111111;
   1026: result <= 10'b0111111111;
   1027: result <= 10'b0111111111;
   1028: result <= 10'b0111111111;
   1029: result <= 10'b0111111111;
   1030: result <= 10'b0111111111;
   1031: result <= 10'b0111111111;
   1032: result <= 10'b0111111111;
   1033: result <= 10'b0111111111;
   1034: result <= 10'b0111111111;
   1035: result <= 10'b0111111111;
   1036: result <= 10'b0111111111;
   1037: result <= 10'b0111111111;
   1038: result <= 10'b0111111111;
   1039: result <= 10'b0111111111;
   1040: result <= 10'b0111111111;
   1041: result <= 10'b0111111111;
   1042: result <= 10'b0111111111;
   1043: result <= 10'b0111111111;
   1044: result <= 10'b0111111111;
   1045: result <= 10'b0111111111;
   1046: result <= 10'b0111111111;
   1047: result <= 10'b0111111111;
   1048: result <= 10'b0111111111;
   1049: result <= 10'b0111111111;
   1050: result <= 10'b0111111111;
   1051: result <= 10'b0111111111;
   1052: result <= 10'b0111111111;
   1053: result <= 10'b0111111111;
   1054: result <= 10'b0111111111;
   1055: result <= 10'b0111111111;
   1056: result <= 10'b0111111111;
   1057: result <= 10'b0111111111;
   1058: result <= 10'b0111111111;
   1059: result <= 10'b0111111111;
   1060: result <= 10'b0111111111;
   1061: result <= 10'b0111111111;
   1062: result <= 10'b0111111111;
   1063: result <= 10'b0111111111;
   1064: result <= 10'b0111111111;
   1065: result <= 10'b0111111111;
   1066: result <= 10'b0111111111;
   1067: result <= 10'b0111111111;
   1068: result <= 10'b0111111111;
   1069: result <= 10'b0111111111;
   1070: result <= 10'b0111111111;
   1071: result <= 10'b0111111111;
   1072: result <= 10'b0111111111;
   1073: result <= 10'b0111111111;
   1074: result <= 10'b0111111110;
   1075: result <= 10'b0111111110;
   1076: result <= 10'b0111111110;
   1077: result <= 10'b0111111110;
   1078: result <= 10'b0111111110;
   1079: result <= 10'b0111111110;
   1080: result <= 10'b0111111110;
   1081: result <= 10'b0111111110;
   1082: result <= 10'b0111111110;
   1083: result <= 10'b0111111110;
   1084: result <= 10'b0111111110;
   1085: result <= 10'b0111111110;
   1086: result <= 10'b0111111110;
   1087: result <= 10'b0111111110;
   1088: result <= 10'b0111111110;
   1089: result <= 10'b0111111101;
   1090: result <= 10'b0111111101;
   1091: result <= 10'b0111111101;
   1092: result <= 10'b0111111101;
   1093: result <= 10'b0111111101;
   1094: result <= 10'b0111111101;
   1095: result <= 10'b0111111101;
   1096: result <= 10'b0111111101;
   1097: result <= 10'b0111111101;
   1098: result <= 10'b0111111101;
   1099: result <= 10'b0111111101;
   1100: result <= 10'b0111111101;
   1101: result <= 10'b0111111100;
   1102: result <= 10'b0111111100;
   1103: result <= 10'b0111111100;
   1104: result <= 10'b0111111100;
   1105: result <= 10'b0111111100;
   1106: result <= 10'b0111111100;
   1107: result <= 10'b0111111100;
   1108: result <= 10'b0111111100;
   1109: result <= 10'b0111111100;
   1110: result <= 10'b0111111100;
   1111: result <= 10'b0111111011;
   1112: result <= 10'b0111111011;
   1113: result <= 10'b0111111011;
   1114: result <= 10'b0111111011;
   1115: result <= 10'b0111111011;
   1116: result <= 10'b0111111011;
   1117: result <= 10'b0111111011;
   1118: result <= 10'b0111111011;
   1119: result <= 10'b0111111011;
   1120: result <= 10'b0111111010;
   1121: result <= 10'b0111111010;
   1122: result <= 10'b0111111010;
   1123: result <= 10'b0111111010;
   1124: result <= 10'b0111111010;
   1125: result <= 10'b0111111010;
   1126: result <= 10'b0111111010;
   1127: result <= 10'b0111111010;
   1128: result <= 10'b0111111001;
   1129: result <= 10'b0111111001;
   1130: result <= 10'b0111111001;
   1131: result <= 10'b0111111001;
   1132: result <= 10'b0111111001;
   1133: result <= 10'b0111111001;
   1134: result <= 10'b0111111001;
   1135: result <= 10'b0111111001;
   1136: result <= 10'b0111111000;
   1137: result <= 10'b0111111000;
   1138: result <= 10'b0111111000;
   1139: result <= 10'b0111111000;
   1140: result <= 10'b0111111000;
   1141: result <= 10'b0111111000;
   1142: result <= 10'b0111111000;
   1143: result <= 10'b0111110111;
   1144: result <= 10'b0111110111;
   1145: result <= 10'b0111110111;
   1146: result <= 10'b0111110111;
   1147: result <= 10'b0111110111;
   1148: result <= 10'b0111110111;
   1149: result <= 10'b0111110111;
   1150: result <= 10'b0111110110;
   1151: result <= 10'b0111110110;
   1152: result <= 10'b0111110110;
   1153: result <= 10'b0111110110;
   1154: result <= 10'b0111110110;
   1155: result <= 10'b0111110110;
   1156: result <= 10'b0111110110;
   1157: result <= 10'b0111110101;
   1158: result <= 10'b0111110101;
   1159: result <= 10'b0111110101;
   1160: result <= 10'b0111110101;
   1161: result <= 10'b0111110101;
   1162: result <= 10'b0111110101;
   1163: result <= 10'b0111110100;
   1164: result <= 10'b0111110100;
   1165: result <= 10'b0111110100;
   1166: result <= 10'b0111110100;
   1167: result <= 10'b0111110100;
   1168: result <= 10'b0111110100;
   1169: result <= 10'b0111110011;
   1170: result <= 10'b0111110011;
   1171: result <= 10'b0111110011;
   1172: result <= 10'b0111110011;
   1173: result <= 10'b0111110011;
   1174: result <= 10'b0111110011;
   1175: result <= 10'b0111110010;
   1176: result <= 10'b0111110010;
   1177: result <= 10'b0111110010;
   1178: result <= 10'b0111110010;
   1179: result <= 10'b0111110010;
   1180: result <= 10'b0111110001;
   1181: result <= 10'b0111110001;
   1182: result <= 10'b0111110001;
   1183: result <= 10'b0111110001;
   1184: result <= 10'b0111110001;
   1185: result <= 10'b0111110000;
   1186: result <= 10'b0111110000;
   1187: result <= 10'b0111110000;
   1188: result <= 10'b0111110000;
   1189: result <= 10'b0111110000;
   1190: result <= 10'b0111101111;
   1191: result <= 10'b0111101111;
   1192: result <= 10'b0111101111;
   1193: result <= 10'b0111101111;
   1194: result <= 10'b0111101111;
   1195: result <= 10'b0111101110;
   1196: result <= 10'b0111101110;
   1197: result <= 10'b0111101110;
   1198: result <= 10'b0111101110;
   1199: result <= 10'b0111101110;
   1200: result <= 10'b0111101101;
   1201: result <= 10'b0111101101;
   1202: result <= 10'b0111101101;
   1203: result <= 10'b0111101101;
   1204: result <= 10'b0111101101;
   1205: result <= 10'b0111101100;
   1206: result <= 10'b0111101100;
   1207: result <= 10'b0111101100;
   1208: result <= 10'b0111101100;
   1209: result <= 10'b0111101100;
   1210: result <= 10'b0111101011;
   1211: result <= 10'b0111101011;
   1212: result <= 10'b0111101011;
   1213: result <= 10'b0111101011;
   1214: result <= 10'b0111101010;
   1215: result <= 10'b0111101010;
   1216: result <= 10'b0111101010;
   1217: result <= 10'b0111101010;
   1218: result <= 10'b0111101001;
   1219: result <= 10'b0111101001;
   1220: result <= 10'b0111101001;
   1221: result <= 10'b0111101001;
   1222: result <= 10'b0111101001;
   1223: result <= 10'b0111101000;
   1224: result <= 10'b0111101000;
   1225: result <= 10'b0111101000;
   1226: result <= 10'b0111101000;
   1227: result <= 10'b0111100111;
   1228: result <= 10'b0111100111;
   1229: result <= 10'b0111100111;
   1230: result <= 10'b0111100111;
   1231: result <= 10'b0111100110;
   1232: result <= 10'b0111100110;
   1233: result <= 10'b0111100110;
   1234: result <= 10'b0111100110;
   1235: result <= 10'b0111100101;
   1236: result <= 10'b0111100101;
   1237: result <= 10'b0111100101;
   1238: result <= 10'b0111100101;
   1239: result <= 10'b0111100100;
   1240: result <= 10'b0111100100;
   1241: result <= 10'b0111100100;
   1242: result <= 10'b0111100100;
   1243: result <= 10'b0111100011;
   1244: result <= 10'b0111100011;
   1245: result <= 10'b0111100011;
   1246: result <= 10'b0111100011;
   1247: result <= 10'b0111100010;
   1248: result <= 10'b0111100010;
   1249: result <= 10'b0111100010;
   1250: result <= 10'b0111100010;
   1251: result <= 10'b0111100001;
   1252: result <= 10'b0111100001;
   1253: result <= 10'b0111100001;
   1254: result <= 10'b0111100000;
   1255: result <= 10'b0111100000;
   1256: result <= 10'b0111100000;
   1257: result <= 10'b0111100000;
   1258: result <= 10'b0111011111;
   1259: result <= 10'b0111011111;
   1260: result <= 10'b0111011111;
   1261: result <= 10'b0111011111;
   1262: result <= 10'b0111011110;
   1263: result <= 10'b0111011110;
   1264: result <= 10'b0111011110;
   1265: result <= 10'b0111011101;
   1266: result <= 10'b0111011101;
   1267: result <= 10'b0111011101;
   1268: result <= 10'b0111011101;
   1269: result <= 10'b0111011100;
   1270: result <= 10'b0111011100;
   1271: result <= 10'b0111011100;
   1272: result <= 10'b0111011011;
   1273: result <= 10'b0111011011;
   1274: result <= 10'b0111011011;
   1275: result <= 10'b0111011011;
   1276: result <= 10'b0111011010;
   1277: result <= 10'b0111011010;
   1278: result <= 10'b0111011010;
   1279: result <= 10'b0111011001;
   1280: result <= 10'b0111011001;
   1281: result <= 10'b0111011001;
   1282: result <= 10'b0111011000;
   1283: result <= 10'b0111011000;
   1284: result <= 10'b0111011000;
   1285: result <= 10'b0111011000;
   1286: result <= 10'b0111010111;
   1287: result <= 10'b0111010111;
   1288: result <= 10'b0111010111;
   1289: result <= 10'b0111010110;
   1290: result <= 10'b0111010110;
   1291: result <= 10'b0111010110;
   1292: result <= 10'b0111010101;
   1293: result <= 10'b0111010101;
   1294: result <= 10'b0111010101;
   1295: result <= 10'b0111010100;
   1296: result <= 10'b0111010100;
   1297: result <= 10'b0111010100;
   1298: result <= 10'b0111010011;
   1299: result <= 10'b0111010011;
   1300: result <= 10'b0111010011;
   1301: result <= 10'b0111010010;
   1302: result <= 10'b0111010010;
   1303: result <= 10'b0111010010;
   1304: result <= 10'b0111010001;
   1305: result <= 10'b0111010001;
   1306: result <= 10'b0111010001;
   1307: result <= 10'b0111010001;
   1308: result <= 10'b0111010000;
   1309: result <= 10'b0111010000;
   1310: result <= 10'b0111010000;
   1311: result <= 10'b0111001111;
   1312: result <= 10'b0111001111;
   1313: result <= 10'b0111001111;
   1314: result <= 10'b0111001110;
   1315: result <= 10'b0111001110;
   1316: result <= 10'b0111001101;
   1317: result <= 10'b0111001101;
   1318: result <= 10'b0111001101;
   1319: result <= 10'b0111001100;
   1320: result <= 10'b0111001100;
   1321: result <= 10'b0111001100;
   1322: result <= 10'b0111001011;
   1323: result <= 10'b0111001011;
   1324: result <= 10'b0111001011;
   1325: result <= 10'b0111001010;
   1326: result <= 10'b0111001010;
   1327: result <= 10'b0111001010;
   1328: result <= 10'b0111001001;
   1329: result <= 10'b0111001001;
   1330: result <= 10'b0111001001;
   1331: result <= 10'b0111001000;
   1332: result <= 10'b0111001000;
   1333: result <= 10'b0111001000;
   1334: result <= 10'b0111000111;
   1335: result <= 10'b0111000111;
   1336: result <= 10'b0111000110;
   1337: result <= 10'b0111000110;
   1338: result <= 10'b0111000110;
   1339: result <= 10'b0111000101;
   1340: result <= 10'b0111000101;
   1341: result <= 10'b0111000101;
   1342: result <= 10'b0111000100;
   1343: result <= 10'b0111000100;
   1344: result <= 10'b0111000100;
   1345: result <= 10'b0111000011;
   1346: result <= 10'b0111000011;
   1347: result <= 10'b0111000010;
   1348: result <= 10'b0111000010;
   1349: result <= 10'b0111000010;
   1350: result <= 10'b0111000001;
   1351: result <= 10'b0111000001;
   1352: result <= 10'b0111000001;
   1353: result <= 10'b0111000000;
   1354: result <= 10'b0111000000;
   1355: result <= 10'b0110111111;
   1356: result <= 10'b0110111111;
   1357: result <= 10'b0110111111;
   1358: result <= 10'b0110111110;
   1359: result <= 10'b0110111110;
   1360: result <= 10'b0110111101;
   1361: result <= 10'b0110111101;
   1362: result <= 10'b0110111101;
   1363: result <= 10'b0110111100;
   1364: result <= 10'b0110111100;
   1365: result <= 10'b0110111100;
   1366: result <= 10'b0110111011;
   1367: result <= 10'b0110111011;
   1368: result <= 10'b0110111010;
   1369: result <= 10'b0110111010;
   1370: result <= 10'b0110111010;
   1371: result <= 10'b0110111001;
   1372: result <= 10'b0110111001;
   1373: result <= 10'b0110111000;
   1374: result <= 10'b0110111000;
   1375: result <= 10'b0110111000;
   1376: result <= 10'b0110110111;
   1377: result <= 10'b0110110111;
   1378: result <= 10'b0110110110;
   1379: result <= 10'b0110110110;
   1380: result <= 10'b0110110110;
   1381: result <= 10'b0110110101;
   1382: result <= 10'b0110110101;
   1383: result <= 10'b0110110100;
   1384: result <= 10'b0110110100;
   1385: result <= 10'b0110110011;
   1386: result <= 10'b0110110011;
   1387: result <= 10'b0110110011;
   1388: result <= 10'b0110110010;
   1389: result <= 10'b0110110010;
   1390: result <= 10'b0110110001;
   1391: result <= 10'b0110110001;
   1392: result <= 10'b0110110001;
   1393: result <= 10'b0110110000;
   1394: result <= 10'b0110110000;
   1395: result <= 10'b0110101111;
   1396: result <= 10'b0110101111;
   1397: result <= 10'b0110101110;
   1398: result <= 10'b0110101110;
   1399: result <= 10'b0110101110;
   1400: result <= 10'b0110101101;
   1401: result <= 10'b0110101101;
   1402: result <= 10'b0110101100;
   1403: result <= 10'b0110101100;
   1404: result <= 10'b0110101011;
   1405: result <= 10'b0110101011;
   1406: result <= 10'b0110101011;
   1407: result <= 10'b0110101010;
   1408: result <= 10'b0110101010;
   1409: result <= 10'b0110101001;
   1410: result <= 10'b0110101001;
   1411: result <= 10'b0110101000;
   1412: result <= 10'b0110101000;
   1413: result <= 10'b0110101000;
   1414: result <= 10'b0110100111;
   1415: result <= 10'b0110100111;
   1416: result <= 10'b0110100110;
   1417: result <= 10'b0110100110;
   1418: result <= 10'b0110100101;
   1419: result <= 10'b0110100101;
   1420: result <= 10'b0110100100;
   1421: result <= 10'b0110100100;
   1422: result <= 10'b0110100100;
   1423: result <= 10'b0110100011;
   1424: result <= 10'b0110100011;
   1425: result <= 10'b0110100010;
   1426: result <= 10'b0110100010;
   1427: result <= 10'b0110100001;
   1428: result <= 10'b0110100001;
   1429: result <= 10'b0110100000;
   1430: result <= 10'b0110100000;
   1431: result <= 10'b0110011111;
   1432: result <= 10'b0110011111;
   1433: result <= 10'b0110011110;
   1434: result <= 10'b0110011110;
   1435: result <= 10'b0110011110;
   1436: result <= 10'b0110011101;
   1437: result <= 10'b0110011101;
   1438: result <= 10'b0110011100;
   1439: result <= 10'b0110011100;
   1440: result <= 10'b0110011011;
   1441: result <= 10'b0110011011;
   1442: result <= 10'b0110011010;
   1443: result <= 10'b0110011010;
   1444: result <= 10'b0110011001;
   1445: result <= 10'b0110011001;
   1446: result <= 10'b0110011000;
   1447: result <= 10'b0110011000;
   1448: result <= 10'b0110010111;
   1449: result <= 10'b0110010111;
   1450: result <= 10'b0110010111;
   1451: result <= 10'b0110010110;
   1452: result <= 10'b0110010110;
   1453: result <= 10'b0110010101;
   1454: result <= 10'b0110010101;
   1455: result <= 10'b0110010100;
   1456: result <= 10'b0110010100;
   1457: result <= 10'b0110010011;
   1458: result <= 10'b0110010011;
   1459: result <= 10'b0110010010;
   1460: result <= 10'b0110010010;
   1461: result <= 10'b0110010001;
   1462: result <= 10'b0110010001;
   1463: result <= 10'b0110010000;
   1464: result <= 10'b0110010000;
   1465: result <= 10'b0110001111;
   1466: result <= 10'b0110001111;
   1467: result <= 10'b0110001110;
   1468: result <= 10'b0110001110;
   1469: result <= 10'b0110001101;
   1470: result <= 10'b0110001101;
   1471: result <= 10'b0110001100;
   1472: result <= 10'b0110001100;
   1473: result <= 10'b0110001011;
   1474: result <= 10'b0110001011;
   1475: result <= 10'b0110001010;
   1476: result <= 10'b0110001010;
   1477: result <= 10'b0110001001;
   1478: result <= 10'b0110001001;
   1479: result <= 10'b0110001000;
   1480: result <= 10'b0110001000;
   1481: result <= 10'b0110000111;
   1482: result <= 10'b0110000111;
   1483: result <= 10'b0110000110;
   1484: result <= 10'b0110000110;
   1485: result <= 10'b0110000101;
   1486: result <= 10'b0110000101;
   1487: result <= 10'b0110000100;
   1488: result <= 10'b0110000100;
   1489: result <= 10'b0110000011;
   1490: result <= 10'b0110000011;
   1491: result <= 10'b0110000010;
   1492: result <= 10'b0110000010;
   1493: result <= 10'b0110000001;
   1494: result <= 10'b0110000001;
   1495: result <= 10'b0110000000;
   1496: result <= 10'b0110000000;
   1497: result <= 10'b0101111111;
   1498: result <= 10'b0101111111;
   1499: result <= 10'b0101111110;
   1500: result <= 10'b0101111101;
   1501: result <= 10'b0101111101;
   1502: result <= 10'b0101111100;
   1503: result <= 10'b0101111100;
   1504: result <= 10'b0101111011;
   1505: result <= 10'b0101111011;
   1506: result <= 10'b0101111010;
   1507: result <= 10'b0101111010;
   1508: result <= 10'b0101111001;
   1509: result <= 10'b0101111001;
   1510: result <= 10'b0101111000;
   1511: result <= 10'b0101111000;
   1512: result <= 10'b0101110111;
   1513: result <= 10'b0101110111;
   1514: result <= 10'b0101110110;
   1515: result <= 10'b0101110110;
   1516: result <= 10'b0101110101;
   1517: result <= 10'b0101110100;
   1518: result <= 10'b0101110100;
   1519: result <= 10'b0101110011;
   1520: result <= 10'b0101110011;
   1521: result <= 10'b0101110010;
   1522: result <= 10'b0101110010;
   1523: result <= 10'b0101110001;
   1524: result <= 10'b0101110001;
   1525: result <= 10'b0101110000;
   1526: result <= 10'b0101110000;
   1527: result <= 10'b0101101111;
   1528: result <= 10'b0101101110;
   1529: result <= 10'b0101101110;
   1530: result <= 10'b0101101101;
   1531: result <= 10'b0101101101;
   1532: result <= 10'b0101101100;
   1533: result <= 10'b0101101100;
   1534: result <= 10'b0101101011;
   1535: result <= 10'b0101101011;
   1536: result <= 10'b0101101010;
   1537: result <= 10'b0101101001;
   1538: result <= 10'b0101101001;
   1539: result <= 10'b0101101000;
   1540: result <= 10'b0101101000;
   1541: result <= 10'b0101100111;
   1542: result <= 10'b0101100111;
   1543: result <= 10'b0101100110;
   1544: result <= 10'b0101100110;
   1545: result <= 10'b0101100101;
   1546: result <= 10'b0101100100;
   1547: result <= 10'b0101100100;
   1548: result <= 10'b0101100011;
   1549: result <= 10'b0101100011;
   1550: result <= 10'b0101100010;
   1551: result <= 10'b0101100010;
   1552: result <= 10'b0101100001;
   1553: result <= 10'b0101100000;
   1554: result <= 10'b0101100000;
   1555: result <= 10'b0101011111;
   1556: result <= 10'b0101011111;
   1557: result <= 10'b0101011110;
   1558: result <= 10'b0101011110;
   1559: result <= 10'b0101011101;
   1560: result <= 10'b0101011100;
   1561: result <= 10'b0101011100;
   1562: result <= 10'b0101011011;
   1563: result <= 10'b0101011011;
   1564: result <= 10'b0101011010;
   1565: result <= 10'b0101011010;
   1566: result <= 10'b0101011001;
   1567: result <= 10'b0101011000;
   1568: result <= 10'b0101011000;
   1569: result <= 10'b0101010111;
   1570: result <= 10'b0101010111;
   1571: result <= 10'b0101010110;
   1572: result <= 10'b0101010110;
   1573: result <= 10'b0101010101;
   1574: result <= 10'b0101010100;
   1575: result <= 10'b0101010100;
   1576: result <= 10'b0101010011;
   1577: result <= 10'b0101010011;
   1578: result <= 10'b0101010010;
   1579: result <= 10'b0101010001;
   1580: result <= 10'b0101010001;
   1581: result <= 10'b0101010000;
   1582: result <= 10'b0101010000;
   1583: result <= 10'b0101001111;
   1584: result <= 10'b0101001110;
   1585: result <= 10'b0101001110;
   1586: result <= 10'b0101001101;
   1587: result <= 10'b0101001101;
   1588: result <= 10'b0101001100;
   1589: result <= 10'b0101001011;
   1590: result <= 10'b0101001011;
   1591: result <= 10'b0101001010;
   1592: result <= 10'b0101001010;
   1593: result <= 10'b0101001001;
   1594: result <= 10'b0101001000;
   1595: result <= 10'b0101001000;
   1596: result <= 10'b0101000111;
   1597: result <= 10'b0101000111;
   1598: result <= 10'b0101000110;
   1599: result <= 10'b0101000101;
   1600: result <= 10'b0101000101;
   1601: result <= 10'b0101000100;
   1602: result <= 10'b0101000100;
   1603: result <= 10'b0101000011;
   1604: result <= 10'b0101000010;
   1605: result <= 10'b0101000010;
   1606: result <= 10'b0101000001;
   1607: result <= 10'b0101000001;
   1608: result <= 10'b0101000000;
   1609: result <= 10'b0100111111;
   1610: result <= 10'b0100111111;
   1611: result <= 10'b0100111110;
   1612: result <= 10'b0100111101;
   1613: result <= 10'b0100111101;
   1614: result <= 10'b0100111100;
   1615: result <= 10'b0100111100;
   1616: result <= 10'b0100111011;
   1617: result <= 10'b0100111010;
   1618: result <= 10'b0100111010;
   1619: result <= 10'b0100111001;
   1620: result <= 10'b0100111001;
   1621: result <= 10'b0100111000;
   1622: result <= 10'b0100110111;
   1623: result <= 10'b0100110111;
   1624: result <= 10'b0100110110;
   1625: result <= 10'b0100110101;
   1626: result <= 10'b0100110101;
   1627: result <= 10'b0100110100;
   1628: result <= 10'b0100110100;
   1629: result <= 10'b0100110011;
   1630: result <= 10'b0100110010;
   1631: result <= 10'b0100110010;
   1632: result <= 10'b0100110001;
   1633: result <= 10'b0100110000;
   1634: result <= 10'b0100110000;
   1635: result <= 10'b0100101111;
   1636: result <= 10'b0100101110;
   1637: result <= 10'b0100101110;
   1638: result <= 10'b0100101101;
   1639: result <= 10'b0100101101;
   1640: result <= 10'b0100101100;
   1641: result <= 10'b0100101011;
   1642: result <= 10'b0100101011;
   1643: result <= 10'b0100101010;
   1644: result <= 10'b0100101001;
   1645: result <= 10'b0100101001;
   1646: result <= 10'b0100101000;
   1647: result <= 10'b0100100111;
   1648: result <= 10'b0100100111;
   1649: result <= 10'b0100100110;
   1650: result <= 10'b0100100110;
   1651: result <= 10'b0100100101;
   1652: result <= 10'b0100100100;
   1653: result <= 10'b0100100100;
   1654: result <= 10'b0100100011;
   1655: result <= 10'b0100100010;
   1656: result <= 10'b0100100010;
   1657: result <= 10'b0100100001;
   1658: result <= 10'b0100100000;
   1659: result <= 10'b0100100000;
   1660: result <= 10'b0100011111;
   1661: result <= 10'b0100011110;
   1662: result <= 10'b0100011110;
   1663: result <= 10'b0100011101;
   1664: result <= 10'b0100011100;
   1665: result <= 10'b0100011100;
   1666: result <= 10'b0100011011;
   1667: result <= 10'b0100011010;
   1668: result <= 10'b0100011010;
   1669: result <= 10'b0100011001;
   1670: result <= 10'b0100011001;
   1671: result <= 10'b0100011000;
   1672: result <= 10'b0100010111;
   1673: result <= 10'b0100010111;
   1674: result <= 10'b0100010110;
   1675: result <= 10'b0100010101;
   1676: result <= 10'b0100010101;
   1677: result <= 10'b0100010100;
   1678: result <= 10'b0100010011;
   1679: result <= 10'b0100010011;
   1680: result <= 10'b0100010010;
   1681: result <= 10'b0100010001;
   1682: result <= 10'b0100010001;
   1683: result <= 10'b0100010000;
   1684: result <= 10'b0100001111;
   1685: result <= 10'b0100001111;
   1686: result <= 10'b0100001110;
   1687: result <= 10'b0100001101;
   1688: result <= 10'b0100001101;
   1689: result <= 10'b0100001100;
   1690: result <= 10'b0100001011;
   1691: result <= 10'b0100001011;
   1692: result <= 10'b0100001010;
   1693: result <= 10'b0100001001;
   1694: result <= 10'b0100001001;
   1695: result <= 10'b0100001000;
   1696: result <= 10'b0100000111;
   1697: result <= 10'b0100000111;
   1698: result <= 10'b0100000110;
   1699: result <= 10'b0100000101;
   1700: result <= 10'b0100000101;
   1701: result <= 10'b0100000100;
   1702: result <= 10'b0100000011;
   1703: result <= 10'b0100000010;
   1704: result <= 10'b0100000010;
   1705: result <= 10'b0100000001;
   1706: result <= 10'b0100000000;
   1707: result <= 10'b0100000000;
   1708: result <= 10'b0011111111;
   1709: result <= 10'b0011111110;
   1710: result <= 10'b0011111110;
   1711: result <= 10'b0011111101;
   1712: result <= 10'b0011111100;
   1713: result <= 10'b0011111100;
   1714: result <= 10'b0011111011;
   1715: result <= 10'b0011111010;
   1716: result <= 10'b0011111010;
   1717: result <= 10'b0011111001;
   1718: result <= 10'b0011111000;
   1719: result <= 10'b0011111000;
   1720: result <= 10'b0011110111;
   1721: result <= 10'b0011110110;
   1722: result <= 10'b0011110110;
   1723: result <= 10'b0011110101;
   1724: result <= 10'b0011110100;
   1725: result <= 10'b0011110011;
   1726: result <= 10'b0011110011;
   1727: result <= 10'b0011110010;
   1728: result <= 10'b0011110001;
   1729: result <= 10'b0011110001;
   1730: result <= 10'b0011110000;
   1731: result <= 10'b0011101111;
   1732: result <= 10'b0011101111;
   1733: result <= 10'b0011101110;
   1734: result <= 10'b0011101101;
   1735: result <= 10'b0011101100;
   1736: result <= 10'b0011101100;
   1737: result <= 10'b0011101011;
   1738: result <= 10'b0011101010;
   1739: result <= 10'b0011101010;
   1740: result <= 10'b0011101001;
   1741: result <= 10'b0011101000;
   1742: result <= 10'b0011101000;
   1743: result <= 10'b0011100111;
   1744: result <= 10'b0011100110;
   1745: result <= 10'b0011100101;
   1746: result <= 10'b0011100101;
   1747: result <= 10'b0011100100;
   1748: result <= 10'b0011100011;
   1749: result <= 10'b0011100011;
   1750: result <= 10'b0011100010;
   1751: result <= 10'b0011100001;
   1752: result <= 10'b0011100001;
   1753: result <= 10'b0011100000;
   1754: result <= 10'b0011011111;
   1755: result <= 10'b0011011110;
   1756: result <= 10'b0011011110;
   1757: result <= 10'b0011011101;
   1758: result <= 10'b0011011100;
   1759: result <= 10'b0011011100;
   1760: result <= 10'b0011011011;
   1761: result <= 10'b0011011010;
   1762: result <= 10'b0011011001;
   1763: result <= 10'b0011011001;
   1764: result <= 10'b0011011000;
   1765: result <= 10'b0011010111;
   1766: result <= 10'b0011010111;
   1767: result <= 10'b0011010110;
   1768: result <= 10'b0011010101;
   1769: result <= 10'b0011010100;
   1770: result <= 10'b0011010100;
   1771: result <= 10'b0011010011;
   1772: result <= 10'b0011010010;
   1773: result <= 10'b0011010010;
   1774: result <= 10'b0011010001;
   1775: result <= 10'b0011010000;
   1776: result <= 10'b0011001111;
   1777: result <= 10'b0011001111;
   1778: result <= 10'b0011001110;
   1779: result <= 10'b0011001101;
   1780: result <= 10'b0011001101;
   1781: result <= 10'b0011001100;
   1782: result <= 10'b0011001011;
   1783: result <= 10'b0011001010;
   1784: result <= 10'b0011001010;
   1785: result <= 10'b0011001001;
   1786: result <= 10'b0011001000;
   1787: result <= 10'b0011001000;
   1788: result <= 10'b0011000111;
   1789: result <= 10'b0011000110;
   1790: result <= 10'b0011000101;
   1791: result <= 10'b0011000101;
   1792: result <= 10'b0011000100;
   1793: result <= 10'b0011000011;
   1794: result <= 10'b0011000010;
   1795: result <= 10'b0011000010;
   1796: result <= 10'b0011000001;
   1797: result <= 10'b0011000000;
   1798: result <= 10'b0011000000;
   1799: result <= 10'b0010111111;
   1800: result <= 10'b0010111110;
   1801: result <= 10'b0010111101;
   1802: result <= 10'b0010111101;
   1803: result <= 10'b0010111100;
   1804: result <= 10'b0010111011;
   1805: result <= 10'b0010111010;
   1806: result <= 10'b0010111010;
   1807: result <= 10'b0010111001;
   1808: result <= 10'b0010111000;
   1809: result <= 10'b0010111000;
   1810: result <= 10'b0010110111;
   1811: result <= 10'b0010110110;
   1812: result <= 10'b0010110101;
   1813: result <= 10'b0010110101;
   1814: result <= 10'b0010110100;
   1815: result <= 10'b0010110011;
   1816: result <= 10'b0010110010;
   1817: result <= 10'b0010110010;
   1818: result <= 10'b0010110001;
   1819: result <= 10'b0010110000;
   1820: result <= 10'b0010101111;
   1821: result <= 10'b0010101111;
   1822: result <= 10'b0010101110;
   1823: result <= 10'b0010101101;
   1824: result <= 10'b0010101100;
   1825: result <= 10'b0010101100;
   1826: result <= 10'b0010101011;
   1827: result <= 10'b0010101010;
   1828: result <= 10'b0010101010;
   1829: result <= 10'b0010101001;
   1830: result <= 10'b0010101000;
   1831: result <= 10'b0010100111;
   1832: result <= 10'b0010100111;
   1833: result <= 10'b0010100110;
   1834: result <= 10'b0010100101;
   1835: result <= 10'b0010100100;
   1836: result <= 10'b0010100100;
   1837: result <= 10'b0010100011;
   1838: result <= 10'b0010100010;
   1839: result <= 10'b0010100001;
   1840: result <= 10'b0010100001;
   1841: result <= 10'b0010100000;
   1842: result <= 10'b0010011111;
   1843: result <= 10'b0010011110;
   1844: result <= 10'b0010011110;
   1845: result <= 10'b0010011101;
   1846: result <= 10'b0010011100;
   1847: result <= 10'b0010011011;
   1848: result <= 10'b0010011011;
   1849: result <= 10'b0010011010;
   1850: result <= 10'b0010011001;
   1851: result <= 10'b0010011000;
   1852: result <= 10'b0010011000;
   1853: result <= 10'b0010010111;
   1854: result <= 10'b0010010110;
   1855: result <= 10'b0010010101;
   1856: result <= 10'b0010010101;
   1857: result <= 10'b0010010100;
   1858: result <= 10'b0010010011;
   1859: result <= 10'b0010010010;
   1860: result <= 10'b0010010010;
   1861: result <= 10'b0010010001;
   1862: result <= 10'b0010010000;
   1863: result <= 10'b0010001111;
   1864: result <= 10'b0010001111;
   1865: result <= 10'b0010001110;
   1866: result <= 10'b0010001101;
   1867: result <= 10'b0010001100;
   1868: result <= 10'b0010001100;
   1869: result <= 10'b0010001011;
   1870: result <= 10'b0010001010;
   1871: result <= 10'b0010001001;
   1872: result <= 10'b0010001001;
   1873: result <= 10'b0010001000;
   1874: result <= 10'b0010000111;
   1875: result <= 10'b0010000110;
   1876: result <= 10'b0010000110;
   1877: result <= 10'b0010000101;
   1878: result <= 10'b0010000100;
   1879: result <= 10'b0010000011;
   1880: result <= 10'b0010000010;
   1881: result <= 10'b0010000010;
   1882: result <= 10'b0010000001;
   1883: result <= 10'b0010000000;
   1884: result <= 10'b0001111111;
   1885: result <= 10'b0001111111;
   1886: result <= 10'b0001111110;
   1887: result <= 10'b0001111101;
   1888: result <= 10'b0001111100;
   1889: result <= 10'b0001111100;
   1890: result <= 10'b0001111011;
   1891: result <= 10'b0001111010;
   1892: result <= 10'b0001111001;
   1893: result <= 10'b0001111001;
   1894: result <= 10'b0001111000;
   1895: result <= 10'b0001110111;
   1896: result <= 10'b0001110110;
   1897: result <= 10'b0001110110;
   1898: result <= 10'b0001110101;
   1899: result <= 10'b0001110100;
   1900: result <= 10'b0001110011;
   1901: result <= 10'b0001110010;
   1902: result <= 10'b0001110010;
   1903: result <= 10'b0001110001;
   1904: result <= 10'b0001110000;
   1905: result <= 10'b0001101111;
   1906: result <= 10'b0001101111;
   1907: result <= 10'b0001101110;
   1908: result <= 10'b0001101101;
   1909: result <= 10'b0001101100;
   1910: result <= 10'b0001101100;
   1911: result <= 10'b0001101011;
   1912: result <= 10'b0001101010;
   1913: result <= 10'b0001101001;
   1914: result <= 10'b0001101001;
   1915: result <= 10'b0001101000;
   1916: result <= 10'b0001100111;
   1917: result <= 10'b0001100110;
   1918: result <= 10'b0001100101;
   1919: result <= 10'b0001100101;
   1920: result <= 10'b0001100100;
   1921: result <= 10'b0001100011;
   1922: result <= 10'b0001100010;
   1923: result <= 10'b0001100010;
   1924: result <= 10'b0001100001;
   1925: result <= 10'b0001100000;
   1926: result <= 10'b0001011111;
   1927: result <= 10'b0001011110;
   1928: result <= 10'b0001011110;
   1929: result <= 10'b0001011101;
   1930: result <= 10'b0001011100;
   1931: result <= 10'b0001011011;
   1932: result <= 10'b0001011011;
   1933: result <= 10'b0001011010;
   1934: result <= 10'b0001011001;
   1935: result <= 10'b0001011000;
   1936: result <= 10'b0001011000;
   1937: result <= 10'b0001010111;
   1938: result <= 10'b0001010110;
   1939: result <= 10'b0001010101;
   1940: result <= 10'b0001010100;
   1941: result <= 10'b0001010100;
   1942: result <= 10'b0001010011;
   1943: result <= 10'b0001010010;
   1944: result <= 10'b0001010001;
   1945: result <= 10'b0001010001;
   1946: result <= 10'b0001010000;
   1947: result <= 10'b0001001111;
   1948: result <= 10'b0001001110;
   1949: result <= 10'b0001001101;
   1950: result <= 10'b0001001101;
   1951: result <= 10'b0001001100;
   1952: result <= 10'b0001001011;
   1953: result <= 10'b0001001010;
   1954: result <= 10'b0001001010;
   1955: result <= 10'b0001001001;
   1956: result <= 10'b0001001000;
   1957: result <= 10'b0001000111;
   1958: result <= 10'b0001000110;
   1959: result <= 10'b0001000110;
   1960: result <= 10'b0001000101;
   1961: result <= 10'b0001000100;
   1962: result <= 10'b0001000011;
   1963: result <= 10'b0001000011;
   1964: result <= 10'b0001000010;
   1965: result <= 10'b0001000001;
   1966: result <= 10'b0001000000;
   1967: result <= 10'b0000111111;
   1968: result <= 10'b0000111111;
   1969: result <= 10'b0000111110;
   1970: result <= 10'b0000111101;
   1971: result <= 10'b0000111100;
   1972: result <= 10'b0000111100;
   1973: result <= 10'b0000111011;
   1974: result <= 10'b0000111010;
   1975: result <= 10'b0000111001;
   1976: result <= 10'b0000111000;
   1977: result <= 10'b0000111000;
   1978: result <= 10'b0000110111;
   1979: result <= 10'b0000110110;
   1980: result <= 10'b0000110101;
   1981: result <= 10'b0000110101;
   1982: result <= 10'b0000110100;
   1983: result <= 10'b0000110011;
   1984: result <= 10'b0000110010;
   1985: result <= 10'b0000110001;
   1986: result <= 10'b0000110001;
   1987: result <= 10'b0000110000;
   1988: result <= 10'b0000101111;
   1989: result <= 10'b0000101110;
   1990: result <= 10'b0000101101;
   1991: result <= 10'b0000101101;
   1992: result <= 10'b0000101100;
   1993: result <= 10'b0000101011;
   1994: result <= 10'b0000101010;
   1995: result <= 10'b0000101010;
   1996: result <= 10'b0000101001;
   1997: result <= 10'b0000101000;
   1998: result <= 10'b0000100111;
   1999: result <= 10'b0000100110;
   2000: result <= 10'b0000100110;
   2001: result <= 10'b0000100101;
   2002: result <= 10'b0000100100;
   2003: result <= 10'b0000100011;
   2004: result <= 10'b0000100011;
   2005: result <= 10'b0000100010;
   2006: result <= 10'b0000100001;
   2007: result <= 10'b0000100000;
   2008: result <= 10'b0000011111;
   2009: result <= 10'b0000011111;
   2010: result <= 10'b0000011110;
   2011: result <= 10'b0000011101;
   2012: result <= 10'b0000011100;
   2013: result <= 10'b0000011011;
   2014: result <= 10'b0000011011;
   2015: result <= 10'b0000011010;
   2016: result <= 10'b0000011001;
   2017: result <= 10'b0000011000;
   2018: result <= 10'b0000011000;
   2019: result <= 10'b0000010111;
   2020: result <= 10'b0000010110;
   2021: result <= 10'b0000010101;
   2022: result <= 10'b0000010100;
   2023: result <= 10'b0000010100;
   2024: result <= 10'b0000010011;
   2025: result <= 10'b0000010010;
   2026: result <= 10'b0000010001;
   2027: result <= 10'b0000010000;
   2028: result <= 10'b0000010000;
   2029: result <= 10'b0000001111;
   2030: result <= 10'b0000001110;
   2031: result <= 10'b0000001101;
   2032: result <= 10'b0000001101;
   2033: result <= 10'b0000001100;
   2034: result <= 10'b0000001011;
   2035: result <= 10'b0000001010;
   2036: result <= 10'b0000001001;
   2037: result <= 10'b0000001001;
   2038: result <= 10'b0000001000;
   2039: result <= 10'b0000000111;
   2040: result <= 10'b0000000110;
   2041: result <= 10'b0000000101;
   2042: result <= 10'b0000000101;
   2043: result <= 10'b0000000100;
   2044: result <= 10'b0000000011;
   2045: result <= 10'b0000000010;
   2046: result <= 10'b0000000010;
   2047: result <= 10'b0000000001;
   2048: result <= 10'b0000000000;
   2049: result <= 10'b1111111111;
   2050: result <= 10'b1111111110;
   2051: result <= 10'b1111111110;
   2052: result <= 10'b1111111101;
   2053: result <= 10'b1111111100;
   2054: result <= 10'b1111111011;
   2055: result <= 10'b1111111011;
   2056: result <= 10'b1111111010;
   2057: result <= 10'b1111111001;
   2058: result <= 10'b1111111000;
   2059: result <= 10'b1111110111;
   2060: result <= 10'b1111110111;
   2061: result <= 10'b1111110110;
   2062: result <= 10'b1111110101;
   2063: result <= 10'b1111110100;
   2064: result <= 10'b1111110011;
   2065: result <= 10'b1111110011;
   2066: result <= 10'b1111110010;
   2067: result <= 10'b1111110001;
   2068: result <= 10'b1111110000;
   2069: result <= 10'b1111110000;
   2070: result <= 10'b1111101111;
   2071: result <= 10'b1111101110;
   2072: result <= 10'b1111101101;
   2073: result <= 10'b1111101100;
   2074: result <= 10'b1111101100;
   2075: result <= 10'b1111101011;
   2076: result <= 10'b1111101010;
   2077: result <= 10'b1111101001;
   2078: result <= 10'b1111101000;
   2079: result <= 10'b1111101000;
   2080: result <= 10'b1111100111;
   2081: result <= 10'b1111100110;
   2082: result <= 10'b1111100101;
   2083: result <= 10'b1111100101;
   2084: result <= 10'b1111100100;
   2085: result <= 10'b1111100011;
   2086: result <= 10'b1111100010;
   2087: result <= 10'b1111100001;
   2088: result <= 10'b1111100001;
   2089: result <= 10'b1111100000;
   2090: result <= 10'b1111011111;
   2091: result <= 10'b1111011110;
   2092: result <= 10'b1111011101;
   2093: result <= 10'b1111011101;
   2094: result <= 10'b1111011100;
   2095: result <= 10'b1111011011;
   2096: result <= 10'b1111011010;
   2097: result <= 10'b1111011010;
   2098: result <= 10'b1111011001;
   2099: result <= 10'b1111011000;
   2100: result <= 10'b1111010111;
   2101: result <= 10'b1111010110;
   2102: result <= 10'b1111010110;
   2103: result <= 10'b1111010101;
   2104: result <= 10'b1111010100;
   2105: result <= 10'b1111010011;
   2106: result <= 10'b1111010011;
   2107: result <= 10'b1111010010;
   2108: result <= 10'b1111010001;
   2109: result <= 10'b1111010000;
   2110: result <= 10'b1111001111;
   2111: result <= 10'b1111001111;
   2112: result <= 10'b1111001110;
   2113: result <= 10'b1111001101;
   2114: result <= 10'b1111001100;
   2115: result <= 10'b1111001011;
   2116: result <= 10'b1111001011;
   2117: result <= 10'b1111001010;
   2118: result <= 10'b1111001001;
   2119: result <= 10'b1111001000;
   2120: result <= 10'b1111001000;
   2121: result <= 10'b1111000111;
   2122: result <= 10'b1111000110;
   2123: result <= 10'b1111000101;
   2124: result <= 10'b1111000100;
   2125: result <= 10'b1111000100;
   2126: result <= 10'b1111000011;
   2127: result <= 10'b1111000010;
   2128: result <= 10'b1111000001;
   2129: result <= 10'b1111000001;
   2130: result <= 10'b1111000000;
   2131: result <= 10'b1110111111;
   2132: result <= 10'b1110111110;
   2133: result <= 10'b1110111101;
   2134: result <= 10'b1110111101;
   2135: result <= 10'b1110111100;
   2136: result <= 10'b1110111011;
   2137: result <= 10'b1110111010;
   2138: result <= 10'b1110111010;
   2139: result <= 10'b1110111001;
   2140: result <= 10'b1110111000;
   2141: result <= 10'b1110110111;
   2142: result <= 10'b1110110110;
   2143: result <= 10'b1110110110;
   2144: result <= 10'b1110110101;
   2145: result <= 10'b1110110100;
   2146: result <= 10'b1110110011;
   2147: result <= 10'b1110110011;
   2148: result <= 10'b1110110010;
   2149: result <= 10'b1110110001;
   2150: result <= 10'b1110110000;
   2151: result <= 10'b1110101111;
   2152: result <= 10'b1110101111;
   2153: result <= 10'b1110101110;
   2154: result <= 10'b1110101101;
   2155: result <= 10'b1110101100;
   2156: result <= 10'b1110101100;
   2157: result <= 10'b1110101011;
   2158: result <= 10'b1110101010;
   2159: result <= 10'b1110101001;
   2160: result <= 10'b1110101000;
   2161: result <= 10'b1110101000;
   2162: result <= 10'b1110100111;
   2163: result <= 10'b1110100110;
   2164: result <= 10'b1110100101;
   2165: result <= 10'b1110100101;
   2166: result <= 10'b1110100100;
   2167: result <= 10'b1110100011;
   2168: result <= 10'b1110100010;
   2169: result <= 10'b1110100010;
   2170: result <= 10'b1110100001;
   2171: result <= 10'b1110100000;
   2172: result <= 10'b1110011111;
   2173: result <= 10'b1110011110;
   2174: result <= 10'b1110011110;
   2175: result <= 10'b1110011101;
   2176: result <= 10'b1110011100;
   2177: result <= 10'b1110011011;
   2178: result <= 10'b1110011011;
   2179: result <= 10'b1110011010;
   2180: result <= 10'b1110011001;
   2181: result <= 10'b1110011000;
   2182: result <= 10'b1110010111;
   2183: result <= 10'b1110010111;
   2184: result <= 10'b1110010110;
   2185: result <= 10'b1110010101;
   2186: result <= 10'b1110010100;
   2187: result <= 10'b1110010100;
   2188: result <= 10'b1110010011;
   2189: result <= 10'b1110010010;
   2190: result <= 10'b1110010001;
   2191: result <= 10'b1110010001;
   2192: result <= 10'b1110010000;
   2193: result <= 10'b1110001111;
   2194: result <= 10'b1110001110;
   2195: result <= 10'b1110001110;
   2196: result <= 10'b1110001101;
   2197: result <= 10'b1110001100;
   2198: result <= 10'b1110001011;
   2199: result <= 10'b1110001010;
   2200: result <= 10'b1110001010;
   2201: result <= 10'b1110001001;
   2202: result <= 10'b1110001000;
   2203: result <= 10'b1110000111;
   2204: result <= 10'b1110000111;
   2205: result <= 10'b1110000110;
   2206: result <= 10'b1110000101;
   2207: result <= 10'b1110000100;
   2208: result <= 10'b1110000100;
   2209: result <= 10'b1110000011;
   2210: result <= 10'b1110000010;
   2211: result <= 10'b1110000001;
   2212: result <= 10'b1110000001;
   2213: result <= 10'b1110000000;
   2214: result <= 10'b1101111111;
   2215: result <= 10'b1101111110;
   2216: result <= 10'b1101111110;
   2217: result <= 10'b1101111101;
   2218: result <= 10'b1101111100;
   2219: result <= 10'b1101111011;
   2220: result <= 10'b1101111010;
   2221: result <= 10'b1101111010;
   2222: result <= 10'b1101111001;
   2223: result <= 10'b1101111000;
   2224: result <= 10'b1101110111;
   2225: result <= 10'b1101110111;
   2226: result <= 10'b1101110110;
   2227: result <= 10'b1101110101;
   2228: result <= 10'b1101110100;
   2229: result <= 10'b1101110100;
   2230: result <= 10'b1101110011;
   2231: result <= 10'b1101110010;
   2232: result <= 10'b1101110001;
   2233: result <= 10'b1101110001;
   2234: result <= 10'b1101110000;
   2235: result <= 10'b1101101111;
   2236: result <= 10'b1101101110;
   2237: result <= 10'b1101101110;
   2238: result <= 10'b1101101101;
   2239: result <= 10'b1101101100;
   2240: result <= 10'b1101101011;
   2241: result <= 10'b1101101011;
   2242: result <= 10'b1101101010;
   2243: result <= 10'b1101101001;
   2244: result <= 10'b1101101000;
   2245: result <= 10'b1101101000;
   2246: result <= 10'b1101100111;
   2247: result <= 10'b1101100110;
   2248: result <= 10'b1101100101;
   2249: result <= 10'b1101100101;
   2250: result <= 10'b1101100100;
   2251: result <= 10'b1101100011;
   2252: result <= 10'b1101100010;
   2253: result <= 10'b1101100010;
   2254: result <= 10'b1101100001;
   2255: result <= 10'b1101100000;
   2256: result <= 10'b1101011111;
   2257: result <= 10'b1101011111;
   2258: result <= 10'b1101011110;
   2259: result <= 10'b1101011101;
   2260: result <= 10'b1101011100;
   2261: result <= 10'b1101011100;
   2262: result <= 10'b1101011011;
   2263: result <= 10'b1101011010;
   2264: result <= 10'b1101011001;
   2265: result <= 10'b1101011001;
   2266: result <= 10'b1101011000;
   2267: result <= 10'b1101010111;
   2268: result <= 10'b1101010110;
   2269: result <= 10'b1101010110;
   2270: result <= 10'b1101010101;
   2271: result <= 10'b1101010100;
   2272: result <= 10'b1101010100;
   2273: result <= 10'b1101010011;
   2274: result <= 10'b1101010010;
   2275: result <= 10'b1101010001;
   2276: result <= 10'b1101010001;
   2277: result <= 10'b1101010000;
   2278: result <= 10'b1101001111;
   2279: result <= 10'b1101001110;
   2280: result <= 10'b1101001110;
   2281: result <= 10'b1101001101;
   2282: result <= 10'b1101001100;
   2283: result <= 10'b1101001011;
   2284: result <= 10'b1101001011;
   2285: result <= 10'b1101001010;
   2286: result <= 10'b1101001001;
   2287: result <= 10'b1101001000;
   2288: result <= 10'b1101001000;
   2289: result <= 10'b1101000111;
   2290: result <= 10'b1101000110;
   2291: result <= 10'b1101000110;
   2292: result <= 10'b1101000101;
   2293: result <= 10'b1101000100;
   2294: result <= 10'b1101000011;
   2295: result <= 10'b1101000011;
   2296: result <= 10'b1101000010;
   2297: result <= 10'b1101000001;
   2298: result <= 10'b1101000000;
   2299: result <= 10'b1101000000;
   2300: result <= 10'b1100111111;
   2301: result <= 10'b1100111110;
   2302: result <= 10'b1100111110;
   2303: result <= 10'b1100111101;
   2304: result <= 10'b1100111100;
   2305: result <= 10'b1100111011;
   2306: result <= 10'b1100111011;
   2307: result <= 10'b1100111010;
   2308: result <= 10'b1100111001;
   2309: result <= 10'b1100111000;
   2310: result <= 10'b1100111000;
   2311: result <= 10'b1100110111;
   2312: result <= 10'b1100110110;
   2313: result <= 10'b1100110110;
   2314: result <= 10'b1100110101;
   2315: result <= 10'b1100110100;
   2316: result <= 10'b1100110011;
   2317: result <= 10'b1100110011;
   2318: result <= 10'b1100110010;
   2319: result <= 10'b1100110001;
   2320: result <= 10'b1100110001;
   2321: result <= 10'b1100110000;
   2322: result <= 10'b1100101111;
   2323: result <= 10'b1100101110;
   2324: result <= 10'b1100101110;
   2325: result <= 10'b1100101101;
   2326: result <= 10'b1100101100;
   2327: result <= 10'b1100101100;
   2328: result <= 10'b1100101011;
   2329: result <= 10'b1100101010;
   2330: result <= 10'b1100101001;
   2331: result <= 10'b1100101001;
   2332: result <= 10'b1100101000;
   2333: result <= 10'b1100100111;
   2334: result <= 10'b1100100111;
   2335: result <= 10'b1100100110;
   2336: result <= 10'b1100100101;
   2337: result <= 10'b1100100100;
   2338: result <= 10'b1100100100;
   2339: result <= 10'b1100100011;
   2340: result <= 10'b1100100010;
   2341: result <= 10'b1100100010;
   2342: result <= 10'b1100100001;
   2343: result <= 10'b1100100000;
   2344: result <= 10'b1100011111;
   2345: result <= 10'b1100011111;
   2346: result <= 10'b1100011110;
   2347: result <= 10'b1100011101;
   2348: result <= 10'b1100011101;
   2349: result <= 10'b1100011100;
   2350: result <= 10'b1100011011;
   2351: result <= 10'b1100011011;
   2352: result <= 10'b1100011010;
   2353: result <= 10'b1100011001;
   2354: result <= 10'b1100011000;
   2355: result <= 10'b1100011000;
   2356: result <= 10'b1100010111;
   2357: result <= 10'b1100010110;
   2358: result <= 10'b1100010110;
   2359: result <= 10'b1100010101;
   2360: result <= 10'b1100010100;
   2361: result <= 10'b1100010100;
   2362: result <= 10'b1100010011;
   2363: result <= 10'b1100010010;
   2364: result <= 10'b1100010001;
   2365: result <= 10'b1100010001;
   2366: result <= 10'b1100010000;
   2367: result <= 10'b1100001111;
   2368: result <= 10'b1100001111;
   2369: result <= 10'b1100001110;
   2370: result <= 10'b1100001101;
   2371: result <= 10'b1100001101;
   2372: result <= 10'b1100001100;
   2373: result <= 10'b1100001011;
   2374: result <= 10'b1100001010;
   2375: result <= 10'b1100001010;
   2376: result <= 10'b1100001001;
   2377: result <= 10'b1100001000;
   2378: result <= 10'b1100001000;
   2379: result <= 10'b1100000111;
   2380: result <= 10'b1100000110;
   2381: result <= 10'b1100000110;
   2382: result <= 10'b1100000101;
   2383: result <= 10'b1100000100;
   2384: result <= 10'b1100000100;
   2385: result <= 10'b1100000011;
   2386: result <= 10'b1100000010;
   2387: result <= 10'b1100000010;
   2388: result <= 10'b1100000001;
   2389: result <= 10'b1100000000;
   2390: result <= 10'b1100000000;
   2391: result <= 10'b1011111111;
   2392: result <= 10'b1011111110;
   2393: result <= 10'b1011111110;
   2394: result <= 10'b1011111101;
   2395: result <= 10'b1011111100;
   2396: result <= 10'b1011111011;
   2397: result <= 10'b1011111011;
   2398: result <= 10'b1011111010;
   2399: result <= 10'b1011111001;
   2400: result <= 10'b1011111001;
   2401: result <= 10'b1011111000;
   2402: result <= 10'b1011110111;
   2403: result <= 10'b1011110111;
   2404: result <= 10'b1011110110;
   2405: result <= 10'b1011110101;
   2406: result <= 10'b1011110101;
   2407: result <= 10'b1011110100;
   2408: result <= 10'b1011110011;
   2409: result <= 10'b1011110011;
   2410: result <= 10'b1011110010;
   2411: result <= 10'b1011110001;
   2412: result <= 10'b1011110001;
   2413: result <= 10'b1011110000;
   2414: result <= 10'b1011101111;
   2415: result <= 10'b1011101111;
   2416: result <= 10'b1011101110;
   2417: result <= 10'b1011101101;
   2418: result <= 10'b1011101101;
   2419: result <= 10'b1011101100;
   2420: result <= 10'b1011101011;
   2421: result <= 10'b1011101011;
   2422: result <= 10'b1011101010;
   2423: result <= 10'b1011101001;
   2424: result <= 10'b1011101001;
   2425: result <= 10'b1011101000;
   2426: result <= 10'b1011100111;
   2427: result <= 10'b1011100111;
   2428: result <= 10'b1011100110;
   2429: result <= 10'b1011100110;
   2430: result <= 10'b1011100101;
   2431: result <= 10'b1011100100;
   2432: result <= 10'b1011100100;
   2433: result <= 10'b1011100011;
   2434: result <= 10'b1011100010;
   2435: result <= 10'b1011100010;
   2436: result <= 10'b1011100001;
   2437: result <= 10'b1011100000;
   2438: result <= 10'b1011100000;
   2439: result <= 10'b1011011111;
   2440: result <= 10'b1011011110;
   2441: result <= 10'b1011011110;
   2442: result <= 10'b1011011101;
   2443: result <= 10'b1011011100;
   2444: result <= 10'b1011011100;
   2445: result <= 10'b1011011011;
   2446: result <= 10'b1011011010;
   2447: result <= 10'b1011011010;
   2448: result <= 10'b1011011001;
   2449: result <= 10'b1011011001;
   2450: result <= 10'b1011011000;
   2451: result <= 10'b1011010111;
   2452: result <= 10'b1011010111;
   2453: result <= 10'b1011010110;
   2454: result <= 10'b1011010101;
   2455: result <= 10'b1011010101;
   2456: result <= 10'b1011010100;
   2457: result <= 10'b1011010011;
   2458: result <= 10'b1011010011;
   2459: result <= 10'b1011010010;
   2460: result <= 10'b1011010010;
   2461: result <= 10'b1011010001;
   2462: result <= 10'b1011010000;
   2463: result <= 10'b1011010000;
   2464: result <= 10'b1011001111;
   2465: result <= 10'b1011001110;
   2466: result <= 10'b1011001110;
   2467: result <= 10'b1011001101;
   2468: result <= 10'b1011001100;
   2469: result <= 10'b1011001100;
   2470: result <= 10'b1011001011;
   2471: result <= 10'b1011001011;
   2472: result <= 10'b1011001010;
   2473: result <= 10'b1011001001;
   2474: result <= 10'b1011001001;
   2475: result <= 10'b1011001000;
   2476: result <= 10'b1011000111;
   2477: result <= 10'b1011000111;
   2478: result <= 10'b1011000110;
   2479: result <= 10'b1011000110;
   2480: result <= 10'b1011000101;
   2481: result <= 10'b1011000100;
   2482: result <= 10'b1011000100;
   2483: result <= 10'b1011000011;
   2484: result <= 10'b1011000011;
   2485: result <= 10'b1011000010;
   2486: result <= 10'b1011000001;
   2487: result <= 10'b1011000001;
   2488: result <= 10'b1011000000;
   2489: result <= 10'b1010111111;
   2490: result <= 10'b1010111111;
   2491: result <= 10'b1010111110;
   2492: result <= 10'b1010111110;
   2493: result <= 10'b1010111101;
   2494: result <= 10'b1010111100;
   2495: result <= 10'b1010111100;
   2496: result <= 10'b1010111011;
   2497: result <= 10'b1010111011;
   2498: result <= 10'b1010111010;
   2499: result <= 10'b1010111001;
   2500: result <= 10'b1010111001;
   2501: result <= 10'b1010111000;
   2502: result <= 10'b1010111000;
   2503: result <= 10'b1010110111;
   2504: result <= 10'b1010110110;
   2505: result <= 10'b1010110110;
   2506: result <= 10'b1010110101;
   2507: result <= 10'b1010110101;
   2508: result <= 10'b1010110100;
   2509: result <= 10'b1010110011;
   2510: result <= 10'b1010110011;
   2511: result <= 10'b1010110010;
   2512: result <= 10'b1010110010;
   2513: result <= 10'b1010110001;
   2514: result <= 10'b1010110000;
   2515: result <= 10'b1010110000;
   2516: result <= 10'b1010101111;
   2517: result <= 10'b1010101111;
   2518: result <= 10'b1010101110;
   2519: result <= 10'b1010101101;
   2520: result <= 10'b1010101101;
   2521: result <= 10'b1010101100;
   2522: result <= 10'b1010101100;
   2523: result <= 10'b1010101011;
   2524: result <= 10'b1010101010;
   2525: result <= 10'b1010101010;
   2526: result <= 10'b1010101001;
   2527: result <= 10'b1010101001;
   2528: result <= 10'b1010101000;
   2529: result <= 10'b1010101000;
   2530: result <= 10'b1010100111;
   2531: result <= 10'b1010100110;
   2532: result <= 10'b1010100110;
   2533: result <= 10'b1010100101;
   2534: result <= 10'b1010100101;
   2535: result <= 10'b1010100100;
   2536: result <= 10'b1010100100;
   2537: result <= 10'b1010100011;
   2538: result <= 10'b1010100010;
   2539: result <= 10'b1010100010;
   2540: result <= 10'b1010100001;
   2541: result <= 10'b1010100001;
   2542: result <= 10'b1010100000;
   2543: result <= 10'b1010100000;
   2544: result <= 10'b1010011111;
   2545: result <= 10'b1010011110;
   2546: result <= 10'b1010011110;
   2547: result <= 10'b1010011101;
   2548: result <= 10'b1010011101;
   2549: result <= 10'b1010011100;
   2550: result <= 10'b1010011100;
   2551: result <= 10'b1010011011;
   2552: result <= 10'b1010011010;
   2553: result <= 10'b1010011010;
   2554: result <= 10'b1010011001;
   2555: result <= 10'b1010011001;
   2556: result <= 10'b1010011000;
   2557: result <= 10'b1010011000;
   2558: result <= 10'b1010010111;
   2559: result <= 10'b1010010111;
   2560: result <= 10'b1010010110;
   2561: result <= 10'b1010010101;
   2562: result <= 10'b1010010101;
   2563: result <= 10'b1010010100;
   2564: result <= 10'b1010010100;
   2565: result <= 10'b1010010011;
   2566: result <= 10'b1010010011;
   2567: result <= 10'b1010010010;
   2568: result <= 10'b1010010010;
   2569: result <= 10'b1010010001;
   2570: result <= 10'b1010010000;
   2571: result <= 10'b1010010000;
   2572: result <= 10'b1010001111;
   2573: result <= 10'b1010001111;
   2574: result <= 10'b1010001110;
   2575: result <= 10'b1010001110;
   2576: result <= 10'b1010001101;
   2577: result <= 10'b1010001101;
   2578: result <= 10'b1010001100;
   2579: result <= 10'b1010001100;
   2580: result <= 10'b1010001011;
   2581: result <= 10'b1010001010;
   2582: result <= 10'b1010001010;
   2583: result <= 10'b1010001001;
   2584: result <= 10'b1010001001;
   2585: result <= 10'b1010001000;
   2586: result <= 10'b1010001000;
   2587: result <= 10'b1010000111;
   2588: result <= 10'b1010000111;
   2589: result <= 10'b1010000110;
   2590: result <= 10'b1010000110;
   2591: result <= 10'b1010000101;
   2592: result <= 10'b1010000101;
   2593: result <= 10'b1010000100;
   2594: result <= 10'b1010000100;
   2595: result <= 10'b1010000011;
   2596: result <= 10'b1010000011;
   2597: result <= 10'b1010000010;
   2598: result <= 10'b1010000001;
   2599: result <= 10'b1010000001;
   2600: result <= 10'b1010000000;
   2601: result <= 10'b1010000000;
   2602: result <= 10'b1001111111;
   2603: result <= 10'b1001111111;
   2604: result <= 10'b1001111110;
   2605: result <= 10'b1001111110;
   2606: result <= 10'b1001111101;
   2607: result <= 10'b1001111101;
   2608: result <= 10'b1001111100;
   2609: result <= 10'b1001111100;
   2610: result <= 10'b1001111011;
   2611: result <= 10'b1001111011;
   2612: result <= 10'b1001111010;
   2613: result <= 10'b1001111010;
   2614: result <= 10'b1001111001;
   2615: result <= 10'b1001111001;
   2616: result <= 10'b1001111000;
   2617: result <= 10'b1001111000;
   2618: result <= 10'b1001110111;
   2619: result <= 10'b1001110111;
   2620: result <= 10'b1001110110;
   2621: result <= 10'b1001110110;
   2622: result <= 10'b1001110101;
   2623: result <= 10'b1001110101;
   2624: result <= 10'b1001110100;
   2625: result <= 10'b1001110100;
   2626: result <= 10'b1001110011;
   2627: result <= 10'b1001110011;
   2628: result <= 10'b1001110010;
   2629: result <= 10'b1001110010;
   2630: result <= 10'b1001110001;
   2631: result <= 10'b1001110001;
   2632: result <= 10'b1001110000;
   2633: result <= 10'b1001110000;
   2634: result <= 10'b1001101111;
   2635: result <= 10'b1001101111;
   2636: result <= 10'b1001101110;
   2637: result <= 10'b1001101110;
   2638: result <= 10'b1001101101;
   2639: result <= 10'b1001101101;
   2640: result <= 10'b1001101100;
   2641: result <= 10'b1001101100;
   2642: result <= 10'b1001101011;
   2643: result <= 10'b1001101011;
   2644: result <= 10'b1001101010;
   2645: result <= 10'b1001101010;
   2646: result <= 10'b1001101001;
   2647: result <= 10'b1001101001;
   2648: result <= 10'b1001101001;
   2649: result <= 10'b1001101000;
   2650: result <= 10'b1001101000;
   2651: result <= 10'b1001100111;
   2652: result <= 10'b1001100111;
   2653: result <= 10'b1001100110;
   2654: result <= 10'b1001100110;
   2655: result <= 10'b1001100101;
   2656: result <= 10'b1001100101;
   2657: result <= 10'b1001100100;
   2658: result <= 10'b1001100100;
   2659: result <= 10'b1001100011;
   2660: result <= 10'b1001100011;
   2661: result <= 10'b1001100010;
   2662: result <= 10'b1001100010;
   2663: result <= 10'b1001100010;
   2664: result <= 10'b1001100001;
   2665: result <= 10'b1001100001;
   2666: result <= 10'b1001100000;
   2667: result <= 10'b1001100000;
   2668: result <= 10'b1001011111;
   2669: result <= 10'b1001011111;
   2670: result <= 10'b1001011110;
   2671: result <= 10'b1001011110;
   2672: result <= 10'b1001011101;
   2673: result <= 10'b1001011101;
   2674: result <= 10'b1001011100;
   2675: result <= 10'b1001011100;
   2676: result <= 10'b1001011100;
   2677: result <= 10'b1001011011;
   2678: result <= 10'b1001011011;
   2679: result <= 10'b1001011010;
   2680: result <= 10'b1001011010;
   2681: result <= 10'b1001011001;
   2682: result <= 10'b1001011001;
   2683: result <= 10'b1001011000;
   2684: result <= 10'b1001011000;
   2685: result <= 10'b1001011000;
   2686: result <= 10'b1001010111;
   2687: result <= 10'b1001010111;
   2688: result <= 10'b1001010110;
   2689: result <= 10'b1001010110;
   2690: result <= 10'b1001010101;
   2691: result <= 10'b1001010101;
   2692: result <= 10'b1001010101;
   2693: result <= 10'b1001010100;
   2694: result <= 10'b1001010100;
   2695: result <= 10'b1001010011;
   2696: result <= 10'b1001010011;
   2697: result <= 10'b1001010010;
   2698: result <= 10'b1001010010;
   2699: result <= 10'b1001010010;
   2700: result <= 10'b1001010001;
   2701: result <= 10'b1001010001;
   2702: result <= 10'b1001010000;
   2703: result <= 10'b1001010000;
   2704: result <= 10'b1001001111;
   2705: result <= 10'b1001001111;
   2706: result <= 10'b1001001111;
   2707: result <= 10'b1001001110;
   2708: result <= 10'b1001001110;
   2709: result <= 10'b1001001101;
   2710: result <= 10'b1001001101;
   2711: result <= 10'b1001001101;
   2712: result <= 10'b1001001100;
   2713: result <= 10'b1001001100;
   2714: result <= 10'b1001001011;
   2715: result <= 10'b1001001011;
   2716: result <= 10'b1001001010;
   2717: result <= 10'b1001001010;
   2718: result <= 10'b1001001010;
   2719: result <= 10'b1001001001;
   2720: result <= 10'b1001001001;
   2721: result <= 10'b1001001000;
   2722: result <= 10'b1001001000;
   2723: result <= 10'b1001001000;
   2724: result <= 10'b1001000111;
   2725: result <= 10'b1001000111;
   2726: result <= 10'b1001000110;
   2727: result <= 10'b1001000110;
   2728: result <= 10'b1001000110;
   2729: result <= 10'b1001000101;
   2730: result <= 10'b1001000101;
   2731: result <= 10'b1001000100;
   2732: result <= 10'b1001000100;
   2733: result <= 10'b1001000100;
   2734: result <= 10'b1001000011;
   2735: result <= 10'b1001000011;
   2736: result <= 10'b1001000011;
   2737: result <= 10'b1001000010;
   2738: result <= 10'b1001000010;
   2739: result <= 10'b1001000001;
   2740: result <= 10'b1001000001;
   2741: result <= 10'b1001000001;
   2742: result <= 10'b1001000000;
   2743: result <= 10'b1001000000;
   2744: result <= 10'b1000111111;
   2745: result <= 10'b1000111111;
   2746: result <= 10'b1000111111;
   2747: result <= 10'b1000111110;
   2748: result <= 10'b1000111110;
   2749: result <= 10'b1000111110;
   2750: result <= 10'b1000111101;
   2751: result <= 10'b1000111101;
   2752: result <= 10'b1000111100;
   2753: result <= 10'b1000111100;
   2754: result <= 10'b1000111100;
   2755: result <= 10'b1000111011;
   2756: result <= 10'b1000111011;
   2757: result <= 10'b1000111011;
   2758: result <= 10'b1000111010;
   2759: result <= 10'b1000111010;
   2760: result <= 10'b1000111010;
   2761: result <= 10'b1000111001;
   2762: result <= 10'b1000111001;
   2763: result <= 10'b1000111000;
   2764: result <= 10'b1000111000;
   2765: result <= 10'b1000111000;
   2766: result <= 10'b1000110111;
   2767: result <= 10'b1000110111;
   2768: result <= 10'b1000110111;
   2769: result <= 10'b1000110110;
   2770: result <= 10'b1000110110;
   2771: result <= 10'b1000110110;
   2772: result <= 10'b1000110101;
   2773: result <= 10'b1000110101;
   2774: result <= 10'b1000110101;
   2775: result <= 10'b1000110100;
   2776: result <= 10'b1000110100;
   2777: result <= 10'b1000110100;
   2778: result <= 10'b1000110011;
   2779: result <= 10'b1000110011;
   2780: result <= 10'b1000110011;
   2781: result <= 10'b1000110010;
   2782: result <= 10'b1000110010;
   2783: result <= 10'b1000110001;
   2784: result <= 10'b1000110001;
   2785: result <= 10'b1000110001;
   2786: result <= 10'b1000110000;
   2787: result <= 10'b1000110000;
   2788: result <= 10'b1000110000;
   2789: result <= 10'b1000101111;
   2790: result <= 10'b1000101111;
   2791: result <= 10'b1000101111;
   2792: result <= 10'b1000101111;
   2793: result <= 10'b1000101110;
   2794: result <= 10'b1000101110;
   2795: result <= 10'b1000101110;
   2796: result <= 10'b1000101101;
   2797: result <= 10'b1000101101;
   2798: result <= 10'b1000101101;
   2799: result <= 10'b1000101100;
   2800: result <= 10'b1000101100;
   2801: result <= 10'b1000101100;
   2802: result <= 10'b1000101011;
   2803: result <= 10'b1000101011;
   2804: result <= 10'b1000101011;
   2805: result <= 10'b1000101010;
   2806: result <= 10'b1000101010;
   2807: result <= 10'b1000101010;
   2808: result <= 10'b1000101001;
   2809: result <= 10'b1000101001;
   2810: result <= 10'b1000101001;
   2811: result <= 10'b1000101000;
   2812: result <= 10'b1000101000;
   2813: result <= 10'b1000101000;
   2814: result <= 10'b1000101000;
   2815: result <= 10'b1000100111;
   2816: result <= 10'b1000100111;
   2817: result <= 10'b1000100111;
   2818: result <= 10'b1000100110;
   2819: result <= 10'b1000100110;
   2820: result <= 10'b1000100110;
   2821: result <= 10'b1000100101;
   2822: result <= 10'b1000100101;
   2823: result <= 10'b1000100101;
   2824: result <= 10'b1000100101;
   2825: result <= 10'b1000100100;
   2826: result <= 10'b1000100100;
   2827: result <= 10'b1000100100;
   2828: result <= 10'b1000100011;
   2829: result <= 10'b1000100011;
   2830: result <= 10'b1000100011;
   2831: result <= 10'b1000100011;
   2832: result <= 10'b1000100010;
   2833: result <= 10'b1000100010;
   2834: result <= 10'b1000100010;
   2835: result <= 10'b1000100001;
   2836: result <= 10'b1000100001;
   2837: result <= 10'b1000100001;
   2838: result <= 10'b1000100001;
   2839: result <= 10'b1000100000;
   2840: result <= 10'b1000100000;
   2841: result <= 10'b1000100000;
   2842: result <= 10'b1000100000;
   2843: result <= 10'b1000011111;
   2844: result <= 10'b1000011111;
   2845: result <= 10'b1000011111;
   2846: result <= 10'b1000011110;
   2847: result <= 10'b1000011110;
   2848: result <= 10'b1000011110;
   2849: result <= 10'b1000011110;
   2850: result <= 10'b1000011101;
   2851: result <= 10'b1000011101;
   2852: result <= 10'b1000011101;
   2853: result <= 10'b1000011101;
   2854: result <= 10'b1000011100;
   2855: result <= 10'b1000011100;
   2856: result <= 10'b1000011100;
   2857: result <= 10'b1000011100;
   2858: result <= 10'b1000011011;
   2859: result <= 10'b1000011011;
   2860: result <= 10'b1000011011;
   2861: result <= 10'b1000011011;
   2862: result <= 10'b1000011010;
   2863: result <= 10'b1000011010;
   2864: result <= 10'b1000011010;
   2865: result <= 10'b1000011010;
   2866: result <= 10'b1000011001;
   2867: result <= 10'b1000011001;
   2868: result <= 10'b1000011001;
   2869: result <= 10'b1000011001;
   2870: result <= 10'b1000011000;
   2871: result <= 10'b1000011000;
   2872: result <= 10'b1000011000;
   2873: result <= 10'b1000011000;
   2874: result <= 10'b1000010111;
   2875: result <= 10'b1000010111;
   2876: result <= 10'b1000010111;
   2877: result <= 10'b1000010111;
   2878: result <= 10'b1000010111;
   2879: result <= 10'b1000010110;
   2880: result <= 10'b1000010110;
   2881: result <= 10'b1000010110;
   2882: result <= 10'b1000010110;
   2883: result <= 10'b1000010101;
   2884: result <= 10'b1000010101;
   2885: result <= 10'b1000010101;
   2886: result <= 10'b1000010101;
   2887: result <= 10'b1000010100;
   2888: result <= 10'b1000010100;
   2889: result <= 10'b1000010100;
   2890: result <= 10'b1000010100;
   2891: result <= 10'b1000010100;
   2892: result <= 10'b1000010011;
   2893: result <= 10'b1000010011;
   2894: result <= 10'b1000010011;
   2895: result <= 10'b1000010011;
   2896: result <= 10'b1000010011;
   2897: result <= 10'b1000010010;
   2898: result <= 10'b1000010010;
   2899: result <= 10'b1000010010;
   2900: result <= 10'b1000010010;
   2901: result <= 10'b1000010010;
   2902: result <= 10'b1000010001;
   2903: result <= 10'b1000010001;
   2904: result <= 10'b1000010001;
   2905: result <= 10'b1000010001;
   2906: result <= 10'b1000010001;
   2907: result <= 10'b1000010000;
   2908: result <= 10'b1000010000;
   2909: result <= 10'b1000010000;
   2910: result <= 10'b1000010000;
   2911: result <= 10'b1000010000;
   2912: result <= 10'b1000001111;
   2913: result <= 10'b1000001111;
   2914: result <= 10'b1000001111;
   2915: result <= 10'b1000001111;
   2916: result <= 10'b1000001111;
   2917: result <= 10'b1000001110;
   2918: result <= 10'b1000001110;
   2919: result <= 10'b1000001110;
   2920: result <= 10'b1000001110;
   2921: result <= 10'b1000001110;
   2922: result <= 10'b1000001101;
   2923: result <= 10'b1000001101;
   2924: result <= 10'b1000001101;
   2925: result <= 10'b1000001101;
   2926: result <= 10'b1000001101;
   2927: result <= 10'b1000001101;
   2928: result <= 10'b1000001100;
   2929: result <= 10'b1000001100;
   2930: result <= 10'b1000001100;
   2931: result <= 10'b1000001100;
   2932: result <= 10'b1000001100;
   2933: result <= 10'b1000001100;
   2934: result <= 10'b1000001011;
   2935: result <= 10'b1000001011;
   2936: result <= 10'b1000001011;
   2937: result <= 10'b1000001011;
   2938: result <= 10'b1000001011;
   2939: result <= 10'b1000001011;
   2940: result <= 10'b1000001010;
   2941: result <= 10'b1000001010;
   2942: result <= 10'b1000001010;
   2943: result <= 10'b1000001010;
   2944: result <= 10'b1000001010;
   2945: result <= 10'b1000001010;
   2946: result <= 10'b1000001010;
   2947: result <= 10'b1000001001;
   2948: result <= 10'b1000001001;
   2949: result <= 10'b1000001001;
   2950: result <= 10'b1000001001;
   2951: result <= 10'b1000001001;
   2952: result <= 10'b1000001001;
   2953: result <= 10'b1000001001;
   2954: result <= 10'b1000001000;
   2955: result <= 10'b1000001000;
   2956: result <= 10'b1000001000;
   2957: result <= 10'b1000001000;
   2958: result <= 10'b1000001000;
   2959: result <= 10'b1000001000;
   2960: result <= 10'b1000001000;
   2961: result <= 10'b1000000111;
   2962: result <= 10'b1000000111;
   2963: result <= 10'b1000000111;
   2964: result <= 10'b1000000111;
   2965: result <= 10'b1000000111;
   2966: result <= 10'b1000000111;
   2967: result <= 10'b1000000111;
   2968: result <= 10'b1000000111;
   2969: result <= 10'b1000000110;
   2970: result <= 10'b1000000110;
   2971: result <= 10'b1000000110;
   2972: result <= 10'b1000000110;
   2973: result <= 10'b1000000110;
   2974: result <= 10'b1000000110;
   2975: result <= 10'b1000000110;
   2976: result <= 10'b1000000110;
   2977: result <= 10'b1000000101;
   2978: result <= 10'b1000000101;
   2979: result <= 10'b1000000101;
   2980: result <= 10'b1000000101;
   2981: result <= 10'b1000000101;
   2982: result <= 10'b1000000101;
   2983: result <= 10'b1000000101;
   2984: result <= 10'b1000000101;
   2985: result <= 10'b1000000101;
   2986: result <= 10'b1000000100;
   2987: result <= 10'b1000000100;
   2988: result <= 10'b1000000100;
   2989: result <= 10'b1000000100;
   2990: result <= 10'b1000000100;
   2991: result <= 10'b1000000100;
   2992: result <= 10'b1000000100;
   2993: result <= 10'b1000000100;
   2994: result <= 10'b1000000100;
   2995: result <= 10'b1000000100;
   2996: result <= 10'b1000000011;
   2997: result <= 10'b1000000011;
   2998: result <= 10'b1000000011;
   2999: result <= 10'b1000000011;
   3000: result <= 10'b1000000011;
   3001: result <= 10'b1000000011;
   3002: result <= 10'b1000000011;
   3003: result <= 10'b1000000011;
   3004: result <= 10'b1000000011;
   3005: result <= 10'b1000000011;
   3006: result <= 10'b1000000011;
   3007: result <= 10'b1000000011;
   3008: result <= 10'b1000000010;
   3009: result <= 10'b1000000010;
   3010: result <= 10'b1000000010;
   3011: result <= 10'b1000000010;
   3012: result <= 10'b1000000010;
   3013: result <= 10'b1000000010;
   3014: result <= 10'b1000000010;
   3015: result <= 10'b1000000010;
   3016: result <= 10'b1000000010;
   3017: result <= 10'b1000000010;
   3018: result <= 10'b1000000010;
   3019: result <= 10'b1000000010;
   3020: result <= 10'b1000000010;
   3021: result <= 10'b1000000010;
   3022: result <= 10'b1000000010;
   3023: result <= 10'b1000000001;
   3024: result <= 10'b1000000001;
   3025: result <= 10'b1000000001;
   3026: result <= 10'b1000000001;
   3027: result <= 10'b1000000001;
   3028: result <= 10'b1000000001;
   3029: result <= 10'b1000000001;
   3030: result <= 10'b1000000001;
   3031: result <= 10'b1000000001;
   3032: result <= 10'b1000000001;
   3033: result <= 10'b1000000001;
   3034: result <= 10'b1000000001;
   3035: result <= 10'b1000000001;
   3036: result <= 10'b1000000001;
   3037: result <= 10'b1000000001;
   3038: result <= 10'b1000000001;
   3039: result <= 10'b1000000001;
   3040: result <= 10'b1000000001;
   3041: result <= 10'b1000000001;
   3042: result <= 10'b1000000001;
   3043: result <= 10'b1000000001;
   3044: result <= 10'b1000000000;
   3045: result <= 10'b1000000000;
   3046: result <= 10'b1000000000;
   3047: result <= 10'b1000000000;
   3048: result <= 10'b1000000000;
   3049: result <= 10'b1000000000;
   3050: result <= 10'b1000000000;
   3051: result <= 10'b1000000000;
   3052: result <= 10'b1000000000;
   3053: result <= 10'b1000000000;
   3054: result <= 10'b1000000000;
   3055: result <= 10'b1000000000;
   3056: result <= 10'b1000000000;
   3057: result <= 10'b1000000000;
   3058: result <= 10'b1000000000;
   3059: result <= 10'b1000000000;
   3060: result <= 10'b1000000000;
   3061: result <= 10'b1000000000;
   3062: result <= 10'b1000000000;
   3063: result <= 10'b1000000000;
   3064: result <= 10'b1000000000;
   3065: result <= 10'b1000000000;
   3066: result <= 10'b1000000000;
   3067: result <= 10'b1000000000;
   3068: result <= 10'b1000000000;
   3069: result <= 10'b1000000000;
   3070: result <= 10'b1000000000;
   3071: result <= 10'b1000000000;
   3072: result <= 10'b1000000000;
   3073: result <= 10'b1000000000;
   3074: result <= 10'b1000000000;
   3075: result <= 10'b1000000000;
   3076: result <= 10'b1000000000;
   3077: result <= 10'b1000000000;
   3078: result <= 10'b1000000000;
   3079: result <= 10'b1000000000;
   3080: result <= 10'b1000000000;
   3081: result <= 10'b1000000000;
   3082: result <= 10'b1000000000;
   3083: result <= 10'b1000000000;
   3084: result <= 10'b1000000000;
   3085: result <= 10'b1000000000;
   3086: result <= 10'b1000000000;
   3087: result <= 10'b1000000000;
   3088: result <= 10'b1000000000;
   3089: result <= 10'b1000000000;
   3090: result <= 10'b1000000000;
   3091: result <= 10'b1000000000;
   3092: result <= 10'b1000000000;
   3093: result <= 10'b1000000000;
   3094: result <= 10'b1000000000;
   3095: result <= 10'b1000000000;
   3096: result <= 10'b1000000000;
   3097: result <= 10'b1000000000;
   3098: result <= 10'b1000000000;
   3099: result <= 10'b1000000000;
   3100: result <= 10'b1000000000;
   3101: result <= 10'b1000000001;
   3102: result <= 10'b1000000001;
   3103: result <= 10'b1000000001;
   3104: result <= 10'b1000000001;
   3105: result <= 10'b1000000001;
   3106: result <= 10'b1000000001;
   3107: result <= 10'b1000000001;
   3108: result <= 10'b1000000001;
   3109: result <= 10'b1000000001;
   3110: result <= 10'b1000000001;
   3111: result <= 10'b1000000001;
   3112: result <= 10'b1000000001;
   3113: result <= 10'b1000000001;
   3114: result <= 10'b1000000001;
   3115: result <= 10'b1000000001;
   3116: result <= 10'b1000000001;
   3117: result <= 10'b1000000001;
   3118: result <= 10'b1000000001;
   3119: result <= 10'b1000000001;
   3120: result <= 10'b1000000001;
   3121: result <= 10'b1000000001;
   3122: result <= 10'b1000000010;
   3123: result <= 10'b1000000010;
   3124: result <= 10'b1000000010;
   3125: result <= 10'b1000000010;
   3126: result <= 10'b1000000010;
   3127: result <= 10'b1000000010;
   3128: result <= 10'b1000000010;
   3129: result <= 10'b1000000010;
   3130: result <= 10'b1000000010;
   3131: result <= 10'b1000000010;
   3132: result <= 10'b1000000010;
   3133: result <= 10'b1000000010;
   3134: result <= 10'b1000000010;
   3135: result <= 10'b1000000010;
   3136: result <= 10'b1000000010;
   3137: result <= 10'b1000000011;
   3138: result <= 10'b1000000011;
   3139: result <= 10'b1000000011;
   3140: result <= 10'b1000000011;
   3141: result <= 10'b1000000011;
   3142: result <= 10'b1000000011;
   3143: result <= 10'b1000000011;
   3144: result <= 10'b1000000011;
   3145: result <= 10'b1000000011;
   3146: result <= 10'b1000000011;
   3147: result <= 10'b1000000011;
   3148: result <= 10'b1000000011;
   3149: result <= 10'b1000000100;
   3150: result <= 10'b1000000100;
   3151: result <= 10'b1000000100;
   3152: result <= 10'b1000000100;
   3153: result <= 10'b1000000100;
   3154: result <= 10'b1000000100;
   3155: result <= 10'b1000000100;
   3156: result <= 10'b1000000100;
   3157: result <= 10'b1000000100;
   3158: result <= 10'b1000000100;
   3159: result <= 10'b1000000101;
   3160: result <= 10'b1000000101;
   3161: result <= 10'b1000000101;
   3162: result <= 10'b1000000101;
   3163: result <= 10'b1000000101;
   3164: result <= 10'b1000000101;
   3165: result <= 10'b1000000101;
   3166: result <= 10'b1000000101;
   3167: result <= 10'b1000000101;
   3168: result <= 10'b1000000110;
   3169: result <= 10'b1000000110;
   3170: result <= 10'b1000000110;
   3171: result <= 10'b1000000110;
   3172: result <= 10'b1000000110;
   3173: result <= 10'b1000000110;
   3174: result <= 10'b1000000110;
   3175: result <= 10'b1000000110;
   3176: result <= 10'b1000000111;
   3177: result <= 10'b1000000111;
   3178: result <= 10'b1000000111;
   3179: result <= 10'b1000000111;
   3180: result <= 10'b1000000111;
   3181: result <= 10'b1000000111;
   3182: result <= 10'b1000000111;
   3183: result <= 10'b1000000111;
   3184: result <= 10'b1000001000;
   3185: result <= 10'b1000001000;
   3186: result <= 10'b1000001000;
   3187: result <= 10'b1000001000;
   3188: result <= 10'b1000001000;
   3189: result <= 10'b1000001000;
   3190: result <= 10'b1000001000;
   3191: result <= 10'b1000001001;
   3192: result <= 10'b1000001001;
   3193: result <= 10'b1000001001;
   3194: result <= 10'b1000001001;
   3195: result <= 10'b1000001001;
   3196: result <= 10'b1000001001;
   3197: result <= 10'b1000001001;
   3198: result <= 10'b1000001010;
   3199: result <= 10'b1000001010;
   3200: result <= 10'b1000001010;
   3201: result <= 10'b1000001010;
   3202: result <= 10'b1000001010;
   3203: result <= 10'b1000001010;
   3204: result <= 10'b1000001010;
   3205: result <= 10'b1000001011;
   3206: result <= 10'b1000001011;
   3207: result <= 10'b1000001011;
   3208: result <= 10'b1000001011;
   3209: result <= 10'b1000001011;
   3210: result <= 10'b1000001011;
   3211: result <= 10'b1000001100;
   3212: result <= 10'b1000001100;
   3213: result <= 10'b1000001100;
   3214: result <= 10'b1000001100;
   3215: result <= 10'b1000001100;
   3216: result <= 10'b1000001100;
   3217: result <= 10'b1000001101;
   3218: result <= 10'b1000001101;
   3219: result <= 10'b1000001101;
   3220: result <= 10'b1000001101;
   3221: result <= 10'b1000001101;
   3222: result <= 10'b1000001101;
   3223: result <= 10'b1000001110;
   3224: result <= 10'b1000001110;
   3225: result <= 10'b1000001110;
   3226: result <= 10'b1000001110;
   3227: result <= 10'b1000001110;
   3228: result <= 10'b1000001111;
   3229: result <= 10'b1000001111;
   3230: result <= 10'b1000001111;
   3231: result <= 10'b1000001111;
   3232: result <= 10'b1000001111;
   3233: result <= 10'b1000010000;
   3234: result <= 10'b1000010000;
   3235: result <= 10'b1000010000;
   3236: result <= 10'b1000010000;
   3237: result <= 10'b1000010000;
   3238: result <= 10'b1000010001;
   3239: result <= 10'b1000010001;
   3240: result <= 10'b1000010001;
   3241: result <= 10'b1000010001;
   3242: result <= 10'b1000010001;
   3243: result <= 10'b1000010010;
   3244: result <= 10'b1000010010;
   3245: result <= 10'b1000010010;
   3246: result <= 10'b1000010010;
   3247: result <= 10'b1000010010;
   3248: result <= 10'b1000010011;
   3249: result <= 10'b1000010011;
   3250: result <= 10'b1000010011;
   3251: result <= 10'b1000010011;
   3252: result <= 10'b1000010011;
   3253: result <= 10'b1000010100;
   3254: result <= 10'b1000010100;
   3255: result <= 10'b1000010100;
   3256: result <= 10'b1000010100;
   3257: result <= 10'b1000010100;
   3258: result <= 10'b1000010101;
   3259: result <= 10'b1000010101;
   3260: result <= 10'b1000010101;
   3261: result <= 10'b1000010101;
   3262: result <= 10'b1000010110;
   3263: result <= 10'b1000010110;
   3264: result <= 10'b1000010110;
   3265: result <= 10'b1000010110;
   3266: result <= 10'b1000010111;
   3267: result <= 10'b1000010111;
   3268: result <= 10'b1000010111;
   3269: result <= 10'b1000010111;
   3270: result <= 10'b1000010111;
   3271: result <= 10'b1000011000;
   3272: result <= 10'b1000011000;
   3273: result <= 10'b1000011000;
   3274: result <= 10'b1000011000;
   3275: result <= 10'b1000011001;
   3276: result <= 10'b1000011001;
   3277: result <= 10'b1000011001;
   3278: result <= 10'b1000011001;
   3279: result <= 10'b1000011010;
   3280: result <= 10'b1000011010;
   3281: result <= 10'b1000011010;
   3282: result <= 10'b1000011010;
   3283: result <= 10'b1000011011;
   3284: result <= 10'b1000011011;
   3285: result <= 10'b1000011011;
   3286: result <= 10'b1000011011;
   3287: result <= 10'b1000011100;
   3288: result <= 10'b1000011100;
   3289: result <= 10'b1000011100;
   3290: result <= 10'b1000011100;
   3291: result <= 10'b1000011101;
   3292: result <= 10'b1000011101;
   3293: result <= 10'b1000011101;
   3294: result <= 10'b1000011101;
   3295: result <= 10'b1000011110;
   3296: result <= 10'b1000011110;
   3297: result <= 10'b1000011110;
   3298: result <= 10'b1000011110;
   3299: result <= 10'b1000011111;
   3300: result <= 10'b1000011111;
   3301: result <= 10'b1000011111;
   3302: result <= 10'b1000100000;
   3303: result <= 10'b1000100000;
   3304: result <= 10'b1000100000;
   3305: result <= 10'b1000100000;
   3306: result <= 10'b1000100001;
   3307: result <= 10'b1000100001;
   3308: result <= 10'b1000100001;
   3309: result <= 10'b1000100001;
   3310: result <= 10'b1000100010;
   3311: result <= 10'b1000100010;
   3312: result <= 10'b1000100010;
   3313: result <= 10'b1000100011;
   3314: result <= 10'b1000100011;
   3315: result <= 10'b1000100011;
   3316: result <= 10'b1000100011;
   3317: result <= 10'b1000100100;
   3318: result <= 10'b1000100100;
   3319: result <= 10'b1000100100;
   3320: result <= 10'b1000100101;
   3321: result <= 10'b1000100101;
   3322: result <= 10'b1000100101;
   3323: result <= 10'b1000100101;
   3324: result <= 10'b1000100110;
   3325: result <= 10'b1000100110;
   3326: result <= 10'b1000100110;
   3327: result <= 10'b1000100111;
   3328: result <= 10'b1000100111;
   3329: result <= 10'b1000100111;
   3330: result <= 10'b1000101000;
   3331: result <= 10'b1000101000;
   3332: result <= 10'b1000101000;
   3333: result <= 10'b1000101000;
   3334: result <= 10'b1000101001;
   3335: result <= 10'b1000101001;
   3336: result <= 10'b1000101001;
   3337: result <= 10'b1000101010;
   3338: result <= 10'b1000101010;
   3339: result <= 10'b1000101010;
   3340: result <= 10'b1000101011;
   3341: result <= 10'b1000101011;
   3342: result <= 10'b1000101011;
   3343: result <= 10'b1000101100;
   3344: result <= 10'b1000101100;
   3345: result <= 10'b1000101100;
   3346: result <= 10'b1000101101;
   3347: result <= 10'b1000101101;
   3348: result <= 10'b1000101101;
   3349: result <= 10'b1000101110;
   3350: result <= 10'b1000101110;
   3351: result <= 10'b1000101110;
   3352: result <= 10'b1000101111;
   3353: result <= 10'b1000101111;
   3354: result <= 10'b1000101111;
   3355: result <= 10'b1000101111;
   3356: result <= 10'b1000110000;
   3357: result <= 10'b1000110000;
   3358: result <= 10'b1000110000;
   3359: result <= 10'b1000110001;
   3360: result <= 10'b1000110001;
   3361: result <= 10'b1000110001;
   3362: result <= 10'b1000110010;
   3363: result <= 10'b1000110010;
   3364: result <= 10'b1000110011;
   3365: result <= 10'b1000110011;
   3366: result <= 10'b1000110011;
   3367: result <= 10'b1000110100;
   3368: result <= 10'b1000110100;
   3369: result <= 10'b1000110100;
   3370: result <= 10'b1000110101;
   3371: result <= 10'b1000110101;
   3372: result <= 10'b1000110101;
   3373: result <= 10'b1000110110;
   3374: result <= 10'b1000110110;
   3375: result <= 10'b1000110110;
   3376: result <= 10'b1000110111;
   3377: result <= 10'b1000110111;
   3378: result <= 10'b1000110111;
   3379: result <= 10'b1000111000;
   3380: result <= 10'b1000111000;
   3381: result <= 10'b1000111000;
   3382: result <= 10'b1000111001;
   3383: result <= 10'b1000111001;
   3384: result <= 10'b1000111010;
   3385: result <= 10'b1000111010;
   3386: result <= 10'b1000111010;
   3387: result <= 10'b1000111011;
   3388: result <= 10'b1000111011;
   3389: result <= 10'b1000111011;
   3390: result <= 10'b1000111100;
   3391: result <= 10'b1000111100;
   3392: result <= 10'b1000111100;
   3393: result <= 10'b1000111101;
   3394: result <= 10'b1000111101;
   3395: result <= 10'b1000111110;
   3396: result <= 10'b1000111110;
   3397: result <= 10'b1000111110;
   3398: result <= 10'b1000111111;
   3399: result <= 10'b1000111111;
   3400: result <= 10'b1000111111;
   3401: result <= 10'b1001000000;
   3402: result <= 10'b1001000000;
   3403: result <= 10'b1001000001;
   3404: result <= 10'b1001000001;
   3405: result <= 10'b1001000001;
   3406: result <= 10'b1001000010;
   3407: result <= 10'b1001000010;
   3408: result <= 10'b1001000011;
   3409: result <= 10'b1001000011;
   3410: result <= 10'b1001000011;
   3411: result <= 10'b1001000100;
   3412: result <= 10'b1001000100;
   3413: result <= 10'b1001000100;
   3414: result <= 10'b1001000101;
   3415: result <= 10'b1001000101;
   3416: result <= 10'b1001000110;
   3417: result <= 10'b1001000110;
   3418: result <= 10'b1001000110;
   3419: result <= 10'b1001000111;
   3420: result <= 10'b1001000111;
   3421: result <= 10'b1001001000;
   3422: result <= 10'b1001001000;
   3423: result <= 10'b1001001000;
   3424: result <= 10'b1001001001;
   3425: result <= 10'b1001001001;
   3426: result <= 10'b1001001010;
   3427: result <= 10'b1001001010;
   3428: result <= 10'b1001001010;
   3429: result <= 10'b1001001011;
   3430: result <= 10'b1001001011;
   3431: result <= 10'b1001001100;
   3432: result <= 10'b1001001100;
   3433: result <= 10'b1001001101;
   3434: result <= 10'b1001001101;
   3435: result <= 10'b1001001101;
   3436: result <= 10'b1001001110;
   3437: result <= 10'b1001001110;
   3438: result <= 10'b1001001111;
   3439: result <= 10'b1001001111;
   3440: result <= 10'b1001001111;
   3441: result <= 10'b1001010000;
   3442: result <= 10'b1001010000;
   3443: result <= 10'b1001010001;
   3444: result <= 10'b1001010001;
   3445: result <= 10'b1001010010;
   3446: result <= 10'b1001010010;
   3447: result <= 10'b1001010010;
   3448: result <= 10'b1001010011;
   3449: result <= 10'b1001010011;
   3450: result <= 10'b1001010100;
   3451: result <= 10'b1001010100;
   3452: result <= 10'b1001010101;
   3453: result <= 10'b1001010101;
   3454: result <= 10'b1001010101;
   3455: result <= 10'b1001010110;
   3456: result <= 10'b1001010110;
   3457: result <= 10'b1001010111;
   3458: result <= 10'b1001010111;
   3459: result <= 10'b1001011000;
   3460: result <= 10'b1001011000;
   3461: result <= 10'b1001011000;
   3462: result <= 10'b1001011001;
   3463: result <= 10'b1001011001;
   3464: result <= 10'b1001011010;
   3465: result <= 10'b1001011010;
   3466: result <= 10'b1001011011;
   3467: result <= 10'b1001011011;
   3468: result <= 10'b1001011100;
   3469: result <= 10'b1001011100;
   3470: result <= 10'b1001011100;
   3471: result <= 10'b1001011101;
   3472: result <= 10'b1001011101;
   3473: result <= 10'b1001011110;
   3474: result <= 10'b1001011110;
   3475: result <= 10'b1001011111;
   3476: result <= 10'b1001011111;
   3477: result <= 10'b1001100000;
   3478: result <= 10'b1001100000;
   3479: result <= 10'b1001100001;
   3480: result <= 10'b1001100001;
   3481: result <= 10'b1001100010;
   3482: result <= 10'b1001100010;
   3483: result <= 10'b1001100010;
   3484: result <= 10'b1001100011;
   3485: result <= 10'b1001100011;
   3486: result <= 10'b1001100100;
   3487: result <= 10'b1001100100;
   3488: result <= 10'b1001100101;
   3489: result <= 10'b1001100101;
   3490: result <= 10'b1001100110;
   3491: result <= 10'b1001100110;
   3492: result <= 10'b1001100111;
   3493: result <= 10'b1001100111;
   3494: result <= 10'b1001101000;
   3495: result <= 10'b1001101000;
   3496: result <= 10'b1001101001;
   3497: result <= 10'b1001101001;
   3498: result <= 10'b1001101001;
   3499: result <= 10'b1001101010;
   3500: result <= 10'b1001101010;
   3501: result <= 10'b1001101011;
   3502: result <= 10'b1001101011;
   3503: result <= 10'b1001101100;
   3504: result <= 10'b1001101100;
   3505: result <= 10'b1001101101;
   3506: result <= 10'b1001101101;
   3507: result <= 10'b1001101110;
   3508: result <= 10'b1001101110;
   3509: result <= 10'b1001101111;
   3510: result <= 10'b1001101111;
   3511: result <= 10'b1001110000;
   3512: result <= 10'b1001110000;
   3513: result <= 10'b1001110001;
   3514: result <= 10'b1001110001;
   3515: result <= 10'b1001110010;
   3516: result <= 10'b1001110010;
   3517: result <= 10'b1001110011;
   3518: result <= 10'b1001110011;
   3519: result <= 10'b1001110100;
   3520: result <= 10'b1001110100;
   3521: result <= 10'b1001110101;
   3522: result <= 10'b1001110101;
   3523: result <= 10'b1001110110;
   3524: result <= 10'b1001110110;
   3525: result <= 10'b1001110111;
   3526: result <= 10'b1001110111;
   3527: result <= 10'b1001111000;
   3528: result <= 10'b1001111000;
   3529: result <= 10'b1001111001;
   3530: result <= 10'b1001111001;
   3531: result <= 10'b1001111010;
   3532: result <= 10'b1001111010;
   3533: result <= 10'b1001111011;
   3534: result <= 10'b1001111011;
   3535: result <= 10'b1001111100;
   3536: result <= 10'b1001111100;
   3537: result <= 10'b1001111101;
   3538: result <= 10'b1001111101;
   3539: result <= 10'b1001111110;
   3540: result <= 10'b1001111110;
   3541: result <= 10'b1001111111;
   3542: result <= 10'b1001111111;
   3543: result <= 10'b1010000000;
   3544: result <= 10'b1010000000;
   3545: result <= 10'b1010000001;
   3546: result <= 10'b1010000001;
   3547: result <= 10'b1010000010;
   3548: result <= 10'b1010000011;
   3549: result <= 10'b1010000011;
   3550: result <= 10'b1010000100;
   3551: result <= 10'b1010000100;
   3552: result <= 10'b1010000101;
   3553: result <= 10'b1010000101;
   3554: result <= 10'b1010000110;
   3555: result <= 10'b1010000110;
   3556: result <= 10'b1010000111;
   3557: result <= 10'b1010000111;
   3558: result <= 10'b1010001000;
   3559: result <= 10'b1010001000;
   3560: result <= 10'b1010001001;
   3561: result <= 10'b1010001001;
   3562: result <= 10'b1010001010;
   3563: result <= 10'b1010001010;
   3564: result <= 10'b1010001011;
   3565: result <= 10'b1010001100;
   3566: result <= 10'b1010001100;
   3567: result <= 10'b1010001101;
   3568: result <= 10'b1010001101;
   3569: result <= 10'b1010001110;
   3570: result <= 10'b1010001110;
   3571: result <= 10'b1010001111;
   3572: result <= 10'b1010001111;
   3573: result <= 10'b1010010000;
   3574: result <= 10'b1010010000;
   3575: result <= 10'b1010010001;
   3576: result <= 10'b1010010010;
   3577: result <= 10'b1010010010;
   3578: result <= 10'b1010010011;
   3579: result <= 10'b1010010011;
   3580: result <= 10'b1010010100;
   3581: result <= 10'b1010010100;
   3582: result <= 10'b1010010101;
   3583: result <= 10'b1010010101;
   3584: result <= 10'b1010010110;
   3585: result <= 10'b1010010111;
   3586: result <= 10'b1010010111;
   3587: result <= 10'b1010011000;
   3588: result <= 10'b1010011000;
   3589: result <= 10'b1010011001;
   3590: result <= 10'b1010011001;
   3591: result <= 10'b1010011010;
   3592: result <= 10'b1010011010;
   3593: result <= 10'b1010011011;
   3594: result <= 10'b1010011100;
   3595: result <= 10'b1010011100;
   3596: result <= 10'b1010011101;
   3597: result <= 10'b1010011101;
   3598: result <= 10'b1010011110;
   3599: result <= 10'b1010011110;
   3600: result <= 10'b1010011111;
   3601: result <= 10'b1010100000;
   3602: result <= 10'b1010100000;
   3603: result <= 10'b1010100001;
   3604: result <= 10'b1010100001;
   3605: result <= 10'b1010100010;
   3606: result <= 10'b1010100010;
   3607: result <= 10'b1010100011;
   3608: result <= 10'b1010100100;
   3609: result <= 10'b1010100100;
   3610: result <= 10'b1010100101;
   3611: result <= 10'b1010100101;
   3612: result <= 10'b1010100110;
   3613: result <= 10'b1010100110;
   3614: result <= 10'b1010100111;
   3615: result <= 10'b1010101000;
   3616: result <= 10'b1010101000;
   3617: result <= 10'b1010101001;
   3618: result <= 10'b1010101001;
   3619: result <= 10'b1010101010;
   3620: result <= 10'b1010101010;
   3621: result <= 10'b1010101011;
   3622: result <= 10'b1010101100;
   3623: result <= 10'b1010101100;
   3624: result <= 10'b1010101101;
   3625: result <= 10'b1010101101;
   3626: result <= 10'b1010101110;
   3627: result <= 10'b1010101111;
   3628: result <= 10'b1010101111;
   3629: result <= 10'b1010110000;
   3630: result <= 10'b1010110000;
   3631: result <= 10'b1010110001;
   3632: result <= 10'b1010110010;
   3633: result <= 10'b1010110010;
   3634: result <= 10'b1010110011;
   3635: result <= 10'b1010110011;
   3636: result <= 10'b1010110100;
   3637: result <= 10'b1010110101;
   3638: result <= 10'b1010110101;
   3639: result <= 10'b1010110110;
   3640: result <= 10'b1010110110;
   3641: result <= 10'b1010110111;
   3642: result <= 10'b1010111000;
   3643: result <= 10'b1010111000;
   3644: result <= 10'b1010111001;
   3645: result <= 10'b1010111001;
   3646: result <= 10'b1010111010;
   3647: result <= 10'b1010111011;
   3648: result <= 10'b1010111011;
   3649: result <= 10'b1010111100;
   3650: result <= 10'b1010111100;
   3651: result <= 10'b1010111101;
   3652: result <= 10'b1010111110;
   3653: result <= 10'b1010111110;
   3654: result <= 10'b1010111111;
   3655: result <= 10'b1010111111;
   3656: result <= 10'b1011000000;
   3657: result <= 10'b1011000001;
   3658: result <= 10'b1011000001;
   3659: result <= 10'b1011000010;
   3660: result <= 10'b1011000011;
   3661: result <= 10'b1011000011;
   3662: result <= 10'b1011000100;
   3663: result <= 10'b1011000100;
   3664: result <= 10'b1011000101;
   3665: result <= 10'b1011000110;
   3666: result <= 10'b1011000110;
   3667: result <= 10'b1011000111;
   3668: result <= 10'b1011000111;
   3669: result <= 10'b1011001000;
   3670: result <= 10'b1011001001;
   3671: result <= 10'b1011001001;
   3672: result <= 10'b1011001010;
   3673: result <= 10'b1011001011;
   3674: result <= 10'b1011001011;
   3675: result <= 10'b1011001100;
   3676: result <= 10'b1011001100;
   3677: result <= 10'b1011001101;
   3678: result <= 10'b1011001110;
   3679: result <= 10'b1011001110;
   3680: result <= 10'b1011001111;
   3681: result <= 10'b1011010000;
   3682: result <= 10'b1011010000;
   3683: result <= 10'b1011010001;
   3684: result <= 10'b1011010010;
   3685: result <= 10'b1011010010;
   3686: result <= 10'b1011010011;
   3687: result <= 10'b1011010011;
   3688: result <= 10'b1011010100;
   3689: result <= 10'b1011010101;
   3690: result <= 10'b1011010101;
   3691: result <= 10'b1011010110;
   3692: result <= 10'b1011010111;
   3693: result <= 10'b1011010111;
   3694: result <= 10'b1011011000;
   3695: result <= 10'b1011011001;
   3696: result <= 10'b1011011001;
   3697: result <= 10'b1011011010;
   3698: result <= 10'b1011011010;
   3699: result <= 10'b1011011011;
   3700: result <= 10'b1011011100;
   3701: result <= 10'b1011011100;
   3702: result <= 10'b1011011101;
   3703: result <= 10'b1011011110;
   3704: result <= 10'b1011011110;
   3705: result <= 10'b1011011111;
   3706: result <= 10'b1011100000;
   3707: result <= 10'b1011100000;
   3708: result <= 10'b1011100001;
   3709: result <= 10'b1011100010;
   3710: result <= 10'b1011100010;
   3711: result <= 10'b1011100011;
   3712: result <= 10'b1011100100;
   3713: result <= 10'b1011100100;
   3714: result <= 10'b1011100101;
   3715: result <= 10'b1011100110;
   3716: result <= 10'b1011100110;
   3717: result <= 10'b1011100111;
   3718: result <= 10'b1011100111;
   3719: result <= 10'b1011101000;
   3720: result <= 10'b1011101001;
   3721: result <= 10'b1011101001;
   3722: result <= 10'b1011101010;
   3723: result <= 10'b1011101011;
   3724: result <= 10'b1011101011;
   3725: result <= 10'b1011101100;
   3726: result <= 10'b1011101101;
   3727: result <= 10'b1011101101;
   3728: result <= 10'b1011101110;
   3729: result <= 10'b1011101111;
   3730: result <= 10'b1011101111;
   3731: result <= 10'b1011110000;
   3732: result <= 10'b1011110001;
   3733: result <= 10'b1011110001;
   3734: result <= 10'b1011110010;
   3735: result <= 10'b1011110011;
   3736: result <= 10'b1011110011;
   3737: result <= 10'b1011110100;
   3738: result <= 10'b1011110101;
   3739: result <= 10'b1011110101;
   3740: result <= 10'b1011110110;
   3741: result <= 10'b1011110111;
   3742: result <= 10'b1011110111;
   3743: result <= 10'b1011111000;
   3744: result <= 10'b1011111001;
   3745: result <= 10'b1011111001;
   3746: result <= 10'b1011111010;
   3747: result <= 10'b1011111011;
   3748: result <= 10'b1011111011;
   3749: result <= 10'b1011111100;
   3750: result <= 10'b1011111101;
   3751: result <= 10'b1011111110;
   3752: result <= 10'b1011111110;
   3753: result <= 10'b1011111111;
   3754: result <= 10'b1100000000;
   3755: result <= 10'b1100000000;
   3756: result <= 10'b1100000001;
   3757: result <= 10'b1100000010;
   3758: result <= 10'b1100000010;
   3759: result <= 10'b1100000011;
   3760: result <= 10'b1100000100;
   3761: result <= 10'b1100000100;
   3762: result <= 10'b1100000101;
   3763: result <= 10'b1100000110;
   3764: result <= 10'b1100000110;
   3765: result <= 10'b1100000111;
   3766: result <= 10'b1100001000;
   3767: result <= 10'b1100001000;
   3768: result <= 10'b1100001001;
   3769: result <= 10'b1100001010;
   3770: result <= 10'b1100001010;
   3771: result <= 10'b1100001011;
   3772: result <= 10'b1100001100;
   3773: result <= 10'b1100001101;
   3774: result <= 10'b1100001101;
   3775: result <= 10'b1100001110;
   3776: result <= 10'b1100001111;
   3777: result <= 10'b1100001111;
   3778: result <= 10'b1100010000;
   3779: result <= 10'b1100010001;
   3780: result <= 10'b1100010001;
   3781: result <= 10'b1100010010;
   3782: result <= 10'b1100010011;
   3783: result <= 10'b1100010100;
   3784: result <= 10'b1100010100;
   3785: result <= 10'b1100010101;
   3786: result <= 10'b1100010110;
   3787: result <= 10'b1100010110;
   3788: result <= 10'b1100010111;
   3789: result <= 10'b1100011000;
   3790: result <= 10'b1100011000;
   3791: result <= 10'b1100011001;
   3792: result <= 10'b1100011010;
   3793: result <= 10'b1100011011;
   3794: result <= 10'b1100011011;
   3795: result <= 10'b1100011100;
   3796: result <= 10'b1100011101;
   3797: result <= 10'b1100011101;
   3798: result <= 10'b1100011110;
   3799: result <= 10'b1100011111;
   3800: result <= 10'b1100011111;
   3801: result <= 10'b1100100000;
   3802: result <= 10'b1100100001;
   3803: result <= 10'b1100100010;
   3804: result <= 10'b1100100010;
   3805: result <= 10'b1100100011;
   3806: result <= 10'b1100100100;
   3807: result <= 10'b1100100100;
   3808: result <= 10'b1100100101;
   3809: result <= 10'b1100100110;
   3810: result <= 10'b1100100111;
   3811: result <= 10'b1100100111;
   3812: result <= 10'b1100101000;
   3813: result <= 10'b1100101001;
   3814: result <= 10'b1100101001;
   3815: result <= 10'b1100101010;
   3816: result <= 10'b1100101011;
   3817: result <= 10'b1100101100;
   3818: result <= 10'b1100101100;
   3819: result <= 10'b1100101101;
   3820: result <= 10'b1100101110;
   3821: result <= 10'b1100101110;
   3822: result <= 10'b1100101111;
   3823: result <= 10'b1100110000;
   3824: result <= 10'b1100110001;
   3825: result <= 10'b1100110001;
   3826: result <= 10'b1100110010;
   3827: result <= 10'b1100110011;
   3828: result <= 10'b1100110011;
   3829: result <= 10'b1100110100;
   3830: result <= 10'b1100110101;
   3831: result <= 10'b1100110110;
   3832: result <= 10'b1100110110;
   3833: result <= 10'b1100110111;
   3834: result <= 10'b1100111000;
   3835: result <= 10'b1100111000;
   3836: result <= 10'b1100111001;
   3837: result <= 10'b1100111010;
   3838: result <= 10'b1100111011;
   3839: result <= 10'b1100111011;
   3840: result <= 10'b1100111100;
   3841: result <= 10'b1100111101;
   3842: result <= 10'b1100111110;
   3843: result <= 10'b1100111110;
   3844: result <= 10'b1100111111;
   3845: result <= 10'b1101000000;
   3846: result <= 10'b1101000000;
   3847: result <= 10'b1101000001;
   3848: result <= 10'b1101000010;
   3849: result <= 10'b1101000011;
   3850: result <= 10'b1101000011;
   3851: result <= 10'b1101000100;
   3852: result <= 10'b1101000101;
   3853: result <= 10'b1101000110;
   3854: result <= 10'b1101000110;
   3855: result <= 10'b1101000111;
   3856: result <= 10'b1101001000;
   3857: result <= 10'b1101001000;
   3858: result <= 10'b1101001001;
   3859: result <= 10'b1101001010;
   3860: result <= 10'b1101001011;
   3861: result <= 10'b1101001011;
   3862: result <= 10'b1101001100;
   3863: result <= 10'b1101001101;
   3864: result <= 10'b1101001110;
   3865: result <= 10'b1101001110;
   3866: result <= 10'b1101001111;
   3867: result <= 10'b1101010000;
   3868: result <= 10'b1101010001;
   3869: result <= 10'b1101010001;
   3870: result <= 10'b1101010010;
   3871: result <= 10'b1101010011;
   3872: result <= 10'b1101010100;
   3873: result <= 10'b1101010100;
   3874: result <= 10'b1101010101;
   3875: result <= 10'b1101010110;
   3876: result <= 10'b1101010110;
   3877: result <= 10'b1101010111;
   3878: result <= 10'b1101011000;
   3879: result <= 10'b1101011001;
   3880: result <= 10'b1101011001;
   3881: result <= 10'b1101011010;
   3882: result <= 10'b1101011011;
   3883: result <= 10'b1101011100;
   3884: result <= 10'b1101011100;
   3885: result <= 10'b1101011101;
   3886: result <= 10'b1101011110;
   3887: result <= 10'b1101011111;
   3888: result <= 10'b1101011111;
   3889: result <= 10'b1101100000;
   3890: result <= 10'b1101100001;
   3891: result <= 10'b1101100010;
   3892: result <= 10'b1101100010;
   3893: result <= 10'b1101100011;
   3894: result <= 10'b1101100100;
   3895: result <= 10'b1101100101;
   3896: result <= 10'b1101100101;
   3897: result <= 10'b1101100110;
   3898: result <= 10'b1101100111;
   3899: result <= 10'b1101101000;
   3900: result <= 10'b1101101000;
   3901: result <= 10'b1101101001;
   3902: result <= 10'b1101101010;
   3903: result <= 10'b1101101011;
   3904: result <= 10'b1101101011;
   3905: result <= 10'b1101101100;
   3906: result <= 10'b1101101101;
   3907: result <= 10'b1101101110;
   3908: result <= 10'b1101101110;
   3909: result <= 10'b1101101111;
   3910: result <= 10'b1101110000;
   3911: result <= 10'b1101110001;
   3912: result <= 10'b1101110001;
   3913: result <= 10'b1101110010;
   3914: result <= 10'b1101110011;
   3915: result <= 10'b1101110100;
   3916: result <= 10'b1101110100;
   3917: result <= 10'b1101110101;
   3918: result <= 10'b1101110110;
   3919: result <= 10'b1101110111;
   3920: result <= 10'b1101110111;
   3921: result <= 10'b1101111000;
   3922: result <= 10'b1101111001;
   3923: result <= 10'b1101111010;
   3924: result <= 10'b1101111010;
   3925: result <= 10'b1101111011;
   3926: result <= 10'b1101111100;
   3927: result <= 10'b1101111101;
   3928: result <= 10'b1101111110;
   3929: result <= 10'b1101111110;
   3930: result <= 10'b1101111111;
   3931: result <= 10'b1110000000;
   3932: result <= 10'b1110000001;
   3933: result <= 10'b1110000001;
   3934: result <= 10'b1110000010;
   3935: result <= 10'b1110000011;
   3936: result <= 10'b1110000100;
   3937: result <= 10'b1110000100;
   3938: result <= 10'b1110000101;
   3939: result <= 10'b1110000110;
   3940: result <= 10'b1110000111;
   3941: result <= 10'b1110000111;
   3942: result <= 10'b1110001000;
   3943: result <= 10'b1110001001;
   3944: result <= 10'b1110001010;
   3945: result <= 10'b1110001010;
   3946: result <= 10'b1110001011;
   3947: result <= 10'b1110001100;
   3948: result <= 10'b1110001101;
   3949: result <= 10'b1110001110;
   3950: result <= 10'b1110001110;
   3951: result <= 10'b1110001111;
   3952: result <= 10'b1110010000;
   3953: result <= 10'b1110010001;
   3954: result <= 10'b1110010001;
   3955: result <= 10'b1110010010;
   3956: result <= 10'b1110010011;
   3957: result <= 10'b1110010100;
   3958: result <= 10'b1110010100;
   3959: result <= 10'b1110010101;
   3960: result <= 10'b1110010110;
   3961: result <= 10'b1110010111;
   3962: result <= 10'b1110010111;
   3963: result <= 10'b1110011000;
   3964: result <= 10'b1110011001;
   3965: result <= 10'b1110011010;
   3966: result <= 10'b1110011011;
   3967: result <= 10'b1110011011;
   3968: result <= 10'b1110011100;
   3969: result <= 10'b1110011101;
   3970: result <= 10'b1110011110;
   3971: result <= 10'b1110011110;
   3972: result <= 10'b1110011111;
   3973: result <= 10'b1110100000;
   3974: result <= 10'b1110100001;
   3975: result <= 10'b1110100010;
   3976: result <= 10'b1110100010;
   3977: result <= 10'b1110100011;
   3978: result <= 10'b1110100100;
   3979: result <= 10'b1110100101;
   3980: result <= 10'b1110100101;
   3981: result <= 10'b1110100110;
   3982: result <= 10'b1110100111;
   3983: result <= 10'b1110101000;
   3984: result <= 10'b1110101000;
   3985: result <= 10'b1110101001;
   3986: result <= 10'b1110101010;
   3987: result <= 10'b1110101011;
   3988: result <= 10'b1110101100;
   3989: result <= 10'b1110101100;
   3990: result <= 10'b1110101101;
   3991: result <= 10'b1110101110;
   3992: result <= 10'b1110101111;
   3993: result <= 10'b1110101111;
   3994: result <= 10'b1110110000;
   3995: result <= 10'b1110110001;
   3996: result <= 10'b1110110010;
   3997: result <= 10'b1110110011;
   3998: result <= 10'b1110110011;
   3999: result <= 10'b1110110100;
   4000: result <= 10'b1110110101;
   4001: result <= 10'b1110110110;
   4002: result <= 10'b1110110110;
   4003: result <= 10'b1110110111;
   4004: result <= 10'b1110111000;
   4005: result <= 10'b1110111001;
   4006: result <= 10'b1110111010;
   4007: result <= 10'b1110111010;
   4008: result <= 10'b1110111011;
   4009: result <= 10'b1110111100;
   4010: result <= 10'b1110111101;
   4011: result <= 10'b1110111101;
   4012: result <= 10'b1110111110;
   4013: result <= 10'b1110111111;
   4014: result <= 10'b1111000000;
   4015: result <= 10'b1111000001;
   4016: result <= 10'b1111000001;
   4017: result <= 10'b1111000010;
   4018: result <= 10'b1111000011;
   4019: result <= 10'b1111000100;
   4020: result <= 10'b1111000100;
   4021: result <= 10'b1111000101;
   4022: result <= 10'b1111000110;
   4023: result <= 10'b1111000111;
   4024: result <= 10'b1111001000;
   4025: result <= 10'b1111001000;
   4026: result <= 10'b1111001001;
   4027: result <= 10'b1111001010;
   4028: result <= 10'b1111001011;
   4029: result <= 10'b1111001011;
   4030: result <= 10'b1111001100;
   4031: result <= 10'b1111001101;
   4032: result <= 10'b1111001110;
   4033: result <= 10'b1111001111;
   4034: result <= 10'b1111001111;
   4035: result <= 10'b1111010000;
   4036: result <= 10'b1111010001;
   4037: result <= 10'b1111010010;
   4038: result <= 10'b1111010011;
   4039: result <= 10'b1111010011;
   4040: result <= 10'b1111010100;
   4041: result <= 10'b1111010101;
   4042: result <= 10'b1111010110;
   4043: result <= 10'b1111010110;
   4044: result <= 10'b1111010111;
   4045: result <= 10'b1111011000;
   4046: result <= 10'b1111011001;
   4047: result <= 10'b1111011010;
   4048: result <= 10'b1111011010;
   4049: result <= 10'b1111011011;
   4050: result <= 10'b1111011100;
   4051: result <= 10'b1111011101;
   4052: result <= 10'b1111011101;
   4053: result <= 10'b1111011110;
   4054: result <= 10'b1111011111;
   4055: result <= 10'b1111100000;
   4056: result <= 10'b1111100001;
   4057: result <= 10'b1111100001;
   4058: result <= 10'b1111100010;
   4059: result <= 10'b1111100011;
   4060: result <= 10'b1111100100;
   4061: result <= 10'b1111100101;
   4062: result <= 10'b1111100101;
   4063: result <= 10'b1111100110;
   4064: result <= 10'b1111100111;
   4065: result <= 10'b1111101000;
   4066: result <= 10'b1111101000;
   4067: result <= 10'b1111101001;
   4068: result <= 10'b1111101010;
   4069: result <= 10'b1111101011;
   4070: result <= 10'b1111101100;
   4071: result <= 10'b1111101100;
   4072: result <= 10'b1111101101;
   4073: result <= 10'b1111101110;
   4074: result <= 10'b1111101111;
   4075: result <= 10'b1111110000;
   4076: result <= 10'b1111110000;
   4077: result <= 10'b1111110001;
   4078: result <= 10'b1111110010;
   4079: result <= 10'b1111110011;
   4080: result <= 10'b1111110011;
   4081: result <= 10'b1111110100;
   4082: result <= 10'b1111110101;
   4083: result <= 10'b1111110110;
   4084: result <= 10'b1111110111;
   4085: result <= 10'b1111110111;
   4086: result <= 10'b1111111000;
   4087: result <= 10'b1111111001;
   4088: result <= 10'b1111111010;
   4089: result <= 10'b1111111011;
   4090: result <= 10'b1111111011;
   4091: result <= 10'b1111111100;
   4092: result <= 10'b1111111101;
   4093: result <= 10'b1111111110;
   4094: result <= 10'b1111111110;
   4095: result <= 10'b1111111111;
   endcase
endmodule
