`timescale 1ns / 1ps
`default_nettype none


//Created by script createsinelookup.py
module sinetable(input wire [13:0] phase, output reg [11:0] result);

always @(*)
  case(phase)
   0: result <= 12'b000000000000;
   1: result <= 12'b000000000001;
   2: result <= 12'b000000000010;
   3: result <= 12'b000000000010;
   4: result <= 12'b000000000011;
   5: result <= 12'b000000000100;
   6: result <= 12'b000000000101;
   7: result <= 12'b000000000101;
   8: result <= 12'b000000000110;
   9: result <= 12'b000000000111;
   10: result <= 12'b000000001000;
   11: result <= 12'b000000001001;
   12: result <= 12'b000000001001;
   13: result <= 12'b000000001010;
   14: result <= 12'b000000001011;
   15: result <= 12'b000000001100;
   16: result <= 12'b000000001101;
   17: result <= 12'b000000001101;
   18: result <= 12'b000000001110;
   19: result <= 12'b000000001111;
   20: result <= 12'b000000010000;
   21: result <= 12'b000000010000;
   22: result <= 12'b000000010001;
   23: result <= 12'b000000010010;
   24: result <= 12'b000000010011;
   25: result <= 12'b000000010100;
   26: result <= 12'b000000010100;
   27: result <= 12'b000000010101;
   28: result <= 12'b000000010110;
   29: result <= 12'b000000010111;
   30: result <= 12'b000000011000;
   31: result <= 12'b000000011000;
   32: result <= 12'b000000011001;
   33: result <= 12'b000000011010;
   34: result <= 12'b000000011011;
   35: result <= 12'b000000011011;
   36: result <= 12'b000000011100;
   37: result <= 12'b000000011101;
   38: result <= 12'b000000011110;
   39: result <= 12'b000000011111;
   40: result <= 12'b000000011111;
   41: result <= 12'b000000100000;
   42: result <= 12'b000000100001;
   43: result <= 12'b000000100010;
   44: result <= 12'b000000100011;
   45: result <= 12'b000000100011;
   46: result <= 12'b000000100100;
   47: result <= 12'b000000100101;
   48: result <= 12'b000000100110;
   49: result <= 12'b000000100110;
   50: result <= 12'b000000100111;
   51: result <= 12'b000000101000;
   52: result <= 12'b000000101001;
   53: result <= 12'b000000101010;
   54: result <= 12'b000000101010;
   55: result <= 12'b000000101011;
   56: result <= 12'b000000101100;
   57: result <= 12'b000000101101;
   58: result <= 12'b000000101110;
   59: result <= 12'b000000101110;
   60: result <= 12'b000000101111;
   61: result <= 12'b000000110000;
   62: result <= 12'b000000110001;
   63: result <= 12'b000000110001;
   64: result <= 12'b000000110010;
   65: result <= 12'b000000110011;
   66: result <= 12'b000000110100;
   67: result <= 12'b000000110101;
   68: result <= 12'b000000110101;
   69: result <= 12'b000000110110;
   70: result <= 12'b000000110111;
   71: result <= 12'b000000111000;
   72: result <= 12'b000000111001;
   73: result <= 12'b000000111001;
   74: result <= 12'b000000111010;
   75: result <= 12'b000000111011;
   76: result <= 12'b000000111100;
   77: result <= 12'b000000111100;
   78: result <= 12'b000000111101;
   79: result <= 12'b000000111110;
   80: result <= 12'b000000111111;
   81: result <= 12'b000001000000;
   82: result <= 12'b000001000000;
   83: result <= 12'b000001000001;
   84: result <= 12'b000001000010;
   85: result <= 12'b000001000011;
   86: result <= 12'b000001000100;
   87: result <= 12'b000001000100;
   88: result <= 12'b000001000101;
   89: result <= 12'b000001000110;
   90: result <= 12'b000001000111;
   91: result <= 12'b000001000111;
   92: result <= 12'b000001001000;
   93: result <= 12'b000001001001;
   94: result <= 12'b000001001010;
   95: result <= 12'b000001001011;
   96: result <= 12'b000001001011;
   97: result <= 12'b000001001100;
   98: result <= 12'b000001001101;
   99: result <= 12'b000001001110;
   100: result <= 12'b000001001111;
   101: result <= 12'b000001001111;
   102: result <= 12'b000001010000;
   103: result <= 12'b000001010001;
   104: result <= 12'b000001010010;
   105: result <= 12'b000001010010;
   106: result <= 12'b000001010011;
   107: result <= 12'b000001010100;
   108: result <= 12'b000001010101;
   109: result <= 12'b000001010110;
   110: result <= 12'b000001010110;
   111: result <= 12'b000001010111;
   112: result <= 12'b000001011000;
   113: result <= 12'b000001011001;
   114: result <= 12'b000001011010;
   115: result <= 12'b000001011010;
   116: result <= 12'b000001011011;
   117: result <= 12'b000001011100;
   118: result <= 12'b000001011101;
   119: result <= 12'b000001011101;
   120: result <= 12'b000001011110;
   121: result <= 12'b000001011111;
   122: result <= 12'b000001100000;
   123: result <= 12'b000001100001;
   124: result <= 12'b000001100001;
   125: result <= 12'b000001100010;
   126: result <= 12'b000001100011;
   127: result <= 12'b000001100100;
   128: result <= 12'b000001100100;
   129: result <= 12'b000001100101;
   130: result <= 12'b000001100110;
   131: result <= 12'b000001100111;
   132: result <= 12'b000001101000;
   133: result <= 12'b000001101000;
   134: result <= 12'b000001101001;
   135: result <= 12'b000001101010;
   136: result <= 12'b000001101011;
   137: result <= 12'b000001101100;
   138: result <= 12'b000001101100;
   139: result <= 12'b000001101101;
   140: result <= 12'b000001101110;
   141: result <= 12'b000001101111;
   142: result <= 12'b000001101111;
   143: result <= 12'b000001110000;
   144: result <= 12'b000001110001;
   145: result <= 12'b000001110010;
   146: result <= 12'b000001110011;
   147: result <= 12'b000001110011;
   148: result <= 12'b000001110100;
   149: result <= 12'b000001110101;
   150: result <= 12'b000001110110;
   151: result <= 12'b000001110111;
   152: result <= 12'b000001110111;
   153: result <= 12'b000001111000;
   154: result <= 12'b000001111001;
   155: result <= 12'b000001111010;
   156: result <= 12'b000001111010;
   157: result <= 12'b000001111011;
   158: result <= 12'b000001111100;
   159: result <= 12'b000001111101;
   160: result <= 12'b000001111110;
   161: result <= 12'b000001111110;
   162: result <= 12'b000001111111;
   163: result <= 12'b000010000000;
   164: result <= 12'b000010000001;
   165: result <= 12'b000010000010;
   166: result <= 12'b000010000010;
   167: result <= 12'b000010000011;
   168: result <= 12'b000010000100;
   169: result <= 12'b000010000101;
   170: result <= 12'b000010000101;
   171: result <= 12'b000010000110;
   172: result <= 12'b000010000111;
   173: result <= 12'b000010001000;
   174: result <= 12'b000010001001;
   175: result <= 12'b000010001001;
   176: result <= 12'b000010001010;
   177: result <= 12'b000010001011;
   178: result <= 12'b000010001100;
   179: result <= 12'b000010001100;
   180: result <= 12'b000010001101;
   181: result <= 12'b000010001110;
   182: result <= 12'b000010001111;
   183: result <= 12'b000010010000;
   184: result <= 12'b000010010000;
   185: result <= 12'b000010010001;
   186: result <= 12'b000010010010;
   187: result <= 12'b000010010011;
   188: result <= 12'b000010010100;
   189: result <= 12'b000010010100;
   190: result <= 12'b000010010101;
   191: result <= 12'b000010010110;
   192: result <= 12'b000010010111;
   193: result <= 12'b000010010111;
   194: result <= 12'b000010011000;
   195: result <= 12'b000010011001;
   196: result <= 12'b000010011010;
   197: result <= 12'b000010011011;
   198: result <= 12'b000010011011;
   199: result <= 12'b000010011100;
   200: result <= 12'b000010011101;
   201: result <= 12'b000010011110;
   202: result <= 12'b000010011110;
   203: result <= 12'b000010011111;
   204: result <= 12'b000010100000;
   205: result <= 12'b000010100001;
   206: result <= 12'b000010100010;
   207: result <= 12'b000010100010;
   208: result <= 12'b000010100011;
   209: result <= 12'b000010100100;
   210: result <= 12'b000010100101;
   211: result <= 12'b000010100110;
   212: result <= 12'b000010100110;
   213: result <= 12'b000010100111;
   214: result <= 12'b000010101000;
   215: result <= 12'b000010101001;
   216: result <= 12'b000010101001;
   217: result <= 12'b000010101010;
   218: result <= 12'b000010101011;
   219: result <= 12'b000010101100;
   220: result <= 12'b000010101101;
   221: result <= 12'b000010101101;
   222: result <= 12'b000010101110;
   223: result <= 12'b000010101111;
   224: result <= 12'b000010110000;
   225: result <= 12'b000010110000;
   226: result <= 12'b000010110001;
   227: result <= 12'b000010110010;
   228: result <= 12'b000010110011;
   229: result <= 12'b000010110100;
   230: result <= 12'b000010110100;
   231: result <= 12'b000010110101;
   232: result <= 12'b000010110110;
   233: result <= 12'b000010110111;
   234: result <= 12'b000010111000;
   235: result <= 12'b000010111000;
   236: result <= 12'b000010111001;
   237: result <= 12'b000010111010;
   238: result <= 12'b000010111011;
   239: result <= 12'b000010111011;
   240: result <= 12'b000010111100;
   241: result <= 12'b000010111101;
   242: result <= 12'b000010111110;
   243: result <= 12'b000010111111;
   244: result <= 12'b000010111111;
   245: result <= 12'b000011000000;
   246: result <= 12'b000011000001;
   247: result <= 12'b000011000010;
   248: result <= 12'b000011000010;
   249: result <= 12'b000011000011;
   250: result <= 12'b000011000100;
   251: result <= 12'b000011000101;
   252: result <= 12'b000011000110;
   253: result <= 12'b000011000110;
   254: result <= 12'b000011000111;
   255: result <= 12'b000011001000;
   256: result <= 12'b000011001001;
   257: result <= 12'b000011001010;
   258: result <= 12'b000011001010;
   259: result <= 12'b000011001011;
   260: result <= 12'b000011001100;
   261: result <= 12'b000011001101;
   262: result <= 12'b000011001101;
   263: result <= 12'b000011001110;
   264: result <= 12'b000011001111;
   265: result <= 12'b000011010000;
   266: result <= 12'b000011010001;
   267: result <= 12'b000011010001;
   268: result <= 12'b000011010010;
   269: result <= 12'b000011010011;
   270: result <= 12'b000011010100;
   271: result <= 12'b000011010100;
   272: result <= 12'b000011010101;
   273: result <= 12'b000011010110;
   274: result <= 12'b000011010111;
   275: result <= 12'b000011011000;
   276: result <= 12'b000011011000;
   277: result <= 12'b000011011001;
   278: result <= 12'b000011011010;
   279: result <= 12'b000011011011;
   280: result <= 12'b000011011011;
   281: result <= 12'b000011011100;
   282: result <= 12'b000011011101;
   283: result <= 12'b000011011110;
   284: result <= 12'b000011011111;
   285: result <= 12'b000011011111;
   286: result <= 12'b000011100000;
   287: result <= 12'b000011100001;
   288: result <= 12'b000011100010;
   289: result <= 12'b000011100011;
   290: result <= 12'b000011100011;
   291: result <= 12'b000011100100;
   292: result <= 12'b000011100101;
   293: result <= 12'b000011100110;
   294: result <= 12'b000011100110;
   295: result <= 12'b000011100111;
   296: result <= 12'b000011101000;
   297: result <= 12'b000011101001;
   298: result <= 12'b000011101010;
   299: result <= 12'b000011101010;
   300: result <= 12'b000011101011;
   301: result <= 12'b000011101100;
   302: result <= 12'b000011101101;
   303: result <= 12'b000011101101;
   304: result <= 12'b000011101110;
   305: result <= 12'b000011101111;
   306: result <= 12'b000011110000;
   307: result <= 12'b000011110001;
   308: result <= 12'b000011110001;
   309: result <= 12'b000011110010;
   310: result <= 12'b000011110011;
   311: result <= 12'b000011110100;
   312: result <= 12'b000011110100;
   313: result <= 12'b000011110101;
   314: result <= 12'b000011110110;
   315: result <= 12'b000011110111;
   316: result <= 12'b000011111000;
   317: result <= 12'b000011111000;
   318: result <= 12'b000011111001;
   319: result <= 12'b000011111010;
   320: result <= 12'b000011111011;
   321: result <= 12'b000011111011;
   322: result <= 12'b000011111100;
   323: result <= 12'b000011111101;
   324: result <= 12'b000011111110;
   325: result <= 12'b000011111111;
   326: result <= 12'b000011111111;
   327: result <= 12'b000100000000;
   328: result <= 12'b000100000001;
   329: result <= 12'b000100000010;
   330: result <= 12'b000100000010;
   331: result <= 12'b000100000011;
   332: result <= 12'b000100000100;
   333: result <= 12'b000100000101;
   334: result <= 12'b000100000110;
   335: result <= 12'b000100000110;
   336: result <= 12'b000100000111;
   337: result <= 12'b000100001000;
   338: result <= 12'b000100001001;
   339: result <= 12'b000100001010;
   340: result <= 12'b000100001010;
   341: result <= 12'b000100001011;
   342: result <= 12'b000100001100;
   343: result <= 12'b000100001101;
   344: result <= 12'b000100001101;
   345: result <= 12'b000100001110;
   346: result <= 12'b000100001111;
   347: result <= 12'b000100010000;
   348: result <= 12'b000100010001;
   349: result <= 12'b000100010001;
   350: result <= 12'b000100010010;
   351: result <= 12'b000100010011;
   352: result <= 12'b000100010100;
   353: result <= 12'b000100010100;
   354: result <= 12'b000100010101;
   355: result <= 12'b000100010110;
   356: result <= 12'b000100010111;
   357: result <= 12'b000100011000;
   358: result <= 12'b000100011000;
   359: result <= 12'b000100011001;
   360: result <= 12'b000100011010;
   361: result <= 12'b000100011011;
   362: result <= 12'b000100011011;
   363: result <= 12'b000100011100;
   364: result <= 12'b000100011101;
   365: result <= 12'b000100011110;
   366: result <= 12'b000100011111;
   367: result <= 12'b000100011111;
   368: result <= 12'b000100100000;
   369: result <= 12'b000100100001;
   370: result <= 12'b000100100010;
   371: result <= 12'b000100100010;
   372: result <= 12'b000100100011;
   373: result <= 12'b000100100100;
   374: result <= 12'b000100100101;
   375: result <= 12'b000100100110;
   376: result <= 12'b000100100110;
   377: result <= 12'b000100100111;
   378: result <= 12'b000100101000;
   379: result <= 12'b000100101001;
   380: result <= 12'b000100101001;
   381: result <= 12'b000100101010;
   382: result <= 12'b000100101011;
   383: result <= 12'b000100101100;
   384: result <= 12'b000100101101;
   385: result <= 12'b000100101101;
   386: result <= 12'b000100101110;
   387: result <= 12'b000100101111;
   388: result <= 12'b000100110000;
   389: result <= 12'b000100110000;
   390: result <= 12'b000100110001;
   391: result <= 12'b000100110010;
   392: result <= 12'b000100110011;
   393: result <= 12'b000100110011;
   394: result <= 12'b000100110100;
   395: result <= 12'b000100110101;
   396: result <= 12'b000100110110;
   397: result <= 12'b000100110111;
   398: result <= 12'b000100110111;
   399: result <= 12'b000100111000;
   400: result <= 12'b000100111001;
   401: result <= 12'b000100111010;
   402: result <= 12'b000100111010;
   403: result <= 12'b000100111011;
   404: result <= 12'b000100111100;
   405: result <= 12'b000100111101;
   406: result <= 12'b000100111110;
   407: result <= 12'b000100111110;
   408: result <= 12'b000100111111;
   409: result <= 12'b000101000000;
   410: result <= 12'b000101000001;
   411: result <= 12'b000101000001;
   412: result <= 12'b000101000010;
   413: result <= 12'b000101000011;
   414: result <= 12'b000101000100;
   415: result <= 12'b000101000101;
   416: result <= 12'b000101000101;
   417: result <= 12'b000101000110;
   418: result <= 12'b000101000111;
   419: result <= 12'b000101001000;
   420: result <= 12'b000101001000;
   421: result <= 12'b000101001001;
   422: result <= 12'b000101001010;
   423: result <= 12'b000101001011;
   424: result <= 12'b000101001100;
   425: result <= 12'b000101001100;
   426: result <= 12'b000101001101;
   427: result <= 12'b000101001110;
   428: result <= 12'b000101001111;
   429: result <= 12'b000101001111;
   430: result <= 12'b000101010000;
   431: result <= 12'b000101010001;
   432: result <= 12'b000101010010;
   433: result <= 12'b000101010011;
   434: result <= 12'b000101010011;
   435: result <= 12'b000101010100;
   436: result <= 12'b000101010101;
   437: result <= 12'b000101010110;
   438: result <= 12'b000101010110;
   439: result <= 12'b000101010111;
   440: result <= 12'b000101011000;
   441: result <= 12'b000101011001;
   442: result <= 12'b000101011001;
   443: result <= 12'b000101011010;
   444: result <= 12'b000101011011;
   445: result <= 12'b000101011100;
   446: result <= 12'b000101011101;
   447: result <= 12'b000101011101;
   448: result <= 12'b000101011110;
   449: result <= 12'b000101011111;
   450: result <= 12'b000101100000;
   451: result <= 12'b000101100000;
   452: result <= 12'b000101100001;
   453: result <= 12'b000101100010;
   454: result <= 12'b000101100011;
   455: result <= 12'b000101100100;
   456: result <= 12'b000101100100;
   457: result <= 12'b000101100101;
   458: result <= 12'b000101100110;
   459: result <= 12'b000101100111;
   460: result <= 12'b000101100111;
   461: result <= 12'b000101101000;
   462: result <= 12'b000101101001;
   463: result <= 12'b000101101010;
   464: result <= 12'b000101101011;
   465: result <= 12'b000101101011;
   466: result <= 12'b000101101100;
   467: result <= 12'b000101101101;
   468: result <= 12'b000101101110;
   469: result <= 12'b000101101110;
   470: result <= 12'b000101101111;
   471: result <= 12'b000101110000;
   472: result <= 12'b000101110001;
   473: result <= 12'b000101110001;
   474: result <= 12'b000101110010;
   475: result <= 12'b000101110011;
   476: result <= 12'b000101110100;
   477: result <= 12'b000101110101;
   478: result <= 12'b000101110101;
   479: result <= 12'b000101110110;
   480: result <= 12'b000101110111;
   481: result <= 12'b000101111000;
   482: result <= 12'b000101111000;
   483: result <= 12'b000101111001;
   484: result <= 12'b000101111010;
   485: result <= 12'b000101111011;
   486: result <= 12'b000101111011;
   487: result <= 12'b000101111100;
   488: result <= 12'b000101111101;
   489: result <= 12'b000101111110;
   490: result <= 12'b000101111111;
   491: result <= 12'b000101111111;
   492: result <= 12'b000110000000;
   493: result <= 12'b000110000001;
   494: result <= 12'b000110000010;
   495: result <= 12'b000110000010;
   496: result <= 12'b000110000011;
   497: result <= 12'b000110000100;
   498: result <= 12'b000110000101;
   499: result <= 12'b000110000110;
   500: result <= 12'b000110000110;
   501: result <= 12'b000110000111;
   502: result <= 12'b000110001000;
   503: result <= 12'b000110001001;
   504: result <= 12'b000110001001;
   505: result <= 12'b000110001010;
   506: result <= 12'b000110001011;
   507: result <= 12'b000110001100;
   508: result <= 12'b000110001100;
   509: result <= 12'b000110001101;
   510: result <= 12'b000110001110;
   511: result <= 12'b000110001111;
   512: result <= 12'b000110010000;
   513: result <= 12'b000110010000;
   514: result <= 12'b000110010001;
   515: result <= 12'b000110010010;
   516: result <= 12'b000110010011;
   517: result <= 12'b000110010011;
   518: result <= 12'b000110010100;
   519: result <= 12'b000110010101;
   520: result <= 12'b000110010110;
   521: result <= 12'b000110010110;
   522: result <= 12'b000110010111;
   523: result <= 12'b000110011000;
   524: result <= 12'b000110011001;
   525: result <= 12'b000110011010;
   526: result <= 12'b000110011010;
   527: result <= 12'b000110011011;
   528: result <= 12'b000110011100;
   529: result <= 12'b000110011101;
   530: result <= 12'b000110011101;
   531: result <= 12'b000110011110;
   532: result <= 12'b000110011111;
   533: result <= 12'b000110100000;
   534: result <= 12'b000110100000;
   535: result <= 12'b000110100001;
   536: result <= 12'b000110100010;
   537: result <= 12'b000110100011;
   538: result <= 12'b000110100100;
   539: result <= 12'b000110100100;
   540: result <= 12'b000110100101;
   541: result <= 12'b000110100110;
   542: result <= 12'b000110100111;
   543: result <= 12'b000110100111;
   544: result <= 12'b000110101000;
   545: result <= 12'b000110101001;
   546: result <= 12'b000110101010;
   547: result <= 12'b000110101010;
   548: result <= 12'b000110101011;
   549: result <= 12'b000110101100;
   550: result <= 12'b000110101101;
   551: result <= 12'b000110101110;
   552: result <= 12'b000110101110;
   553: result <= 12'b000110101111;
   554: result <= 12'b000110110000;
   555: result <= 12'b000110110001;
   556: result <= 12'b000110110001;
   557: result <= 12'b000110110010;
   558: result <= 12'b000110110011;
   559: result <= 12'b000110110100;
   560: result <= 12'b000110110100;
   561: result <= 12'b000110110101;
   562: result <= 12'b000110110110;
   563: result <= 12'b000110110111;
   564: result <= 12'b000110111000;
   565: result <= 12'b000110111000;
   566: result <= 12'b000110111001;
   567: result <= 12'b000110111010;
   568: result <= 12'b000110111011;
   569: result <= 12'b000110111011;
   570: result <= 12'b000110111100;
   571: result <= 12'b000110111101;
   572: result <= 12'b000110111110;
   573: result <= 12'b000110111110;
   574: result <= 12'b000110111111;
   575: result <= 12'b000111000000;
   576: result <= 12'b000111000001;
   577: result <= 12'b000111000001;
   578: result <= 12'b000111000010;
   579: result <= 12'b000111000011;
   580: result <= 12'b000111000100;
   581: result <= 12'b000111000101;
   582: result <= 12'b000111000101;
   583: result <= 12'b000111000110;
   584: result <= 12'b000111000111;
   585: result <= 12'b000111001000;
   586: result <= 12'b000111001000;
   587: result <= 12'b000111001001;
   588: result <= 12'b000111001010;
   589: result <= 12'b000111001011;
   590: result <= 12'b000111001011;
   591: result <= 12'b000111001100;
   592: result <= 12'b000111001101;
   593: result <= 12'b000111001110;
   594: result <= 12'b000111001111;
   595: result <= 12'b000111001111;
   596: result <= 12'b000111010000;
   597: result <= 12'b000111010001;
   598: result <= 12'b000111010010;
   599: result <= 12'b000111010010;
   600: result <= 12'b000111010011;
   601: result <= 12'b000111010100;
   602: result <= 12'b000111010101;
   603: result <= 12'b000111010101;
   604: result <= 12'b000111010110;
   605: result <= 12'b000111010111;
   606: result <= 12'b000111011000;
   607: result <= 12'b000111011000;
   608: result <= 12'b000111011001;
   609: result <= 12'b000111011010;
   610: result <= 12'b000111011011;
   611: result <= 12'b000111011011;
   612: result <= 12'b000111011100;
   613: result <= 12'b000111011101;
   614: result <= 12'b000111011110;
   615: result <= 12'b000111011111;
   616: result <= 12'b000111011111;
   617: result <= 12'b000111100000;
   618: result <= 12'b000111100001;
   619: result <= 12'b000111100010;
   620: result <= 12'b000111100010;
   621: result <= 12'b000111100011;
   622: result <= 12'b000111100100;
   623: result <= 12'b000111100101;
   624: result <= 12'b000111100101;
   625: result <= 12'b000111100110;
   626: result <= 12'b000111100111;
   627: result <= 12'b000111101000;
   628: result <= 12'b000111101000;
   629: result <= 12'b000111101001;
   630: result <= 12'b000111101010;
   631: result <= 12'b000111101011;
   632: result <= 12'b000111101100;
   633: result <= 12'b000111101100;
   634: result <= 12'b000111101101;
   635: result <= 12'b000111101110;
   636: result <= 12'b000111101111;
   637: result <= 12'b000111101111;
   638: result <= 12'b000111110000;
   639: result <= 12'b000111110001;
   640: result <= 12'b000111110010;
   641: result <= 12'b000111110010;
   642: result <= 12'b000111110011;
   643: result <= 12'b000111110100;
   644: result <= 12'b000111110101;
   645: result <= 12'b000111110101;
   646: result <= 12'b000111110110;
   647: result <= 12'b000111110111;
   648: result <= 12'b000111111000;
   649: result <= 12'b000111111000;
   650: result <= 12'b000111111001;
   651: result <= 12'b000111111010;
   652: result <= 12'b000111111011;
   653: result <= 12'b000111111100;
   654: result <= 12'b000111111100;
   655: result <= 12'b000111111101;
   656: result <= 12'b000111111110;
   657: result <= 12'b000111111111;
   658: result <= 12'b000111111111;
   659: result <= 12'b001000000000;
   660: result <= 12'b001000000001;
   661: result <= 12'b001000000010;
   662: result <= 12'b001000000010;
   663: result <= 12'b001000000011;
   664: result <= 12'b001000000100;
   665: result <= 12'b001000000101;
   666: result <= 12'b001000000101;
   667: result <= 12'b001000000110;
   668: result <= 12'b001000000111;
   669: result <= 12'b001000001000;
   670: result <= 12'b001000001000;
   671: result <= 12'b001000001001;
   672: result <= 12'b001000001010;
   673: result <= 12'b001000001011;
   674: result <= 12'b001000001011;
   675: result <= 12'b001000001100;
   676: result <= 12'b001000001101;
   677: result <= 12'b001000001110;
   678: result <= 12'b001000001111;
   679: result <= 12'b001000001111;
   680: result <= 12'b001000010000;
   681: result <= 12'b001000010001;
   682: result <= 12'b001000010010;
   683: result <= 12'b001000010010;
   684: result <= 12'b001000010011;
   685: result <= 12'b001000010100;
   686: result <= 12'b001000010101;
   687: result <= 12'b001000010101;
   688: result <= 12'b001000010110;
   689: result <= 12'b001000010111;
   690: result <= 12'b001000011000;
   691: result <= 12'b001000011000;
   692: result <= 12'b001000011001;
   693: result <= 12'b001000011010;
   694: result <= 12'b001000011011;
   695: result <= 12'b001000011011;
   696: result <= 12'b001000011100;
   697: result <= 12'b001000011101;
   698: result <= 12'b001000011110;
   699: result <= 12'b001000011110;
   700: result <= 12'b001000011111;
   701: result <= 12'b001000100000;
   702: result <= 12'b001000100001;
   703: result <= 12'b001000100001;
   704: result <= 12'b001000100010;
   705: result <= 12'b001000100011;
   706: result <= 12'b001000100100;
   707: result <= 12'b001000100100;
   708: result <= 12'b001000100101;
   709: result <= 12'b001000100110;
   710: result <= 12'b001000100111;
   711: result <= 12'b001000101000;
   712: result <= 12'b001000101000;
   713: result <= 12'b001000101001;
   714: result <= 12'b001000101010;
   715: result <= 12'b001000101011;
   716: result <= 12'b001000101011;
   717: result <= 12'b001000101100;
   718: result <= 12'b001000101101;
   719: result <= 12'b001000101110;
   720: result <= 12'b001000101110;
   721: result <= 12'b001000101111;
   722: result <= 12'b001000110000;
   723: result <= 12'b001000110001;
   724: result <= 12'b001000110001;
   725: result <= 12'b001000110010;
   726: result <= 12'b001000110011;
   727: result <= 12'b001000110100;
   728: result <= 12'b001000110100;
   729: result <= 12'b001000110101;
   730: result <= 12'b001000110110;
   731: result <= 12'b001000110111;
   732: result <= 12'b001000110111;
   733: result <= 12'b001000111000;
   734: result <= 12'b001000111001;
   735: result <= 12'b001000111010;
   736: result <= 12'b001000111010;
   737: result <= 12'b001000111011;
   738: result <= 12'b001000111100;
   739: result <= 12'b001000111101;
   740: result <= 12'b001000111101;
   741: result <= 12'b001000111110;
   742: result <= 12'b001000111111;
   743: result <= 12'b001001000000;
   744: result <= 12'b001001000000;
   745: result <= 12'b001001000001;
   746: result <= 12'b001001000010;
   747: result <= 12'b001001000011;
   748: result <= 12'b001001000011;
   749: result <= 12'b001001000100;
   750: result <= 12'b001001000101;
   751: result <= 12'b001001000110;
   752: result <= 12'b001001000110;
   753: result <= 12'b001001000111;
   754: result <= 12'b001001001000;
   755: result <= 12'b001001001001;
   756: result <= 12'b001001001001;
   757: result <= 12'b001001001010;
   758: result <= 12'b001001001011;
   759: result <= 12'b001001001100;
   760: result <= 12'b001001001100;
   761: result <= 12'b001001001101;
   762: result <= 12'b001001001110;
   763: result <= 12'b001001001111;
   764: result <= 12'b001001001111;
   765: result <= 12'b001001010000;
   766: result <= 12'b001001010001;
   767: result <= 12'b001001010010;
   768: result <= 12'b001001010011;
   769: result <= 12'b001001010011;
   770: result <= 12'b001001010100;
   771: result <= 12'b001001010101;
   772: result <= 12'b001001010110;
   773: result <= 12'b001001010110;
   774: result <= 12'b001001010111;
   775: result <= 12'b001001011000;
   776: result <= 12'b001001011001;
   777: result <= 12'b001001011001;
   778: result <= 12'b001001011010;
   779: result <= 12'b001001011011;
   780: result <= 12'b001001011100;
   781: result <= 12'b001001011100;
   782: result <= 12'b001001011101;
   783: result <= 12'b001001011110;
   784: result <= 12'b001001011111;
   785: result <= 12'b001001011111;
   786: result <= 12'b001001100000;
   787: result <= 12'b001001100001;
   788: result <= 12'b001001100010;
   789: result <= 12'b001001100010;
   790: result <= 12'b001001100011;
   791: result <= 12'b001001100100;
   792: result <= 12'b001001100101;
   793: result <= 12'b001001100101;
   794: result <= 12'b001001100110;
   795: result <= 12'b001001100111;
   796: result <= 12'b001001101000;
   797: result <= 12'b001001101000;
   798: result <= 12'b001001101001;
   799: result <= 12'b001001101010;
   800: result <= 12'b001001101011;
   801: result <= 12'b001001101011;
   802: result <= 12'b001001101100;
   803: result <= 12'b001001101101;
   804: result <= 12'b001001101110;
   805: result <= 12'b001001101110;
   806: result <= 12'b001001101111;
   807: result <= 12'b001001110000;
   808: result <= 12'b001001110000;
   809: result <= 12'b001001110001;
   810: result <= 12'b001001110010;
   811: result <= 12'b001001110011;
   812: result <= 12'b001001110011;
   813: result <= 12'b001001110100;
   814: result <= 12'b001001110101;
   815: result <= 12'b001001110110;
   816: result <= 12'b001001110110;
   817: result <= 12'b001001110111;
   818: result <= 12'b001001111000;
   819: result <= 12'b001001111001;
   820: result <= 12'b001001111001;
   821: result <= 12'b001001111010;
   822: result <= 12'b001001111011;
   823: result <= 12'b001001111100;
   824: result <= 12'b001001111100;
   825: result <= 12'b001001111101;
   826: result <= 12'b001001111110;
   827: result <= 12'b001001111111;
   828: result <= 12'b001001111111;
   829: result <= 12'b001010000000;
   830: result <= 12'b001010000001;
   831: result <= 12'b001010000010;
   832: result <= 12'b001010000010;
   833: result <= 12'b001010000011;
   834: result <= 12'b001010000100;
   835: result <= 12'b001010000101;
   836: result <= 12'b001010000101;
   837: result <= 12'b001010000110;
   838: result <= 12'b001010000111;
   839: result <= 12'b001010001000;
   840: result <= 12'b001010001000;
   841: result <= 12'b001010001001;
   842: result <= 12'b001010001010;
   843: result <= 12'b001010001011;
   844: result <= 12'b001010001011;
   845: result <= 12'b001010001100;
   846: result <= 12'b001010001101;
   847: result <= 12'b001010001110;
   848: result <= 12'b001010001110;
   849: result <= 12'b001010001111;
   850: result <= 12'b001010010000;
   851: result <= 12'b001010010001;
   852: result <= 12'b001010010001;
   853: result <= 12'b001010010010;
   854: result <= 12'b001010010011;
   855: result <= 12'b001010010100;
   856: result <= 12'b001010010100;
   857: result <= 12'b001010010101;
   858: result <= 12'b001010010110;
   859: result <= 12'b001010010111;
   860: result <= 12'b001010010111;
   861: result <= 12'b001010011000;
   862: result <= 12'b001010011001;
   863: result <= 12'b001010011001;
   864: result <= 12'b001010011010;
   865: result <= 12'b001010011011;
   866: result <= 12'b001010011100;
   867: result <= 12'b001010011100;
   868: result <= 12'b001010011101;
   869: result <= 12'b001010011110;
   870: result <= 12'b001010011111;
   871: result <= 12'b001010011111;
   872: result <= 12'b001010100000;
   873: result <= 12'b001010100001;
   874: result <= 12'b001010100010;
   875: result <= 12'b001010100010;
   876: result <= 12'b001010100011;
   877: result <= 12'b001010100100;
   878: result <= 12'b001010100101;
   879: result <= 12'b001010100101;
   880: result <= 12'b001010100110;
   881: result <= 12'b001010100111;
   882: result <= 12'b001010101000;
   883: result <= 12'b001010101000;
   884: result <= 12'b001010101001;
   885: result <= 12'b001010101010;
   886: result <= 12'b001010101011;
   887: result <= 12'b001010101011;
   888: result <= 12'b001010101100;
   889: result <= 12'b001010101101;
   890: result <= 12'b001010101110;
   891: result <= 12'b001010101110;
   892: result <= 12'b001010101111;
   893: result <= 12'b001010110000;
   894: result <= 12'b001010110000;
   895: result <= 12'b001010110001;
   896: result <= 12'b001010110010;
   897: result <= 12'b001010110011;
   898: result <= 12'b001010110011;
   899: result <= 12'b001010110100;
   900: result <= 12'b001010110101;
   901: result <= 12'b001010110110;
   902: result <= 12'b001010110110;
   903: result <= 12'b001010110111;
   904: result <= 12'b001010111000;
   905: result <= 12'b001010111001;
   906: result <= 12'b001010111001;
   907: result <= 12'b001010111010;
   908: result <= 12'b001010111011;
   909: result <= 12'b001010111100;
   910: result <= 12'b001010111100;
   911: result <= 12'b001010111101;
   912: result <= 12'b001010111110;
   913: result <= 12'b001010111111;
   914: result <= 12'b001010111111;
   915: result <= 12'b001011000000;
   916: result <= 12'b001011000001;
   917: result <= 12'b001011000001;
   918: result <= 12'b001011000010;
   919: result <= 12'b001011000011;
   920: result <= 12'b001011000100;
   921: result <= 12'b001011000100;
   922: result <= 12'b001011000101;
   923: result <= 12'b001011000110;
   924: result <= 12'b001011000111;
   925: result <= 12'b001011000111;
   926: result <= 12'b001011001000;
   927: result <= 12'b001011001001;
   928: result <= 12'b001011001010;
   929: result <= 12'b001011001010;
   930: result <= 12'b001011001011;
   931: result <= 12'b001011001100;
   932: result <= 12'b001011001101;
   933: result <= 12'b001011001101;
   934: result <= 12'b001011001110;
   935: result <= 12'b001011001111;
   936: result <= 12'b001011001111;
   937: result <= 12'b001011010000;
   938: result <= 12'b001011010001;
   939: result <= 12'b001011010010;
   940: result <= 12'b001011010010;
   941: result <= 12'b001011010011;
   942: result <= 12'b001011010100;
   943: result <= 12'b001011010101;
   944: result <= 12'b001011010101;
   945: result <= 12'b001011010110;
   946: result <= 12'b001011010111;
   947: result <= 12'b001011011000;
   948: result <= 12'b001011011000;
   949: result <= 12'b001011011001;
   950: result <= 12'b001011011010;
   951: result <= 12'b001011011010;
   952: result <= 12'b001011011011;
   953: result <= 12'b001011011100;
   954: result <= 12'b001011011101;
   955: result <= 12'b001011011101;
   956: result <= 12'b001011011110;
   957: result <= 12'b001011011111;
   958: result <= 12'b001011100000;
   959: result <= 12'b001011100000;
   960: result <= 12'b001011100001;
   961: result <= 12'b001011100010;
   962: result <= 12'b001011100011;
   963: result <= 12'b001011100011;
   964: result <= 12'b001011100100;
   965: result <= 12'b001011100101;
   966: result <= 12'b001011100101;
   967: result <= 12'b001011100110;
   968: result <= 12'b001011100111;
   969: result <= 12'b001011101000;
   970: result <= 12'b001011101000;
   971: result <= 12'b001011101001;
   972: result <= 12'b001011101010;
   973: result <= 12'b001011101011;
   974: result <= 12'b001011101011;
   975: result <= 12'b001011101100;
   976: result <= 12'b001011101101;
   977: result <= 12'b001011101110;
   978: result <= 12'b001011101110;
   979: result <= 12'b001011101111;
   980: result <= 12'b001011110000;
   981: result <= 12'b001011110000;
   982: result <= 12'b001011110001;
   983: result <= 12'b001011110010;
   984: result <= 12'b001011110011;
   985: result <= 12'b001011110011;
   986: result <= 12'b001011110100;
   987: result <= 12'b001011110101;
   988: result <= 12'b001011110110;
   989: result <= 12'b001011110110;
   990: result <= 12'b001011110111;
   991: result <= 12'b001011111000;
   992: result <= 12'b001011111000;
   993: result <= 12'b001011111001;
   994: result <= 12'b001011111010;
   995: result <= 12'b001011111011;
   996: result <= 12'b001011111011;
   997: result <= 12'b001011111100;
   998: result <= 12'b001011111101;
   999: result <= 12'b001011111110;
   1000: result <= 12'b001011111110;
   1001: result <= 12'b001011111111;
   1002: result <= 12'b001100000000;
   1003: result <= 12'b001100000000;
   1004: result <= 12'b001100000001;
   1005: result <= 12'b001100000010;
   1006: result <= 12'b001100000011;
   1007: result <= 12'b001100000011;
   1008: result <= 12'b001100000100;
   1009: result <= 12'b001100000101;
   1010: result <= 12'b001100000110;
   1011: result <= 12'b001100000110;
   1012: result <= 12'b001100000111;
   1013: result <= 12'b001100001000;
   1014: result <= 12'b001100001000;
   1015: result <= 12'b001100001001;
   1016: result <= 12'b001100001010;
   1017: result <= 12'b001100001011;
   1018: result <= 12'b001100001011;
   1019: result <= 12'b001100001100;
   1020: result <= 12'b001100001101;
   1021: result <= 12'b001100001110;
   1022: result <= 12'b001100001110;
   1023: result <= 12'b001100001111;
   1024: result <= 12'b001100010000;
   1025: result <= 12'b001100010000;
   1026: result <= 12'b001100010001;
   1027: result <= 12'b001100010010;
   1028: result <= 12'b001100010011;
   1029: result <= 12'b001100010011;
   1030: result <= 12'b001100010100;
   1031: result <= 12'b001100010101;
   1032: result <= 12'b001100010110;
   1033: result <= 12'b001100010110;
   1034: result <= 12'b001100010111;
   1035: result <= 12'b001100011000;
   1036: result <= 12'b001100011000;
   1037: result <= 12'b001100011001;
   1038: result <= 12'b001100011010;
   1039: result <= 12'b001100011011;
   1040: result <= 12'b001100011011;
   1041: result <= 12'b001100011100;
   1042: result <= 12'b001100011101;
   1043: result <= 12'b001100011110;
   1044: result <= 12'b001100011110;
   1045: result <= 12'b001100011111;
   1046: result <= 12'b001100100000;
   1047: result <= 12'b001100100000;
   1048: result <= 12'b001100100001;
   1049: result <= 12'b001100100010;
   1050: result <= 12'b001100100011;
   1051: result <= 12'b001100100011;
   1052: result <= 12'b001100100100;
   1053: result <= 12'b001100100101;
   1054: result <= 12'b001100100101;
   1055: result <= 12'b001100100110;
   1056: result <= 12'b001100100111;
   1057: result <= 12'b001100101000;
   1058: result <= 12'b001100101000;
   1059: result <= 12'b001100101001;
   1060: result <= 12'b001100101010;
   1061: result <= 12'b001100101011;
   1062: result <= 12'b001100101011;
   1063: result <= 12'b001100101100;
   1064: result <= 12'b001100101101;
   1065: result <= 12'b001100101101;
   1066: result <= 12'b001100101110;
   1067: result <= 12'b001100101111;
   1068: result <= 12'b001100110000;
   1069: result <= 12'b001100110000;
   1070: result <= 12'b001100110001;
   1071: result <= 12'b001100110010;
   1072: result <= 12'b001100110010;
   1073: result <= 12'b001100110011;
   1074: result <= 12'b001100110100;
   1075: result <= 12'b001100110101;
   1076: result <= 12'b001100110101;
   1077: result <= 12'b001100110110;
   1078: result <= 12'b001100110111;
   1079: result <= 12'b001100110111;
   1080: result <= 12'b001100111000;
   1081: result <= 12'b001100111001;
   1082: result <= 12'b001100111010;
   1083: result <= 12'b001100111010;
   1084: result <= 12'b001100111011;
   1085: result <= 12'b001100111100;
   1086: result <= 12'b001100111100;
   1087: result <= 12'b001100111101;
   1088: result <= 12'b001100111110;
   1089: result <= 12'b001100111111;
   1090: result <= 12'b001100111111;
   1091: result <= 12'b001101000000;
   1092: result <= 12'b001101000001;
   1093: result <= 12'b001101000010;
   1094: result <= 12'b001101000010;
   1095: result <= 12'b001101000011;
   1096: result <= 12'b001101000100;
   1097: result <= 12'b001101000100;
   1098: result <= 12'b001101000101;
   1099: result <= 12'b001101000110;
   1100: result <= 12'b001101000111;
   1101: result <= 12'b001101000111;
   1102: result <= 12'b001101001000;
   1103: result <= 12'b001101001001;
   1104: result <= 12'b001101001001;
   1105: result <= 12'b001101001010;
   1106: result <= 12'b001101001011;
   1107: result <= 12'b001101001100;
   1108: result <= 12'b001101001100;
   1109: result <= 12'b001101001101;
   1110: result <= 12'b001101001110;
   1111: result <= 12'b001101001110;
   1112: result <= 12'b001101001111;
   1113: result <= 12'b001101010000;
   1114: result <= 12'b001101010001;
   1115: result <= 12'b001101010001;
   1116: result <= 12'b001101010010;
   1117: result <= 12'b001101010011;
   1118: result <= 12'b001101010011;
   1119: result <= 12'b001101010100;
   1120: result <= 12'b001101010101;
   1121: result <= 12'b001101010110;
   1122: result <= 12'b001101010110;
   1123: result <= 12'b001101010111;
   1124: result <= 12'b001101011000;
   1125: result <= 12'b001101011000;
   1126: result <= 12'b001101011001;
   1127: result <= 12'b001101011010;
   1128: result <= 12'b001101011011;
   1129: result <= 12'b001101011011;
   1130: result <= 12'b001101011100;
   1131: result <= 12'b001101011101;
   1132: result <= 12'b001101011101;
   1133: result <= 12'b001101011110;
   1134: result <= 12'b001101011111;
   1135: result <= 12'b001101100000;
   1136: result <= 12'b001101100000;
   1137: result <= 12'b001101100001;
   1138: result <= 12'b001101100010;
   1139: result <= 12'b001101100010;
   1140: result <= 12'b001101100011;
   1141: result <= 12'b001101100100;
   1142: result <= 12'b001101100101;
   1143: result <= 12'b001101100101;
   1144: result <= 12'b001101100110;
   1145: result <= 12'b001101100111;
   1146: result <= 12'b001101100111;
   1147: result <= 12'b001101101000;
   1148: result <= 12'b001101101001;
   1149: result <= 12'b001101101010;
   1150: result <= 12'b001101101010;
   1151: result <= 12'b001101101011;
   1152: result <= 12'b001101101100;
   1153: result <= 12'b001101101100;
   1154: result <= 12'b001101101101;
   1155: result <= 12'b001101101110;
   1156: result <= 12'b001101101110;
   1157: result <= 12'b001101101111;
   1158: result <= 12'b001101110000;
   1159: result <= 12'b001101110001;
   1160: result <= 12'b001101110001;
   1161: result <= 12'b001101110010;
   1162: result <= 12'b001101110011;
   1163: result <= 12'b001101110011;
   1164: result <= 12'b001101110100;
   1165: result <= 12'b001101110101;
   1166: result <= 12'b001101110110;
   1167: result <= 12'b001101110110;
   1168: result <= 12'b001101110111;
   1169: result <= 12'b001101111000;
   1170: result <= 12'b001101111000;
   1171: result <= 12'b001101111001;
   1172: result <= 12'b001101111010;
   1173: result <= 12'b001101111011;
   1174: result <= 12'b001101111011;
   1175: result <= 12'b001101111100;
   1176: result <= 12'b001101111101;
   1177: result <= 12'b001101111101;
   1178: result <= 12'b001101111110;
   1179: result <= 12'b001101111111;
   1180: result <= 12'b001101111111;
   1181: result <= 12'b001110000000;
   1182: result <= 12'b001110000001;
   1183: result <= 12'b001110000010;
   1184: result <= 12'b001110000010;
   1185: result <= 12'b001110000011;
   1186: result <= 12'b001110000100;
   1187: result <= 12'b001110000100;
   1188: result <= 12'b001110000101;
   1189: result <= 12'b001110000110;
   1190: result <= 12'b001110000111;
   1191: result <= 12'b001110000111;
   1192: result <= 12'b001110001000;
   1193: result <= 12'b001110001001;
   1194: result <= 12'b001110001001;
   1195: result <= 12'b001110001010;
   1196: result <= 12'b001110001011;
   1197: result <= 12'b001110001011;
   1198: result <= 12'b001110001100;
   1199: result <= 12'b001110001101;
   1200: result <= 12'b001110001110;
   1201: result <= 12'b001110001110;
   1202: result <= 12'b001110001111;
   1203: result <= 12'b001110010000;
   1204: result <= 12'b001110010000;
   1205: result <= 12'b001110010001;
   1206: result <= 12'b001110010010;
   1207: result <= 12'b001110010010;
   1208: result <= 12'b001110010011;
   1209: result <= 12'b001110010100;
   1210: result <= 12'b001110010101;
   1211: result <= 12'b001110010101;
   1212: result <= 12'b001110010110;
   1213: result <= 12'b001110010111;
   1214: result <= 12'b001110010111;
   1215: result <= 12'b001110011000;
   1216: result <= 12'b001110011001;
   1217: result <= 12'b001110011010;
   1218: result <= 12'b001110011010;
   1219: result <= 12'b001110011011;
   1220: result <= 12'b001110011100;
   1221: result <= 12'b001110011100;
   1222: result <= 12'b001110011101;
   1223: result <= 12'b001110011110;
   1224: result <= 12'b001110011110;
   1225: result <= 12'b001110011111;
   1226: result <= 12'b001110100000;
   1227: result <= 12'b001110100001;
   1228: result <= 12'b001110100001;
   1229: result <= 12'b001110100010;
   1230: result <= 12'b001110100011;
   1231: result <= 12'b001110100011;
   1232: result <= 12'b001110100100;
   1233: result <= 12'b001110100101;
   1234: result <= 12'b001110100101;
   1235: result <= 12'b001110100110;
   1236: result <= 12'b001110100111;
   1237: result <= 12'b001110101000;
   1238: result <= 12'b001110101000;
   1239: result <= 12'b001110101001;
   1240: result <= 12'b001110101010;
   1241: result <= 12'b001110101010;
   1242: result <= 12'b001110101011;
   1243: result <= 12'b001110101100;
   1244: result <= 12'b001110101100;
   1245: result <= 12'b001110101101;
   1246: result <= 12'b001110101110;
   1247: result <= 12'b001110101110;
   1248: result <= 12'b001110101111;
   1249: result <= 12'b001110110000;
   1250: result <= 12'b001110110001;
   1251: result <= 12'b001110110001;
   1252: result <= 12'b001110110010;
   1253: result <= 12'b001110110011;
   1254: result <= 12'b001110110011;
   1255: result <= 12'b001110110100;
   1256: result <= 12'b001110110101;
   1257: result <= 12'b001110110101;
   1258: result <= 12'b001110110110;
   1259: result <= 12'b001110110111;
   1260: result <= 12'b001110111000;
   1261: result <= 12'b001110111000;
   1262: result <= 12'b001110111001;
   1263: result <= 12'b001110111010;
   1264: result <= 12'b001110111010;
   1265: result <= 12'b001110111011;
   1266: result <= 12'b001110111100;
   1267: result <= 12'b001110111100;
   1268: result <= 12'b001110111101;
   1269: result <= 12'b001110111110;
   1270: result <= 12'b001110111110;
   1271: result <= 12'b001110111111;
   1272: result <= 12'b001111000000;
   1273: result <= 12'b001111000001;
   1274: result <= 12'b001111000001;
   1275: result <= 12'b001111000010;
   1276: result <= 12'b001111000011;
   1277: result <= 12'b001111000011;
   1278: result <= 12'b001111000100;
   1279: result <= 12'b001111000101;
   1280: result <= 12'b001111000101;
   1281: result <= 12'b001111000110;
   1282: result <= 12'b001111000111;
   1283: result <= 12'b001111000111;
   1284: result <= 12'b001111001000;
   1285: result <= 12'b001111001001;
   1286: result <= 12'b001111001010;
   1287: result <= 12'b001111001010;
   1288: result <= 12'b001111001011;
   1289: result <= 12'b001111001100;
   1290: result <= 12'b001111001100;
   1291: result <= 12'b001111001101;
   1292: result <= 12'b001111001110;
   1293: result <= 12'b001111001110;
   1294: result <= 12'b001111001111;
   1295: result <= 12'b001111010000;
   1296: result <= 12'b001111010000;
   1297: result <= 12'b001111010001;
   1298: result <= 12'b001111010010;
   1299: result <= 12'b001111010011;
   1300: result <= 12'b001111010011;
   1301: result <= 12'b001111010100;
   1302: result <= 12'b001111010101;
   1303: result <= 12'b001111010101;
   1304: result <= 12'b001111010110;
   1305: result <= 12'b001111010111;
   1306: result <= 12'b001111010111;
   1307: result <= 12'b001111011000;
   1308: result <= 12'b001111011001;
   1309: result <= 12'b001111011001;
   1310: result <= 12'b001111011010;
   1311: result <= 12'b001111011011;
   1312: result <= 12'b001111011100;
   1313: result <= 12'b001111011100;
   1314: result <= 12'b001111011101;
   1315: result <= 12'b001111011110;
   1316: result <= 12'b001111011110;
   1317: result <= 12'b001111011111;
   1318: result <= 12'b001111100000;
   1319: result <= 12'b001111100000;
   1320: result <= 12'b001111100001;
   1321: result <= 12'b001111100010;
   1322: result <= 12'b001111100010;
   1323: result <= 12'b001111100011;
   1324: result <= 12'b001111100100;
   1325: result <= 12'b001111100100;
   1326: result <= 12'b001111100101;
   1327: result <= 12'b001111100110;
   1328: result <= 12'b001111100111;
   1329: result <= 12'b001111100111;
   1330: result <= 12'b001111101000;
   1331: result <= 12'b001111101001;
   1332: result <= 12'b001111101001;
   1333: result <= 12'b001111101010;
   1334: result <= 12'b001111101011;
   1335: result <= 12'b001111101011;
   1336: result <= 12'b001111101100;
   1337: result <= 12'b001111101101;
   1338: result <= 12'b001111101101;
   1339: result <= 12'b001111101110;
   1340: result <= 12'b001111101111;
   1341: result <= 12'b001111101111;
   1342: result <= 12'b001111110000;
   1343: result <= 12'b001111110001;
   1344: result <= 12'b001111110001;
   1345: result <= 12'b001111110010;
   1346: result <= 12'b001111110011;
   1347: result <= 12'b001111110100;
   1348: result <= 12'b001111110100;
   1349: result <= 12'b001111110101;
   1350: result <= 12'b001111110110;
   1351: result <= 12'b001111110110;
   1352: result <= 12'b001111110111;
   1353: result <= 12'b001111111000;
   1354: result <= 12'b001111111000;
   1355: result <= 12'b001111111001;
   1356: result <= 12'b001111111010;
   1357: result <= 12'b001111111010;
   1358: result <= 12'b001111111011;
   1359: result <= 12'b001111111100;
   1360: result <= 12'b001111111100;
   1361: result <= 12'b001111111101;
   1362: result <= 12'b001111111110;
   1363: result <= 12'b001111111110;
   1364: result <= 12'b001111111111;
   1365: result <= 12'b010000000000;
   1366: result <= 12'b010000000000;
   1367: result <= 12'b010000000001;
   1368: result <= 12'b010000000010;
   1369: result <= 12'b010000000010;
   1370: result <= 12'b010000000011;
   1371: result <= 12'b010000000100;
   1372: result <= 12'b010000000101;
   1373: result <= 12'b010000000101;
   1374: result <= 12'b010000000110;
   1375: result <= 12'b010000000111;
   1376: result <= 12'b010000000111;
   1377: result <= 12'b010000001000;
   1378: result <= 12'b010000001001;
   1379: result <= 12'b010000001001;
   1380: result <= 12'b010000001010;
   1381: result <= 12'b010000001011;
   1382: result <= 12'b010000001011;
   1383: result <= 12'b010000001100;
   1384: result <= 12'b010000001101;
   1385: result <= 12'b010000001101;
   1386: result <= 12'b010000001110;
   1387: result <= 12'b010000001111;
   1388: result <= 12'b010000001111;
   1389: result <= 12'b010000010000;
   1390: result <= 12'b010000010001;
   1391: result <= 12'b010000010001;
   1392: result <= 12'b010000010010;
   1393: result <= 12'b010000010011;
   1394: result <= 12'b010000010011;
   1395: result <= 12'b010000010100;
   1396: result <= 12'b010000010101;
   1397: result <= 12'b010000010101;
   1398: result <= 12'b010000010110;
   1399: result <= 12'b010000010111;
   1400: result <= 12'b010000010111;
   1401: result <= 12'b010000011000;
   1402: result <= 12'b010000011001;
   1403: result <= 12'b010000011010;
   1404: result <= 12'b010000011010;
   1405: result <= 12'b010000011011;
   1406: result <= 12'b010000011100;
   1407: result <= 12'b010000011100;
   1408: result <= 12'b010000011101;
   1409: result <= 12'b010000011110;
   1410: result <= 12'b010000011110;
   1411: result <= 12'b010000011111;
   1412: result <= 12'b010000100000;
   1413: result <= 12'b010000100000;
   1414: result <= 12'b010000100001;
   1415: result <= 12'b010000100010;
   1416: result <= 12'b010000100010;
   1417: result <= 12'b010000100011;
   1418: result <= 12'b010000100100;
   1419: result <= 12'b010000100100;
   1420: result <= 12'b010000100101;
   1421: result <= 12'b010000100110;
   1422: result <= 12'b010000100110;
   1423: result <= 12'b010000100111;
   1424: result <= 12'b010000101000;
   1425: result <= 12'b010000101000;
   1426: result <= 12'b010000101001;
   1427: result <= 12'b010000101010;
   1428: result <= 12'b010000101010;
   1429: result <= 12'b010000101011;
   1430: result <= 12'b010000101100;
   1431: result <= 12'b010000101100;
   1432: result <= 12'b010000101101;
   1433: result <= 12'b010000101110;
   1434: result <= 12'b010000101110;
   1435: result <= 12'b010000101111;
   1436: result <= 12'b010000110000;
   1437: result <= 12'b010000110000;
   1438: result <= 12'b010000110001;
   1439: result <= 12'b010000110010;
   1440: result <= 12'b010000110010;
   1441: result <= 12'b010000110011;
   1442: result <= 12'b010000110100;
   1443: result <= 12'b010000110100;
   1444: result <= 12'b010000110101;
   1445: result <= 12'b010000110110;
   1446: result <= 12'b010000110110;
   1447: result <= 12'b010000110111;
   1448: result <= 12'b010000111000;
   1449: result <= 12'b010000111000;
   1450: result <= 12'b010000111001;
   1451: result <= 12'b010000111010;
   1452: result <= 12'b010000111010;
   1453: result <= 12'b010000111011;
   1454: result <= 12'b010000111100;
   1455: result <= 12'b010000111100;
   1456: result <= 12'b010000111101;
   1457: result <= 12'b010000111110;
   1458: result <= 12'b010000111110;
   1459: result <= 12'b010000111111;
   1460: result <= 12'b010001000000;
   1461: result <= 12'b010001000000;
   1462: result <= 12'b010001000001;
   1463: result <= 12'b010001000010;
   1464: result <= 12'b010001000010;
   1465: result <= 12'b010001000011;
   1466: result <= 12'b010001000100;
   1467: result <= 12'b010001000100;
   1468: result <= 12'b010001000101;
   1469: result <= 12'b010001000110;
   1470: result <= 12'b010001000110;
   1471: result <= 12'b010001000111;
   1472: result <= 12'b010001001000;
   1473: result <= 12'b010001001000;
   1474: result <= 12'b010001001001;
   1475: result <= 12'b010001001010;
   1476: result <= 12'b010001001010;
   1477: result <= 12'b010001001011;
   1478: result <= 12'b010001001100;
   1479: result <= 12'b010001001100;
   1480: result <= 12'b010001001101;
   1481: result <= 12'b010001001110;
   1482: result <= 12'b010001001110;
   1483: result <= 12'b010001001111;
   1484: result <= 12'b010001010000;
   1485: result <= 12'b010001010000;
   1486: result <= 12'b010001010001;
   1487: result <= 12'b010001010010;
   1488: result <= 12'b010001010010;
   1489: result <= 12'b010001010011;
   1490: result <= 12'b010001010100;
   1491: result <= 12'b010001010100;
   1492: result <= 12'b010001010101;
   1493: result <= 12'b010001010110;
   1494: result <= 12'b010001010110;
   1495: result <= 12'b010001010111;
   1496: result <= 12'b010001011000;
   1497: result <= 12'b010001011000;
   1498: result <= 12'b010001011001;
   1499: result <= 12'b010001011010;
   1500: result <= 12'b010001011010;
   1501: result <= 12'b010001011011;
   1502: result <= 12'b010001011100;
   1503: result <= 12'b010001011100;
   1504: result <= 12'b010001011101;
   1505: result <= 12'b010001011101;
   1506: result <= 12'b010001011110;
   1507: result <= 12'b010001011111;
   1508: result <= 12'b010001011111;
   1509: result <= 12'b010001100000;
   1510: result <= 12'b010001100001;
   1511: result <= 12'b010001100001;
   1512: result <= 12'b010001100010;
   1513: result <= 12'b010001100011;
   1514: result <= 12'b010001100011;
   1515: result <= 12'b010001100100;
   1516: result <= 12'b010001100101;
   1517: result <= 12'b010001100101;
   1518: result <= 12'b010001100110;
   1519: result <= 12'b010001100111;
   1520: result <= 12'b010001100111;
   1521: result <= 12'b010001101000;
   1522: result <= 12'b010001101001;
   1523: result <= 12'b010001101001;
   1524: result <= 12'b010001101010;
   1525: result <= 12'b010001101011;
   1526: result <= 12'b010001101011;
   1527: result <= 12'b010001101100;
   1528: result <= 12'b010001101101;
   1529: result <= 12'b010001101101;
   1530: result <= 12'b010001101110;
   1531: result <= 12'b010001101111;
   1532: result <= 12'b010001101111;
   1533: result <= 12'b010001110000;
   1534: result <= 12'b010001110001;
   1535: result <= 12'b010001110001;
   1536: result <= 12'b010001110010;
   1537: result <= 12'b010001110010;
   1538: result <= 12'b010001110011;
   1539: result <= 12'b010001110100;
   1540: result <= 12'b010001110100;
   1541: result <= 12'b010001110101;
   1542: result <= 12'b010001110110;
   1543: result <= 12'b010001110110;
   1544: result <= 12'b010001110111;
   1545: result <= 12'b010001111000;
   1546: result <= 12'b010001111000;
   1547: result <= 12'b010001111001;
   1548: result <= 12'b010001111010;
   1549: result <= 12'b010001111010;
   1550: result <= 12'b010001111011;
   1551: result <= 12'b010001111100;
   1552: result <= 12'b010001111100;
   1553: result <= 12'b010001111101;
   1554: result <= 12'b010001111110;
   1555: result <= 12'b010001111110;
   1556: result <= 12'b010001111111;
   1557: result <= 12'b010001111111;
   1558: result <= 12'b010010000000;
   1559: result <= 12'b010010000001;
   1560: result <= 12'b010010000001;
   1561: result <= 12'b010010000010;
   1562: result <= 12'b010010000011;
   1563: result <= 12'b010010000011;
   1564: result <= 12'b010010000100;
   1565: result <= 12'b010010000101;
   1566: result <= 12'b010010000101;
   1567: result <= 12'b010010000110;
   1568: result <= 12'b010010000111;
   1569: result <= 12'b010010000111;
   1570: result <= 12'b010010001000;
   1571: result <= 12'b010010001001;
   1572: result <= 12'b010010001001;
   1573: result <= 12'b010010001010;
   1574: result <= 12'b010010001011;
   1575: result <= 12'b010010001011;
   1576: result <= 12'b010010001100;
   1577: result <= 12'b010010001100;
   1578: result <= 12'b010010001101;
   1579: result <= 12'b010010001110;
   1580: result <= 12'b010010001110;
   1581: result <= 12'b010010001111;
   1582: result <= 12'b010010010000;
   1583: result <= 12'b010010010000;
   1584: result <= 12'b010010010001;
   1585: result <= 12'b010010010010;
   1586: result <= 12'b010010010010;
   1587: result <= 12'b010010010011;
   1588: result <= 12'b010010010100;
   1589: result <= 12'b010010010100;
   1590: result <= 12'b010010010101;
   1591: result <= 12'b010010010101;
   1592: result <= 12'b010010010110;
   1593: result <= 12'b010010010111;
   1594: result <= 12'b010010010111;
   1595: result <= 12'b010010011000;
   1596: result <= 12'b010010011001;
   1597: result <= 12'b010010011001;
   1598: result <= 12'b010010011010;
   1599: result <= 12'b010010011011;
   1600: result <= 12'b010010011011;
   1601: result <= 12'b010010011100;
   1602: result <= 12'b010010011101;
   1603: result <= 12'b010010011101;
   1604: result <= 12'b010010011110;
   1605: result <= 12'b010010011110;
   1606: result <= 12'b010010011111;
   1607: result <= 12'b010010100000;
   1608: result <= 12'b010010100000;
   1609: result <= 12'b010010100001;
   1610: result <= 12'b010010100010;
   1611: result <= 12'b010010100010;
   1612: result <= 12'b010010100011;
   1613: result <= 12'b010010100100;
   1614: result <= 12'b010010100100;
   1615: result <= 12'b010010100101;
   1616: result <= 12'b010010100110;
   1617: result <= 12'b010010100110;
   1618: result <= 12'b010010100111;
   1619: result <= 12'b010010100111;
   1620: result <= 12'b010010101000;
   1621: result <= 12'b010010101001;
   1622: result <= 12'b010010101001;
   1623: result <= 12'b010010101010;
   1624: result <= 12'b010010101011;
   1625: result <= 12'b010010101011;
   1626: result <= 12'b010010101100;
   1627: result <= 12'b010010101101;
   1628: result <= 12'b010010101101;
   1629: result <= 12'b010010101110;
   1630: result <= 12'b010010101110;
   1631: result <= 12'b010010101111;
   1632: result <= 12'b010010110000;
   1633: result <= 12'b010010110000;
   1634: result <= 12'b010010110001;
   1635: result <= 12'b010010110010;
   1636: result <= 12'b010010110010;
   1637: result <= 12'b010010110011;
   1638: result <= 12'b010010110100;
   1639: result <= 12'b010010110100;
   1640: result <= 12'b010010110101;
   1641: result <= 12'b010010110101;
   1642: result <= 12'b010010110110;
   1643: result <= 12'b010010110111;
   1644: result <= 12'b010010110111;
   1645: result <= 12'b010010111000;
   1646: result <= 12'b010010111001;
   1647: result <= 12'b010010111001;
   1648: result <= 12'b010010111010;
   1649: result <= 12'b010010111011;
   1650: result <= 12'b010010111011;
   1651: result <= 12'b010010111100;
   1652: result <= 12'b010010111100;
   1653: result <= 12'b010010111101;
   1654: result <= 12'b010010111110;
   1655: result <= 12'b010010111110;
   1656: result <= 12'b010010111111;
   1657: result <= 12'b010011000000;
   1658: result <= 12'b010011000000;
   1659: result <= 12'b010011000001;
   1660: result <= 12'b010011000001;
   1661: result <= 12'b010011000010;
   1662: result <= 12'b010011000011;
   1663: result <= 12'b010011000011;
   1664: result <= 12'b010011000100;
   1665: result <= 12'b010011000101;
   1666: result <= 12'b010011000101;
   1667: result <= 12'b010011000110;
   1668: result <= 12'b010011000111;
   1669: result <= 12'b010011000111;
   1670: result <= 12'b010011001000;
   1671: result <= 12'b010011001000;
   1672: result <= 12'b010011001001;
   1673: result <= 12'b010011001010;
   1674: result <= 12'b010011001010;
   1675: result <= 12'b010011001011;
   1676: result <= 12'b010011001100;
   1677: result <= 12'b010011001100;
   1678: result <= 12'b010011001101;
   1679: result <= 12'b010011001101;
   1680: result <= 12'b010011001110;
   1681: result <= 12'b010011001111;
   1682: result <= 12'b010011001111;
   1683: result <= 12'b010011010000;
   1684: result <= 12'b010011010001;
   1685: result <= 12'b010011010001;
   1686: result <= 12'b010011010010;
   1687: result <= 12'b010011010010;
   1688: result <= 12'b010011010011;
   1689: result <= 12'b010011010100;
   1690: result <= 12'b010011010100;
   1691: result <= 12'b010011010101;
   1692: result <= 12'b010011010110;
   1693: result <= 12'b010011010110;
   1694: result <= 12'b010011010111;
   1695: result <= 12'b010011010111;
   1696: result <= 12'b010011011000;
   1697: result <= 12'b010011011001;
   1698: result <= 12'b010011011001;
   1699: result <= 12'b010011011010;
   1700: result <= 12'b010011011011;
   1701: result <= 12'b010011011011;
   1702: result <= 12'b010011011100;
   1703: result <= 12'b010011011100;
   1704: result <= 12'b010011011101;
   1705: result <= 12'b010011011110;
   1706: result <= 12'b010011011110;
   1707: result <= 12'b010011011111;
   1708: result <= 12'b010011100000;
   1709: result <= 12'b010011100000;
   1710: result <= 12'b010011100001;
   1711: result <= 12'b010011100001;
   1712: result <= 12'b010011100010;
   1713: result <= 12'b010011100011;
   1714: result <= 12'b010011100011;
   1715: result <= 12'b010011100100;
   1716: result <= 12'b010011100101;
   1717: result <= 12'b010011100101;
   1718: result <= 12'b010011100110;
   1719: result <= 12'b010011100110;
   1720: result <= 12'b010011100111;
   1721: result <= 12'b010011101000;
   1722: result <= 12'b010011101000;
   1723: result <= 12'b010011101001;
   1724: result <= 12'b010011101010;
   1725: result <= 12'b010011101010;
   1726: result <= 12'b010011101011;
   1727: result <= 12'b010011101011;
   1728: result <= 12'b010011101100;
   1729: result <= 12'b010011101101;
   1730: result <= 12'b010011101101;
   1731: result <= 12'b010011101110;
   1732: result <= 12'b010011101110;
   1733: result <= 12'b010011101111;
   1734: result <= 12'b010011110000;
   1735: result <= 12'b010011110000;
   1736: result <= 12'b010011110001;
   1737: result <= 12'b010011110010;
   1738: result <= 12'b010011110010;
   1739: result <= 12'b010011110011;
   1740: result <= 12'b010011110011;
   1741: result <= 12'b010011110100;
   1742: result <= 12'b010011110101;
   1743: result <= 12'b010011110101;
   1744: result <= 12'b010011110110;
   1745: result <= 12'b010011110110;
   1746: result <= 12'b010011110111;
   1747: result <= 12'b010011111000;
   1748: result <= 12'b010011111000;
   1749: result <= 12'b010011111001;
   1750: result <= 12'b010011111010;
   1751: result <= 12'b010011111010;
   1752: result <= 12'b010011111011;
   1753: result <= 12'b010011111011;
   1754: result <= 12'b010011111100;
   1755: result <= 12'b010011111101;
   1756: result <= 12'b010011111101;
   1757: result <= 12'b010011111110;
   1758: result <= 12'b010011111110;
   1759: result <= 12'b010011111111;
   1760: result <= 12'b010100000000;
   1761: result <= 12'b010100000000;
   1762: result <= 12'b010100000001;
   1763: result <= 12'b010100000010;
   1764: result <= 12'b010100000010;
   1765: result <= 12'b010100000011;
   1766: result <= 12'b010100000011;
   1767: result <= 12'b010100000100;
   1768: result <= 12'b010100000101;
   1769: result <= 12'b010100000101;
   1770: result <= 12'b010100000110;
   1771: result <= 12'b010100000110;
   1772: result <= 12'b010100000111;
   1773: result <= 12'b010100001000;
   1774: result <= 12'b010100001000;
   1775: result <= 12'b010100001001;
   1776: result <= 12'b010100001001;
   1777: result <= 12'b010100001010;
   1778: result <= 12'b010100001011;
   1779: result <= 12'b010100001011;
   1780: result <= 12'b010100001100;
   1781: result <= 12'b010100001101;
   1782: result <= 12'b010100001101;
   1783: result <= 12'b010100001110;
   1784: result <= 12'b010100001110;
   1785: result <= 12'b010100001111;
   1786: result <= 12'b010100010000;
   1787: result <= 12'b010100010000;
   1788: result <= 12'b010100010001;
   1789: result <= 12'b010100010001;
   1790: result <= 12'b010100010010;
   1791: result <= 12'b010100010011;
   1792: result <= 12'b010100010011;
   1793: result <= 12'b010100010100;
   1794: result <= 12'b010100010100;
   1795: result <= 12'b010100010101;
   1796: result <= 12'b010100010110;
   1797: result <= 12'b010100010110;
   1798: result <= 12'b010100010111;
   1799: result <= 12'b010100010111;
   1800: result <= 12'b010100011000;
   1801: result <= 12'b010100011001;
   1802: result <= 12'b010100011001;
   1803: result <= 12'b010100011010;
   1804: result <= 12'b010100011011;
   1805: result <= 12'b010100011011;
   1806: result <= 12'b010100011100;
   1807: result <= 12'b010100011100;
   1808: result <= 12'b010100011101;
   1809: result <= 12'b010100011110;
   1810: result <= 12'b010100011110;
   1811: result <= 12'b010100011111;
   1812: result <= 12'b010100011111;
   1813: result <= 12'b010100100000;
   1814: result <= 12'b010100100001;
   1815: result <= 12'b010100100001;
   1816: result <= 12'b010100100010;
   1817: result <= 12'b010100100010;
   1818: result <= 12'b010100100011;
   1819: result <= 12'b010100100100;
   1820: result <= 12'b010100100100;
   1821: result <= 12'b010100100101;
   1822: result <= 12'b010100100101;
   1823: result <= 12'b010100100110;
   1824: result <= 12'b010100100111;
   1825: result <= 12'b010100100111;
   1826: result <= 12'b010100101000;
   1827: result <= 12'b010100101000;
   1828: result <= 12'b010100101001;
   1829: result <= 12'b010100101010;
   1830: result <= 12'b010100101010;
   1831: result <= 12'b010100101011;
   1832: result <= 12'b010100101011;
   1833: result <= 12'b010100101100;
   1834: result <= 12'b010100101101;
   1835: result <= 12'b010100101101;
   1836: result <= 12'b010100101110;
   1837: result <= 12'b010100101110;
   1838: result <= 12'b010100101111;
   1839: result <= 12'b010100110000;
   1840: result <= 12'b010100110000;
   1841: result <= 12'b010100110001;
   1842: result <= 12'b010100110001;
   1843: result <= 12'b010100110010;
   1844: result <= 12'b010100110011;
   1845: result <= 12'b010100110011;
   1846: result <= 12'b010100110100;
   1847: result <= 12'b010100110100;
   1848: result <= 12'b010100110101;
   1849: result <= 12'b010100110110;
   1850: result <= 12'b010100110110;
   1851: result <= 12'b010100110111;
   1852: result <= 12'b010100110111;
   1853: result <= 12'b010100111000;
   1854: result <= 12'b010100111001;
   1855: result <= 12'b010100111001;
   1856: result <= 12'b010100111010;
   1857: result <= 12'b010100111010;
   1858: result <= 12'b010100111011;
   1859: result <= 12'b010100111011;
   1860: result <= 12'b010100111100;
   1861: result <= 12'b010100111101;
   1862: result <= 12'b010100111101;
   1863: result <= 12'b010100111110;
   1864: result <= 12'b010100111110;
   1865: result <= 12'b010100111111;
   1866: result <= 12'b010101000000;
   1867: result <= 12'b010101000000;
   1868: result <= 12'b010101000001;
   1869: result <= 12'b010101000001;
   1870: result <= 12'b010101000010;
   1871: result <= 12'b010101000011;
   1872: result <= 12'b010101000011;
   1873: result <= 12'b010101000100;
   1874: result <= 12'b010101000100;
   1875: result <= 12'b010101000101;
   1876: result <= 12'b010101000110;
   1877: result <= 12'b010101000110;
   1878: result <= 12'b010101000111;
   1879: result <= 12'b010101000111;
   1880: result <= 12'b010101001000;
   1881: result <= 12'b010101001001;
   1882: result <= 12'b010101001001;
   1883: result <= 12'b010101001010;
   1884: result <= 12'b010101001010;
   1885: result <= 12'b010101001011;
   1886: result <= 12'b010101001011;
   1887: result <= 12'b010101001100;
   1888: result <= 12'b010101001101;
   1889: result <= 12'b010101001101;
   1890: result <= 12'b010101001110;
   1891: result <= 12'b010101001110;
   1892: result <= 12'b010101001111;
   1893: result <= 12'b010101010000;
   1894: result <= 12'b010101010000;
   1895: result <= 12'b010101010001;
   1896: result <= 12'b010101010001;
   1897: result <= 12'b010101010010;
   1898: result <= 12'b010101010011;
   1899: result <= 12'b010101010011;
   1900: result <= 12'b010101010100;
   1901: result <= 12'b010101010100;
   1902: result <= 12'b010101010101;
   1903: result <= 12'b010101010101;
   1904: result <= 12'b010101010110;
   1905: result <= 12'b010101010111;
   1906: result <= 12'b010101010111;
   1907: result <= 12'b010101011000;
   1908: result <= 12'b010101011000;
   1909: result <= 12'b010101011001;
   1910: result <= 12'b010101011010;
   1911: result <= 12'b010101011010;
   1912: result <= 12'b010101011011;
   1913: result <= 12'b010101011011;
   1914: result <= 12'b010101011100;
   1915: result <= 12'b010101011100;
   1916: result <= 12'b010101011101;
   1917: result <= 12'b010101011110;
   1918: result <= 12'b010101011110;
   1919: result <= 12'b010101011111;
   1920: result <= 12'b010101011111;
   1921: result <= 12'b010101100000;
   1922: result <= 12'b010101100001;
   1923: result <= 12'b010101100001;
   1924: result <= 12'b010101100010;
   1925: result <= 12'b010101100010;
   1926: result <= 12'b010101100011;
   1927: result <= 12'b010101100011;
   1928: result <= 12'b010101100100;
   1929: result <= 12'b010101100101;
   1930: result <= 12'b010101100101;
   1931: result <= 12'b010101100110;
   1932: result <= 12'b010101100110;
   1933: result <= 12'b010101100111;
   1934: result <= 12'b010101100111;
   1935: result <= 12'b010101101000;
   1936: result <= 12'b010101101001;
   1937: result <= 12'b010101101001;
   1938: result <= 12'b010101101010;
   1939: result <= 12'b010101101010;
   1940: result <= 12'b010101101011;
   1941: result <= 12'b010101101100;
   1942: result <= 12'b010101101100;
   1943: result <= 12'b010101101101;
   1944: result <= 12'b010101101101;
   1945: result <= 12'b010101101110;
   1946: result <= 12'b010101101110;
   1947: result <= 12'b010101101111;
   1948: result <= 12'b010101110000;
   1949: result <= 12'b010101110000;
   1950: result <= 12'b010101110001;
   1951: result <= 12'b010101110001;
   1952: result <= 12'b010101110010;
   1953: result <= 12'b010101110010;
   1954: result <= 12'b010101110011;
   1955: result <= 12'b010101110100;
   1956: result <= 12'b010101110100;
   1957: result <= 12'b010101110101;
   1958: result <= 12'b010101110101;
   1959: result <= 12'b010101110110;
   1960: result <= 12'b010101110110;
   1961: result <= 12'b010101110111;
   1962: result <= 12'b010101111000;
   1963: result <= 12'b010101111000;
   1964: result <= 12'b010101111001;
   1965: result <= 12'b010101111001;
   1966: result <= 12'b010101111010;
   1967: result <= 12'b010101111010;
   1968: result <= 12'b010101111011;
   1969: result <= 12'b010101111100;
   1970: result <= 12'b010101111100;
   1971: result <= 12'b010101111101;
   1972: result <= 12'b010101111101;
   1973: result <= 12'b010101111110;
   1974: result <= 12'b010101111110;
   1975: result <= 12'b010101111111;
   1976: result <= 12'b010110000000;
   1977: result <= 12'b010110000000;
   1978: result <= 12'b010110000001;
   1979: result <= 12'b010110000001;
   1980: result <= 12'b010110000010;
   1981: result <= 12'b010110000010;
   1982: result <= 12'b010110000011;
   1983: result <= 12'b010110000100;
   1984: result <= 12'b010110000100;
   1985: result <= 12'b010110000101;
   1986: result <= 12'b010110000101;
   1987: result <= 12'b010110000110;
   1988: result <= 12'b010110000110;
   1989: result <= 12'b010110000111;
   1990: result <= 12'b010110001000;
   1991: result <= 12'b010110001000;
   1992: result <= 12'b010110001001;
   1993: result <= 12'b010110001001;
   1994: result <= 12'b010110001010;
   1995: result <= 12'b010110001010;
   1996: result <= 12'b010110001011;
   1997: result <= 12'b010110001100;
   1998: result <= 12'b010110001100;
   1999: result <= 12'b010110001101;
   2000: result <= 12'b010110001101;
   2001: result <= 12'b010110001110;
   2002: result <= 12'b010110001110;
   2003: result <= 12'b010110001111;
   2004: result <= 12'b010110010000;
   2005: result <= 12'b010110010000;
   2006: result <= 12'b010110010001;
   2007: result <= 12'b010110010001;
   2008: result <= 12'b010110010010;
   2009: result <= 12'b010110010010;
   2010: result <= 12'b010110010011;
   2011: result <= 12'b010110010011;
   2012: result <= 12'b010110010100;
   2013: result <= 12'b010110010101;
   2014: result <= 12'b010110010101;
   2015: result <= 12'b010110010110;
   2016: result <= 12'b010110010110;
   2017: result <= 12'b010110010111;
   2018: result <= 12'b010110010111;
   2019: result <= 12'b010110011000;
   2020: result <= 12'b010110011001;
   2021: result <= 12'b010110011001;
   2022: result <= 12'b010110011010;
   2023: result <= 12'b010110011010;
   2024: result <= 12'b010110011011;
   2025: result <= 12'b010110011011;
   2026: result <= 12'b010110011100;
   2027: result <= 12'b010110011100;
   2028: result <= 12'b010110011101;
   2029: result <= 12'b010110011110;
   2030: result <= 12'b010110011110;
   2031: result <= 12'b010110011111;
   2032: result <= 12'b010110011111;
   2033: result <= 12'b010110100000;
   2034: result <= 12'b010110100000;
   2035: result <= 12'b010110100001;
   2036: result <= 12'b010110100001;
   2037: result <= 12'b010110100010;
   2038: result <= 12'b010110100011;
   2039: result <= 12'b010110100011;
   2040: result <= 12'b010110100100;
   2041: result <= 12'b010110100100;
   2042: result <= 12'b010110100101;
   2043: result <= 12'b010110100101;
   2044: result <= 12'b010110100110;
   2045: result <= 12'b010110100110;
   2046: result <= 12'b010110100111;
   2047: result <= 12'b010110101000;
   2048: result <= 12'b010110101000;
   2049: result <= 12'b010110101001;
   2050: result <= 12'b010110101001;
   2051: result <= 12'b010110101010;
   2052: result <= 12'b010110101010;
   2053: result <= 12'b010110101011;
   2054: result <= 12'b010110101011;
   2055: result <= 12'b010110101100;
   2056: result <= 12'b010110101101;
   2057: result <= 12'b010110101101;
   2058: result <= 12'b010110101110;
   2059: result <= 12'b010110101110;
   2060: result <= 12'b010110101111;
   2061: result <= 12'b010110101111;
   2062: result <= 12'b010110110000;
   2063: result <= 12'b010110110000;
   2064: result <= 12'b010110110001;
   2065: result <= 12'b010110110010;
   2066: result <= 12'b010110110010;
   2067: result <= 12'b010110110011;
   2068: result <= 12'b010110110011;
   2069: result <= 12'b010110110100;
   2070: result <= 12'b010110110100;
   2071: result <= 12'b010110110101;
   2072: result <= 12'b010110110101;
   2073: result <= 12'b010110110110;
   2074: result <= 12'b010110110111;
   2075: result <= 12'b010110110111;
   2076: result <= 12'b010110111000;
   2077: result <= 12'b010110111000;
   2078: result <= 12'b010110111001;
   2079: result <= 12'b010110111001;
   2080: result <= 12'b010110111010;
   2081: result <= 12'b010110111010;
   2082: result <= 12'b010110111011;
   2083: result <= 12'b010110111011;
   2084: result <= 12'b010110111100;
   2085: result <= 12'b010110111101;
   2086: result <= 12'b010110111101;
   2087: result <= 12'b010110111110;
   2088: result <= 12'b010110111110;
   2089: result <= 12'b010110111111;
   2090: result <= 12'b010110111111;
   2091: result <= 12'b010111000000;
   2092: result <= 12'b010111000000;
   2093: result <= 12'b010111000001;
   2094: result <= 12'b010111000001;
   2095: result <= 12'b010111000010;
   2096: result <= 12'b010111000011;
   2097: result <= 12'b010111000011;
   2098: result <= 12'b010111000100;
   2099: result <= 12'b010111000100;
   2100: result <= 12'b010111000101;
   2101: result <= 12'b010111000101;
   2102: result <= 12'b010111000110;
   2103: result <= 12'b010111000110;
   2104: result <= 12'b010111000111;
   2105: result <= 12'b010111000111;
   2106: result <= 12'b010111001000;
   2107: result <= 12'b010111001001;
   2108: result <= 12'b010111001001;
   2109: result <= 12'b010111001010;
   2110: result <= 12'b010111001010;
   2111: result <= 12'b010111001011;
   2112: result <= 12'b010111001011;
   2113: result <= 12'b010111001100;
   2114: result <= 12'b010111001100;
   2115: result <= 12'b010111001101;
   2116: result <= 12'b010111001101;
   2117: result <= 12'b010111001110;
   2118: result <= 12'b010111001111;
   2119: result <= 12'b010111001111;
   2120: result <= 12'b010111010000;
   2121: result <= 12'b010111010000;
   2122: result <= 12'b010111010001;
   2123: result <= 12'b010111010001;
   2124: result <= 12'b010111010010;
   2125: result <= 12'b010111010010;
   2126: result <= 12'b010111010011;
   2127: result <= 12'b010111010011;
   2128: result <= 12'b010111010100;
   2129: result <= 12'b010111010100;
   2130: result <= 12'b010111010101;
   2131: result <= 12'b010111010110;
   2132: result <= 12'b010111010110;
   2133: result <= 12'b010111010111;
   2134: result <= 12'b010111010111;
   2135: result <= 12'b010111011000;
   2136: result <= 12'b010111011000;
   2137: result <= 12'b010111011001;
   2138: result <= 12'b010111011001;
   2139: result <= 12'b010111011010;
   2140: result <= 12'b010111011010;
   2141: result <= 12'b010111011011;
   2142: result <= 12'b010111011011;
   2143: result <= 12'b010111011100;
   2144: result <= 12'b010111011100;
   2145: result <= 12'b010111011101;
   2146: result <= 12'b010111011110;
   2147: result <= 12'b010111011110;
   2148: result <= 12'b010111011111;
   2149: result <= 12'b010111011111;
   2150: result <= 12'b010111100000;
   2151: result <= 12'b010111100000;
   2152: result <= 12'b010111100001;
   2153: result <= 12'b010111100001;
   2154: result <= 12'b010111100010;
   2155: result <= 12'b010111100010;
   2156: result <= 12'b010111100011;
   2157: result <= 12'b010111100011;
   2158: result <= 12'b010111100100;
   2159: result <= 12'b010111100100;
   2160: result <= 12'b010111100101;
   2161: result <= 12'b010111100110;
   2162: result <= 12'b010111100110;
   2163: result <= 12'b010111100111;
   2164: result <= 12'b010111100111;
   2165: result <= 12'b010111101000;
   2166: result <= 12'b010111101000;
   2167: result <= 12'b010111101001;
   2168: result <= 12'b010111101001;
   2169: result <= 12'b010111101010;
   2170: result <= 12'b010111101010;
   2171: result <= 12'b010111101011;
   2172: result <= 12'b010111101011;
   2173: result <= 12'b010111101100;
   2174: result <= 12'b010111101100;
   2175: result <= 12'b010111101101;
   2176: result <= 12'b010111101101;
   2177: result <= 12'b010111101110;
   2178: result <= 12'b010111101111;
   2179: result <= 12'b010111101111;
   2180: result <= 12'b010111110000;
   2181: result <= 12'b010111110000;
   2182: result <= 12'b010111110001;
   2183: result <= 12'b010111110001;
   2184: result <= 12'b010111110010;
   2185: result <= 12'b010111110010;
   2186: result <= 12'b010111110011;
   2187: result <= 12'b010111110011;
   2188: result <= 12'b010111110100;
   2189: result <= 12'b010111110100;
   2190: result <= 12'b010111110101;
   2191: result <= 12'b010111110101;
   2192: result <= 12'b010111110110;
   2193: result <= 12'b010111110110;
   2194: result <= 12'b010111110111;
   2195: result <= 12'b010111110111;
   2196: result <= 12'b010111111000;
   2197: result <= 12'b010111111000;
   2198: result <= 12'b010111111001;
   2199: result <= 12'b010111111010;
   2200: result <= 12'b010111111010;
   2201: result <= 12'b010111111011;
   2202: result <= 12'b010111111011;
   2203: result <= 12'b010111111100;
   2204: result <= 12'b010111111100;
   2205: result <= 12'b010111111101;
   2206: result <= 12'b010111111101;
   2207: result <= 12'b010111111110;
   2208: result <= 12'b010111111110;
   2209: result <= 12'b010111111111;
   2210: result <= 12'b010111111111;
   2211: result <= 12'b011000000000;
   2212: result <= 12'b011000000000;
   2213: result <= 12'b011000000001;
   2214: result <= 12'b011000000001;
   2215: result <= 12'b011000000010;
   2216: result <= 12'b011000000010;
   2217: result <= 12'b011000000011;
   2218: result <= 12'b011000000011;
   2219: result <= 12'b011000000100;
   2220: result <= 12'b011000000100;
   2221: result <= 12'b011000000101;
   2222: result <= 12'b011000000101;
   2223: result <= 12'b011000000110;
   2224: result <= 12'b011000000111;
   2225: result <= 12'b011000000111;
   2226: result <= 12'b011000001000;
   2227: result <= 12'b011000001000;
   2228: result <= 12'b011000001001;
   2229: result <= 12'b011000001001;
   2230: result <= 12'b011000001010;
   2231: result <= 12'b011000001010;
   2232: result <= 12'b011000001011;
   2233: result <= 12'b011000001011;
   2234: result <= 12'b011000001100;
   2235: result <= 12'b011000001100;
   2236: result <= 12'b011000001101;
   2237: result <= 12'b011000001101;
   2238: result <= 12'b011000001110;
   2239: result <= 12'b011000001110;
   2240: result <= 12'b011000001111;
   2241: result <= 12'b011000001111;
   2242: result <= 12'b011000010000;
   2243: result <= 12'b011000010000;
   2244: result <= 12'b011000010001;
   2245: result <= 12'b011000010001;
   2246: result <= 12'b011000010010;
   2247: result <= 12'b011000010010;
   2248: result <= 12'b011000010011;
   2249: result <= 12'b011000010011;
   2250: result <= 12'b011000010100;
   2251: result <= 12'b011000010100;
   2252: result <= 12'b011000010101;
   2253: result <= 12'b011000010101;
   2254: result <= 12'b011000010110;
   2255: result <= 12'b011000010110;
   2256: result <= 12'b011000010111;
   2257: result <= 12'b011000010111;
   2258: result <= 12'b011000011000;
   2259: result <= 12'b011000011000;
   2260: result <= 12'b011000011001;
   2261: result <= 12'b011000011001;
   2262: result <= 12'b011000011010;
   2263: result <= 12'b011000011011;
   2264: result <= 12'b011000011011;
   2265: result <= 12'b011000011100;
   2266: result <= 12'b011000011100;
   2267: result <= 12'b011000011101;
   2268: result <= 12'b011000011101;
   2269: result <= 12'b011000011110;
   2270: result <= 12'b011000011110;
   2271: result <= 12'b011000011111;
   2272: result <= 12'b011000011111;
   2273: result <= 12'b011000100000;
   2274: result <= 12'b011000100000;
   2275: result <= 12'b011000100001;
   2276: result <= 12'b011000100001;
   2277: result <= 12'b011000100010;
   2278: result <= 12'b011000100010;
   2279: result <= 12'b011000100011;
   2280: result <= 12'b011000100011;
   2281: result <= 12'b011000100100;
   2282: result <= 12'b011000100100;
   2283: result <= 12'b011000100101;
   2284: result <= 12'b011000100101;
   2285: result <= 12'b011000100110;
   2286: result <= 12'b011000100110;
   2287: result <= 12'b011000100111;
   2288: result <= 12'b011000100111;
   2289: result <= 12'b011000101000;
   2290: result <= 12'b011000101000;
   2291: result <= 12'b011000101001;
   2292: result <= 12'b011000101001;
   2293: result <= 12'b011000101010;
   2294: result <= 12'b011000101010;
   2295: result <= 12'b011000101011;
   2296: result <= 12'b011000101011;
   2297: result <= 12'b011000101100;
   2298: result <= 12'b011000101100;
   2299: result <= 12'b011000101101;
   2300: result <= 12'b011000101101;
   2301: result <= 12'b011000101110;
   2302: result <= 12'b011000101110;
   2303: result <= 12'b011000101111;
   2304: result <= 12'b011000101111;
   2305: result <= 12'b011000110000;
   2306: result <= 12'b011000110000;
   2307: result <= 12'b011000110001;
   2308: result <= 12'b011000110001;
   2309: result <= 12'b011000110010;
   2310: result <= 12'b011000110010;
   2311: result <= 12'b011000110011;
   2312: result <= 12'b011000110011;
   2313: result <= 12'b011000110100;
   2314: result <= 12'b011000110100;
   2315: result <= 12'b011000110101;
   2316: result <= 12'b011000110101;
   2317: result <= 12'b011000110110;
   2318: result <= 12'b011000110110;
   2319: result <= 12'b011000110111;
   2320: result <= 12'b011000110111;
   2321: result <= 12'b011000111000;
   2322: result <= 12'b011000111000;
   2323: result <= 12'b011000111001;
   2324: result <= 12'b011000111001;
   2325: result <= 12'b011000111010;
   2326: result <= 12'b011000111010;
   2327: result <= 12'b011000111011;
   2328: result <= 12'b011000111011;
   2329: result <= 12'b011000111100;
   2330: result <= 12'b011000111100;
   2331: result <= 12'b011000111100;
   2332: result <= 12'b011000111101;
   2333: result <= 12'b011000111101;
   2334: result <= 12'b011000111110;
   2335: result <= 12'b011000111110;
   2336: result <= 12'b011000111111;
   2337: result <= 12'b011000111111;
   2338: result <= 12'b011001000000;
   2339: result <= 12'b011001000000;
   2340: result <= 12'b011001000001;
   2341: result <= 12'b011001000001;
   2342: result <= 12'b011001000010;
   2343: result <= 12'b011001000010;
   2344: result <= 12'b011001000011;
   2345: result <= 12'b011001000011;
   2346: result <= 12'b011001000100;
   2347: result <= 12'b011001000100;
   2348: result <= 12'b011001000101;
   2349: result <= 12'b011001000101;
   2350: result <= 12'b011001000110;
   2351: result <= 12'b011001000110;
   2352: result <= 12'b011001000111;
   2353: result <= 12'b011001000111;
   2354: result <= 12'b011001001000;
   2355: result <= 12'b011001001000;
   2356: result <= 12'b011001001001;
   2357: result <= 12'b011001001001;
   2358: result <= 12'b011001001010;
   2359: result <= 12'b011001001010;
   2360: result <= 12'b011001001011;
   2361: result <= 12'b011001001011;
   2362: result <= 12'b011001001100;
   2363: result <= 12'b011001001100;
   2364: result <= 12'b011001001101;
   2365: result <= 12'b011001001101;
   2366: result <= 12'b011001001110;
   2367: result <= 12'b011001001110;
   2368: result <= 12'b011001001111;
   2369: result <= 12'b011001001111;
   2370: result <= 12'b011001001111;
   2371: result <= 12'b011001010000;
   2372: result <= 12'b011001010000;
   2373: result <= 12'b011001010001;
   2374: result <= 12'b011001010001;
   2375: result <= 12'b011001010010;
   2376: result <= 12'b011001010010;
   2377: result <= 12'b011001010011;
   2378: result <= 12'b011001010011;
   2379: result <= 12'b011001010100;
   2380: result <= 12'b011001010100;
   2381: result <= 12'b011001010101;
   2382: result <= 12'b011001010101;
   2383: result <= 12'b011001010110;
   2384: result <= 12'b011001010110;
   2385: result <= 12'b011001010111;
   2386: result <= 12'b011001010111;
   2387: result <= 12'b011001011000;
   2388: result <= 12'b011001011000;
   2389: result <= 12'b011001011001;
   2390: result <= 12'b011001011001;
   2391: result <= 12'b011001011010;
   2392: result <= 12'b011001011010;
   2393: result <= 12'b011001011011;
   2394: result <= 12'b011001011011;
   2395: result <= 12'b011001011011;
   2396: result <= 12'b011001011100;
   2397: result <= 12'b011001011100;
   2398: result <= 12'b011001011101;
   2399: result <= 12'b011001011101;
   2400: result <= 12'b011001011110;
   2401: result <= 12'b011001011110;
   2402: result <= 12'b011001011111;
   2403: result <= 12'b011001011111;
   2404: result <= 12'b011001100000;
   2405: result <= 12'b011001100000;
   2406: result <= 12'b011001100001;
   2407: result <= 12'b011001100001;
   2408: result <= 12'b011001100010;
   2409: result <= 12'b011001100010;
   2410: result <= 12'b011001100011;
   2411: result <= 12'b011001100011;
   2412: result <= 12'b011001100100;
   2413: result <= 12'b011001100100;
   2414: result <= 12'b011001100101;
   2415: result <= 12'b011001100101;
   2416: result <= 12'b011001100101;
   2417: result <= 12'b011001100110;
   2418: result <= 12'b011001100110;
   2419: result <= 12'b011001100111;
   2420: result <= 12'b011001100111;
   2421: result <= 12'b011001101000;
   2422: result <= 12'b011001101000;
   2423: result <= 12'b011001101001;
   2424: result <= 12'b011001101001;
   2425: result <= 12'b011001101010;
   2426: result <= 12'b011001101010;
   2427: result <= 12'b011001101011;
   2428: result <= 12'b011001101011;
   2429: result <= 12'b011001101100;
   2430: result <= 12'b011001101100;
   2431: result <= 12'b011001101101;
   2432: result <= 12'b011001101101;
   2433: result <= 12'b011001101101;
   2434: result <= 12'b011001101110;
   2435: result <= 12'b011001101110;
   2436: result <= 12'b011001101111;
   2437: result <= 12'b011001101111;
   2438: result <= 12'b011001110000;
   2439: result <= 12'b011001110000;
   2440: result <= 12'b011001110001;
   2441: result <= 12'b011001110001;
   2442: result <= 12'b011001110010;
   2443: result <= 12'b011001110010;
   2444: result <= 12'b011001110011;
   2445: result <= 12'b011001110011;
   2446: result <= 12'b011001110011;
   2447: result <= 12'b011001110100;
   2448: result <= 12'b011001110100;
   2449: result <= 12'b011001110101;
   2450: result <= 12'b011001110101;
   2451: result <= 12'b011001110110;
   2452: result <= 12'b011001110110;
   2453: result <= 12'b011001110111;
   2454: result <= 12'b011001110111;
   2455: result <= 12'b011001111000;
   2456: result <= 12'b011001111000;
   2457: result <= 12'b011001111001;
   2458: result <= 12'b011001111001;
   2459: result <= 12'b011001111010;
   2460: result <= 12'b011001111010;
   2461: result <= 12'b011001111010;
   2462: result <= 12'b011001111011;
   2463: result <= 12'b011001111011;
   2464: result <= 12'b011001111100;
   2465: result <= 12'b011001111100;
   2466: result <= 12'b011001111101;
   2467: result <= 12'b011001111101;
   2468: result <= 12'b011001111110;
   2469: result <= 12'b011001111110;
   2470: result <= 12'b011001111111;
   2471: result <= 12'b011001111111;
   2472: result <= 12'b011001111111;
   2473: result <= 12'b011010000000;
   2474: result <= 12'b011010000000;
   2475: result <= 12'b011010000001;
   2476: result <= 12'b011010000001;
   2477: result <= 12'b011010000010;
   2478: result <= 12'b011010000010;
   2479: result <= 12'b011010000011;
   2480: result <= 12'b011010000011;
   2481: result <= 12'b011010000100;
   2482: result <= 12'b011010000100;
   2483: result <= 12'b011010000101;
   2484: result <= 12'b011010000101;
   2485: result <= 12'b011010000101;
   2486: result <= 12'b011010000110;
   2487: result <= 12'b011010000110;
   2488: result <= 12'b011010000111;
   2489: result <= 12'b011010000111;
   2490: result <= 12'b011010001000;
   2491: result <= 12'b011010001000;
   2492: result <= 12'b011010001001;
   2493: result <= 12'b011010001001;
   2494: result <= 12'b011010001010;
   2495: result <= 12'b011010001010;
   2496: result <= 12'b011010001010;
   2497: result <= 12'b011010001011;
   2498: result <= 12'b011010001011;
   2499: result <= 12'b011010001100;
   2500: result <= 12'b011010001100;
   2501: result <= 12'b011010001101;
   2502: result <= 12'b011010001101;
   2503: result <= 12'b011010001110;
   2504: result <= 12'b011010001110;
   2505: result <= 12'b011010001110;
   2506: result <= 12'b011010001111;
   2507: result <= 12'b011010001111;
   2508: result <= 12'b011010010000;
   2509: result <= 12'b011010010000;
   2510: result <= 12'b011010010001;
   2511: result <= 12'b011010010001;
   2512: result <= 12'b011010010010;
   2513: result <= 12'b011010010010;
   2514: result <= 12'b011010010011;
   2515: result <= 12'b011010010011;
   2516: result <= 12'b011010010011;
   2517: result <= 12'b011010010100;
   2518: result <= 12'b011010010100;
   2519: result <= 12'b011010010101;
   2520: result <= 12'b011010010101;
   2521: result <= 12'b011010010110;
   2522: result <= 12'b011010010110;
   2523: result <= 12'b011010010111;
   2524: result <= 12'b011010010111;
   2525: result <= 12'b011010010111;
   2526: result <= 12'b011010011000;
   2527: result <= 12'b011010011000;
   2528: result <= 12'b011010011001;
   2529: result <= 12'b011010011001;
   2530: result <= 12'b011010011010;
   2531: result <= 12'b011010011010;
   2532: result <= 12'b011010011011;
   2533: result <= 12'b011010011011;
   2534: result <= 12'b011010011011;
   2535: result <= 12'b011010011100;
   2536: result <= 12'b011010011100;
   2537: result <= 12'b011010011101;
   2538: result <= 12'b011010011101;
   2539: result <= 12'b011010011110;
   2540: result <= 12'b011010011110;
   2541: result <= 12'b011010011111;
   2542: result <= 12'b011010011111;
   2543: result <= 12'b011010011111;
   2544: result <= 12'b011010100000;
   2545: result <= 12'b011010100000;
   2546: result <= 12'b011010100001;
   2547: result <= 12'b011010100001;
   2548: result <= 12'b011010100010;
   2549: result <= 12'b011010100010;
   2550: result <= 12'b011010100010;
   2551: result <= 12'b011010100011;
   2552: result <= 12'b011010100011;
   2553: result <= 12'b011010100100;
   2554: result <= 12'b011010100100;
   2555: result <= 12'b011010100101;
   2556: result <= 12'b011010100101;
   2557: result <= 12'b011010100110;
   2558: result <= 12'b011010100110;
   2559: result <= 12'b011010100110;
   2560: result <= 12'b011010100111;
   2561: result <= 12'b011010100111;
   2562: result <= 12'b011010101000;
   2563: result <= 12'b011010101000;
   2564: result <= 12'b011010101001;
   2565: result <= 12'b011010101001;
   2566: result <= 12'b011010101001;
   2567: result <= 12'b011010101010;
   2568: result <= 12'b011010101010;
   2569: result <= 12'b011010101011;
   2570: result <= 12'b011010101011;
   2571: result <= 12'b011010101100;
   2572: result <= 12'b011010101100;
   2573: result <= 12'b011010101101;
   2574: result <= 12'b011010101101;
   2575: result <= 12'b011010101101;
   2576: result <= 12'b011010101110;
   2577: result <= 12'b011010101110;
   2578: result <= 12'b011010101111;
   2579: result <= 12'b011010101111;
   2580: result <= 12'b011010110000;
   2581: result <= 12'b011010110000;
   2582: result <= 12'b011010110000;
   2583: result <= 12'b011010110001;
   2584: result <= 12'b011010110001;
   2585: result <= 12'b011010110010;
   2586: result <= 12'b011010110010;
   2587: result <= 12'b011010110011;
   2588: result <= 12'b011010110011;
   2589: result <= 12'b011010110011;
   2590: result <= 12'b011010110100;
   2591: result <= 12'b011010110100;
   2592: result <= 12'b011010110101;
   2593: result <= 12'b011010110101;
   2594: result <= 12'b011010110110;
   2595: result <= 12'b011010110110;
   2596: result <= 12'b011010110110;
   2597: result <= 12'b011010110111;
   2598: result <= 12'b011010110111;
   2599: result <= 12'b011010111000;
   2600: result <= 12'b011010111000;
   2601: result <= 12'b011010111001;
   2602: result <= 12'b011010111001;
   2603: result <= 12'b011010111001;
   2604: result <= 12'b011010111010;
   2605: result <= 12'b011010111010;
   2606: result <= 12'b011010111011;
   2607: result <= 12'b011010111011;
   2608: result <= 12'b011010111100;
   2609: result <= 12'b011010111100;
   2610: result <= 12'b011010111100;
   2611: result <= 12'b011010111101;
   2612: result <= 12'b011010111101;
   2613: result <= 12'b011010111110;
   2614: result <= 12'b011010111110;
   2615: result <= 12'b011010111110;
   2616: result <= 12'b011010111111;
   2617: result <= 12'b011010111111;
   2618: result <= 12'b011011000000;
   2619: result <= 12'b011011000000;
   2620: result <= 12'b011011000001;
   2621: result <= 12'b011011000001;
   2622: result <= 12'b011011000001;
   2623: result <= 12'b011011000010;
   2624: result <= 12'b011011000010;
   2625: result <= 12'b011011000011;
   2626: result <= 12'b011011000011;
   2627: result <= 12'b011011000100;
   2628: result <= 12'b011011000100;
   2629: result <= 12'b011011000100;
   2630: result <= 12'b011011000101;
   2631: result <= 12'b011011000101;
   2632: result <= 12'b011011000110;
   2633: result <= 12'b011011000110;
   2634: result <= 12'b011011000110;
   2635: result <= 12'b011011000111;
   2636: result <= 12'b011011000111;
   2637: result <= 12'b011011001000;
   2638: result <= 12'b011011001000;
   2639: result <= 12'b011011001001;
   2640: result <= 12'b011011001001;
   2641: result <= 12'b011011001001;
   2642: result <= 12'b011011001010;
   2643: result <= 12'b011011001010;
   2644: result <= 12'b011011001011;
   2645: result <= 12'b011011001011;
   2646: result <= 12'b011011001011;
   2647: result <= 12'b011011001100;
   2648: result <= 12'b011011001100;
   2649: result <= 12'b011011001101;
   2650: result <= 12'b011011001101;
   2651: result <= 12'b011011001110;
   2652: result <= 12'b011011001110;
   2653: result <= 12'b011011001110;
   2654: result <= 12'b011011001111;
   2655: result <= 12'b011011001111;
   2656: result <= 12'b011011010000;
   2657: result <= 12'b011011010000;
   2658: result <= 12'b011011010000;
   2659: result <= 12'b011011010001;
   2660: result <= 12'b011011010001;
   2661: result <= 12'b011011010010;
   2662: result <= 12'b011011010010;
   2663: result <= 12'b011011010010;
   2664: result <= 12'b011011010011;
   2665: result <= 12'b011011010011;
   2666: result <= 12'b011011010100;
   2667: result <= 12'b011011010100;
   2668: result <= 12'b011011010101;
   2669: result <= 12'b011011010101;
   2670: result <= 12'b011011010101;
   2671: result <= 12'b011011010110;
   2672: result <= 12'b011011010110;
   2673: result <= 12'b011011010111;
   2674: result <= 12'b011011010111;
   2675: result <= 12'b011011010111;
   2676: result <= 12'b011011011000;
   2677: result <= 12'b011011011000;
   2678: result <= 12'b011011011001;
   2679: result <= 12'b011011011001;
   2680: result <= 12'b011011011001;
   2681: result <= 12'b011011011010;
   2682: result <= 12'b011011011010;
   2683: result <= 12'b011011011011;
   2684: result <= 12'b011011011011;
   2685: result <= 12'b011011011011;
   2686: result <= 12'b011011011100;
   2687: result <= 12'b011011011100;
   2688: result <= 12'b011011011101;
   2689: result <= 12'b011011011101;
   2690: result <= 12'b011011011101;
   2691: result <= 12'b011011011110;
   2692: result <= 12'b011011011110;
   2693: result <= 12'b011011011111;
   2694: result <= 12'b011011011111;
   2695: result <= 12'b011011011111;
   2696: result <= 12'b011011100000;
   2697: result <= 12'b011011100000;
   2698: result <= 12'b011011100001;
   2699: result <= 12'b011011100001;
   2700: result <= 12'b011011100001;
   2701: result <= 12'b011011100010;
   2702: result <= 12'b011011100010;
   2703: result <= 12'b011011100011;
   2704: result <= 12'b011011100011;
   2705: result <= 12'b011011100011;
   2706: result <= 12'b011011100100;
   2707: result <= 12'b011011100100;
   2708: result <= 12'b011011100101;
   2709: result <= 12'b011011100101;
   2710: result <= 12'b011011100101;
   2711: result <= 12'b011011100110;
   2712: result <= 12'b011011100110;
   2713: result <= 12'b011011100111;
   2714: result <= 12'b011011100111;
   2715: result <= 12'b011011100111;
   2716: result <= 12'b011011101000;
   2717: result <= 12'b011011101000;
   2718: result <= 12'b011011101001;
   2719: result <= 12'b011011101001;
   2720: result <= 12'b011011101001;
   2721: result <= 12'b011011101010;
   2722: result <= 12'b011011101010;
   2723: result <= 12'b011011101011;
   2724: result <= 12'b011011101011;
   2725: result <= 12'b011011101011;
   2726: result <= 12'b011011101100;
   2727: result <= 12'b011011101100;
   2728: result <= 12'b011011101101;
   2729: result <= 12'b011011101101;
   2730: result <= 12'b011011101101;
   2731: result <= 12'b011011101110;
   2732: result <= 12'b011011101110;
   2733: result <= 12'b011011101111;
   2734: result <= 12'b011011101111;
   2735: result <= 12'b011011101111;
   2736: result <= 12'b011011110000;
   2737: result <= 12'b011011110000;
   2738: result <= 12'b011011110000;
   2739: result <= 12'b011011110001;
   2740: result <= 12'b011011110001;
   2741: result <= 12'b011011110010;
   2742: result <= 12'b011011110010;
   2743: result <= 12'b011011110010;
   2744: result <= 12'b011011110011;
   2745: result <= 12'b011011110011;
   2746: result <= 12'b011011110100;
   2747: result <= 12'b011011110100;
   2748: result <= 12'b011011110100;
   2749: result <= 12'b011011110101;
   2750: result <= 12'b011011110101;
   2751: result <= 12'b011011110110;
   2752: result <= 12'b011011110110;
   2753: result <= 12'b011011110110;
   2754: result <= 12'b011011110111;
   2755: result <= 12'b011011110111;
   2756: result <= 12'b011011110111;
   2757: result <= 12'b011011111000;
   2758: result <= 12'b011011111000;
   2759: result <= 12'b011011111001;
   2760: result <= 12'b011011111001;
   2761: result <= 12'b011011111001;
   2762: result <= 12'b011011111010;
   2763: result <= 12'b011011111010;
   2764: result <= 12'b011011111011;
   2765: result <= 12'b011011111011;
   2766: result <= 12'b011011111011;
   2767: result <= 12'b011011111100;
   2768: result <= 12'b011011111100;
   2769: result <= 12'b011011111100;
   2770: result <= 12'b011011111101;
   2771: result <= 12'b011011111101;
   2772: result <= 12'b011011111110;
   2773: result <= 12'b011011111110;
   2774: result <= 12'b011011111110;
   2775: result <= 12'b011011111111;
   2776: result <= 12'b011011111111;
   2777: result <= 12'b011100000000;
   2778: result <= 12'b011100000000;
   2779: result <= 12'b011100000000;
   2780: result <= 12'b011100000001;
   2781: result <= 12'b011100000001;
   2782: result <= 12'b011100000001;
   2783: result <= 12'b011100000010;
   2784: result <= 12'b011100000010;
   2785: result <= 12'b011100000011;
   2786: result <= 12'b011100000011;
   2787: result <= 12'b011100000011;
   2788: result <= 12'b011100000100;
   2789: result <= 12'b011100000100;
   2790: result <= 12'b011100000100;
   2791: result <= 12'b011100000101;
   2792: result <= 12'b011100000101;
   2793: result <= 12'b011100000110;
   2794: result <= 12'b011100000110;
   2795: result <= 12'b011100000110;
   2796: result <= 12'b011100000111;
   2797: result <= 12'b011100000111;
   2798: result <= 12'b011100000111;
   2799: result <= 12'b011100001000;
   2800: result <= 12'b011100001000;
   2801: result <= 12'b011100001001;
   2802: result <= 12'b011100001001;
   2803: result <= 12'b011100001001;
   2804: result <= 12'b011100001010;
   2805: result <= 12'b011100001010;
   2806: result <= 12'b011100001010;
   2807: result <= 12'b011100001011;
   2808: result <= 12'b011100001011;
   2809: result <= 12'b011100001100;
   2810: result <= 12'b011100001100;
   2811: result <= 12'b011100001100;
   2812: result <= 12'b011100001101;
   2813: result <= 12'b011100001101;
   2814: result <= 12'b011100001101;
   2815: result <= 12'b011100001110;
   2816: result <= 12'b011100001110;
   2817: result <= 12'b011100001111;
   2818: result <= 12'b011100001111;
   2819: result <= 12'b011100001111;
   2820: result <= 12'b011100010000;
   2821: result <= 12'b011100010000;
   2822: result <= 12'b011100010000;
   2823: result <= 12'b011100010001;
   2824: result <= 12'b011100010001;
   2825: result <= 12'b011100010001;
   2826: result <= 12'b011100010010;
   2827: result <= 12'b011100010010;
   2828: result <= 12'b011100010011;
   2829: result <= 12'b011100010011;
   2830: result <= 12'b011100010011;
   2831: result <= 12'b011100010100;
   2832: result <= 12'b011100010100;
   2833: result <= 12'b011100010100;
   2834: result <= 12'b011100010101;
   2835: result <= 12'b011100010101;
   2836: result <= 12'b011100010110;
   2837: result <= 12'b011100010110;
   2838: result <= 12'b011100010110;
   2839: result <= 12'b011100010111;
   2840: result <= 12'b011100010111;
   2841: result <= 12'b011100010111;
   2842: result <= 12'b011100011000;
   2843: result <= 12'b011100011000;
   2844: result <= 12'b011100011000;
   2845: result <= 12'b011100011001;
   2846: result <= 12'b011100011001;
   2847: result <= 12'b011100011010;
   2848: result <= 12'b011100011010;
   2849: result <= 12'b011100011010;
   2850: result <= 12'b011100011011;
   2851: result <= 12'b011100011011;
   2852: result <= 12'b011100011011;
   2853: result <= 12'b011100011100;
   2854: result <= 12'b011100011100;
   2855: result <= 12'b011100011100;
   2856: result <= 12'b011100011101;
   2857: result <= 12'b011100011101;
   2858: result <= 12'b011100011101;
   2859: result <= 12'b011100011110;
   2860: result <= 12'b011100011110;
   2861: result <= 12'b011100011111;
   2862: result <= 12'b011100011111;
   2863: result <= 12'b011100011111;
   2864: result <= 12'b011100100000;
   2865: result <= 12'b011100100000;
   2866: result <= 12'b011100100000;
   2867: result <= 12'b011100100001;
   2868: result <= 12'b011100100001;
   2869: result <= 12'b011100100001;
   2870: result <= 12'b011100100010;
   2871: result <= 12'b011100100010;
   2872: result <= 12'b011100100010;
   2873: result <= 12'b011100100011;
   2874: result <= 12'b011100100011;
   2875: result <= 12'b011100100100;
   2876: result <= 12'b011100100100;
   2877: result <= 12'b011100100100;
   2878: result <= 12'b011100100101;
   2879: result <= 12'b011100100101;
   2880: result <= 12'b011100100101;
   2881: result <= 12'b011100100110;
   2882: result <= 12'b011100100110;
   2883: result <= 12'b011100100110;
   2884: result <= 12'b011100100111;
   2885: result <= 12'b011100100111;
   2886: result <= 12'b011100100111;
   2887: result <= 12'b011100101000;
   2888: result <= 12'b011100101000;
   2889: result <= 12'b011100101000;
   2890: result <= 12'b011100101001;
   2891: result <= 12'b011100101001;
   2892: result <= 12'b011100101010;
   2893: result <= 12'b011100101010;
   2894: result <= 12'b011100101010;
   2895: result <= 12'b011100101011;
   2896: result <= 12'b011100101011;
   2897: result <= 12'b011100101011;
   2898: result <= 12'b011100101100;
   2899: result <= 12'b011100101100;
   2900: result <= 12'b011100101100;
   2901: result <= 12'b011100101101;
   2902: result <= 12'b011100101101;
   2903: result <= 12'b011100101101;
   2904: result <= 12'b011100101110;
   2905: result <= 12'b011100101110;
   2906: result <= 12'b011100101110;
   2907: result <= 12'b011100101111;
   2908: result <= 12'b011100101111;
   2909: result <= 12'b011100101111;
   2910: result <= 12'b011100110000;
   2911: result <= 12'b011100110000;
   2912: result <= 12'b011100110000;
   2913: result <= 12'b011100110001;
   2914: result <= 12'b011100110001;
   2915: result <= 12'b011100110010;
   2916: result <= 12'b011100110010;
   2917: result <= 12'b011100110010;
   2918: result <= 12'b011100110011;
   2919: result <= 12'b011100110011;
   2920: result <= 12'b011100110011;
   2921: result <= 12'b011100110100;
   2922: result <= 12'b011100110100;
   2923: result <= 12'b011100110100;
   2924: result <= 12'b011100110101;
   2925: result <= 12'b011100110101;
   2926: result <= 12'b011100110101;
   2927: result <= 12'b011100110110;
   2928: result <= 12'b011100110110;
   2929: result <= 12'b011100110110;
   2930: result <= 12'b011100110111;
   2931: result <= 12'b011100110111;
   2932: result <= 12'b011100110111;
   2933: result <= 12'b011100111000;
   2934: result <= 12'b011100111000;
   2935: result <= 12'b011100111000;
   2936: result <= 12'b011100111001;
   2937: result <= 12'b011100111001;
   2938: result <= 12'b011100111001;
   2939: result <= 12'b011100111010;
   2940: result <= 12'b011100111010;
   2941: result <= 12'b011100111010;
   2942: result <= 12'b011100111011;
   2943: result <= 12'b011100111011;
   2944: result <= 12'b011100111011;
   2945: result <= 12'b011100111100;
   2946: result <= 12'b011100111100;
   2947: result <= 12'b011100111100;
   2948: result <= 12'b011100111101;
   2949: result <= 12'b011100111101;
   2950: result <= 12'b011100111101;
   2951: result <= 12'b011100111110;
   2952: result <= 12'b011100111110;
   2953: result <= 12'b011100111110;
   2954: result <= 12'b011100111111;
   2955: result <= 12'b011100111111;
   2956: result <= 12'b011100111111;
   2957: result <= 12'b011101000000;
   2958: result <= 12'b011101000000;
   2959: result <= 12'b011101000000;
   2960: result <= 12'b011101000001;
   2961: result <= 12'b011101000001;
   2962: result <= 12'b011101000001;
   2963: result <= 12'b011101000010;
   2964: result <= 12'b011101000010;
   2965: result <= 12'b011101000010;
   2966: result <= 12'b011101000011;
   2967: result <= 12'b011101000011;
   2968: result <= 12'b011101000011;
   2969: result <= 12'b011101000100;
   2970: result <= 12'b011101000100;
   2971: result <= 12'b011101000100;
   2972: result <= 12'b011101000101;
   2973: result <= 12'b011101000101;
   2974: result <= 12'b011101000101;
   2975: result <= 12'b011101000110;
   2976: result <= 12'b011101000110;
   2977: result <= 12'b011101000110;
   2978: result <= 12'b011101000111;
   2979: result <= 12'b011101000111;
   2980: result <= 12'b011101000111;
   2981: result <= 12'b011101001000;
   2982: result <= 12'b011101001000;
   2983: result <= 12'b011101001000;
   2984: result <= 12'b011101001001;
   2985: result <= 12'b011101001001;
   2986: result <= 12'b011101001001;
   2987: result <= 12'b011101001010;
   2988: result <= 12'b011101001010;
   2989: result <= 12'b011101001010;
   2990: result <= 12'b011101001011;
   2991: result <= 12'b011101001011;
   2992: result <= 12'b011101001011;
   2993: result <= 12'b011101001011;
   2994: result <= 12'b011101001100;
   2995: result <= 12'b011101001100;
   2996: result <= 12'b011101001100;
   2997: result <= 12'b011101001101;
   2998: result <= 12'b011101001101;
   2999: result <= 12'b011101001101;
   3000: result <= 12'b011101001110;
   3001: result <= 12'b011101001110;
   3002: result <= 12'b011101001110;
   3003: result <= 12'b011101001111;
   3004: result <= 12'b011101001111;
   3005: result <= 12'b011101001111;
   3006: result <= 12'b011101010000;
   3007: result <= 12'b011101010000;
   3008: result <= 12'b011101010000;
   3009: result <= 12'b011101010001;
   3010: result <= 12'b011101010001;
   3011: result <= 12'b011101010001;
   3012: result <= 12'b011101010010;
   3013: result <= 12'b011101010010;
   3014: result <= 12'b011101010010;
   3015: result <= 12'b011101010011;
   3016: result <= 12'b011101010011;
   3017: result <= 12'b011101010011;
   3018: result <= 12'b011101010011;
   3019: result <= 12'b011101010100;
   3020: result <= 12'b011101010100;
   3021: result <= 12'b011101010100;
   3022: result <= 12'b011101010101;
   3023: result <= 12'b011101010101;
   3024: result <= 12'b011101010101;
   3025: result <= 12'b011101010110;
   3026: result <= 12'b011101010110;
   3027: result <= 12'b011101010110;
   3028: result <= 12'b011101010111;
   3029: result <= 12'b011101010111;
   3030: result <= 12'b011101010111;
   3031: result <= 12'b011101011000;
   3032: result <= 12'b011101011000;
   3033: result <= 12'b011101011000;
   3034: result <= 12'b011101011000;
   3035: result <= 12'b011101011001;
   3036: result <= 12'b011101011001;
   3037: result <= 12'b011101011001;
   3038: result <= 12'b011101011010;
   3039: result <= 12'b011101011010;
   3040: result <= 12'b011101011010;
   3041: result <= 12'b011101011011;
   3042: result <= 12'b011101011011;
   3043: result <= 12'b011101011011;
   3044: result <= 12'b011101011100;
   3045: result <= 12'b011101011100;
   3046: result <= 12'b011101011100;
   3047: result <= 12'b011101011101;
   3048: result <= 12'b011101011101;
   3049: result <= 12'b011101011101;
   3050: result <= 12'b011101011101;
   3051: result <= 12'b011101011110;
   3052: result <= 12'b011101011110;
   3053: result <= 12'b011101011110;
   3054: result <= 12'b011101011111;
   3055: result <= 12'b011101011111;
   3056: result <= 12'b011101011111;
   3057: result <= 12'b011101100000;
   3058: result <= 12'b011101100000;
   3059: result <= 12'b011101100000;
   3060: result <= 12'b011101100000;
   3061: result <= 12'b011101100001;
   3062: result <= 12'b011101100001;
   3063: result <= 12'b011101100001;
   3064: result <= 12'b011101100010;
   3065: result <= 12'b011101100010;
   3066: result <= 12'b011101100010;
   3067: result <= 12'b011101100011;
   3068: result <= 12'b011101100011;
   3069: result <= 12'b011101100011;
   3070: result <= 12'b011101100100;
   3071: result <= 12'b011101100100;
   3072: result <= 12'b011101100100;
   3073: result <= 12'b011101100100;
   3074: result <= 12'b011101100101;
   3075: result <= 12'b011101100101;
   3076: result <= 12'b011101100101;
   3077: result <= 12'b011101100110;
   3078: result <= 12'b011101100110;
   3079: result <= 12'b011101100110;
   3080: result <= 12'b011101100111;
   3081: result <= 12'b011101100111;
   3082: result <= 12'b011101100111;
   3083: result <= 12'b011101100111;
   3084: result <= 12'b011101101000;
   3085: result <= 12'b011101101000;
   3086: result <= 12'b011101101000;
   3087: result <= 12'b011101101001;
   3088: result <= 12'b011101101001;
   3089: result <= 12'b011101101001;
   3090: result <= 12'b011101101001;
   3091: result <= 12'b011101101010;
   3092: result <= 12'b011101101010;
   3093: result <= 12'b011101101010;
   3094: result <= 12'b011101101011;
   3095: result <= 12'b011101101011;
   3096: result <= 12'b011101101011;
   3097: result <= 12'b011101101100;
   3098: result <= 12'b011101101100;
   3099: result <= 12'b011101101100;
   3100: result <= 12'b011101101100;
   3101: result <= 12'b011101101101;
   3102: result <= 12'b011101101101;
   3103: result <= 12'b011101101101;
   3104: result <= 12'b011101101110;
   3105: result <= 12'b011101101110;
   3106: result <= 12'b011101101110;
   3107: result <= 12'b011101101110;
   3108: result <= 12'b011101101111;
   3109: result <= 12'b011101101111;
   3110: result <= 12'b011101101111;
   3111: result <= 12'b011101110000;
   3112: result <= 12'b011101110000;
   3113: result <= 12'b011101110000;
   3114: result <= 12'b011101110000;
   3115: result <= 12'b011101110001;
   3116: result <= 12'b011101110001;
   3117: result <= 12'b011101110001;
   3118: result <= 12'b011101110010;
   3119: result <= 12'b011101110010;
   3120: result <= 12'b011101110010;
   3121: result <= 12'b011101110010;
   3122: result <= 12'b011101110011;
   3123: result <= 12'b011101110011;
   3124: result <= 12'b011101110011;
   3125: result <= 12'b011101110100;
   3126: result <= 12'b011101110100;
   3127: result <= 12'b011101110100;
   3128: result <= 12'b011101110100;
   3129: result <= 12'b011101110101;
   3130: result <= 12'b011101110101;
   3131: result <= 12'b011101110101;
   3132: result <= 12'b011101110110;
   3133: result <= 12'b011101110110;
   3134: result <= 12'b011101110110;
   3135: result <= 12'b011101110110;
   3136: result <= 12'b011101110111;
   3137: result <= 12'b011101110111;
   3138: result <= 12'b011101110111;
   3139: result <= 12'b011101111000;
   3140: result <= 12'b011101111000;
   3141: result <= 12'b011101111000;
   3142: result <= 12'b011101111000;
   3143: result <= 12'b011101111001;
   3144: result <= 12'b011101111001;
   3145: result <= 12'b011101111001;
   3146: result <= 12'b011101111010;
   3147: result <= 12'b011101111010;
   3148: result <= 12'b011101111010;
   3149: result <= 12'b011101111010;
   3150: result <= 12'b011101111011;
   3151: result <= 12'b011101111011;
   3152: result <= 12'b011101111011;
   3153: result <= 12'b011101111100;
   3154: result <= 12'b011101111100;
   3155: result <= 12'b011101111100;
   3156: result <= 12'b011101111100;
   3157: result <= 12'b011101111101;
   3158: result <= 12'b011101111101;
   3159: result <= 12'b011101111101;
   3160: result <= 12'b011101111101;
   3161: result <= 12'b011101111110;
   3162: result <= 12'b011101111110;
   3163: result <= 12'b011101111110;
   3164: result <= 12'b011101111111;
   3165: result <= 12'b011101111111;
   3166: result <= 12'b011101111111;
   3167: result <= 12'b011101111111;
   3168: result <= 12'b011110000000;
   3169: result <= 12'b011110000000;
   3170: result <= 12'b011110000000;
   3171: result <= 12'b011110000000;
   3172: result <= 12'b011110000001;
   3173: result <= 12'b011110000001;
   3174: result <= 12'b011110000001;
   3175: result <= 12'b011110000010;
   3176: result <= 12'b011110000010;
   3177: result <= 12'b011110000010;
   3178: result <= 12'b011110000010;
   3179: result <= 12'b011110000011;
   3180: result <= 12'b011110000011;
   3181: result <= 12'b011110000011;
   3182: result <= 12'b011110000011;
   3183: result <= 12'b011110000100;
   3184: result <= 12'b011110000100;
   3185: result <= 12'b011110000100;
   3186: result <= 12'b011110000101;
   3187: result <= 12'b011110000101;
   3188: result <= 12'b011110000101;
   3189: result <= 12'b011110000101;
   3190: result <= 12'b011110000110;
   3191: result <= 12'b011110000110;
   3192: result <= 12'b011110000110;
   3193: result <= 12'b011110000110;
   3194: result <= 12'b011110000111;
   3195: result <= 12'b011110000111;
   3196: result <= 12'b011110000111;
   3197: result <= 12'b011110000111;
   3198: result <= 12'b011110001000;
   3199: result <= 12'b011110001000;
   3200: result <= 12'b011110001000;
   3201: result <= 12'b011110001001;
   3202: result <= 12'b011110001001;
   3203: result <= 12'b011110001001;
   3204: result <= 12'b011110001001;
   3205: result <= 12'b011110001010;
   3206: result <= 12'b011110001010;
   3207: result <= 12'b011110001010;
   3208: result <= 12'b011110001010;
   3209: result <= 12'b011110001011;
   3210: result <= 12'b011110001011;
   3211: result <= 12'b011110001011;
   3212: result <= 12'b011110001011;
   3213: result <= 12'b011110001100;
   3214: result <= 12'b011110001100;
   3215: result <= 12'b011110001100;
   3216: result <= 12'b011110001100;
   3217: result <= 12'b011110001101;
   3218: result <= 12'b011110001101;
   3219: result <= 12'b011110001101;
   3220: result <= 12'b011110001110;
   3221: result <= 12'b011110001110;
   3222: result <= 12'b011110001110;
   3223: result <= 12'b011110001110;
   3224: result <= 12'b011110001111;
   3225: result <= 12'b011110001111;
   3226: result <= 12'b011110001111;
   3227: result <= 12'b011110001111;
   3228: result <= 12'b011110010000;
   3229: result <= 12'b011110010000;
   3230: result <= 12'b011110010000;
   3231: result <= 12'b011110010000;
   3232: result <= 12'b011110010001;
   3233: result <= 12'b011110010001;
   3234: result <= 12'b011110010001;
   3235: result <= 12'b011110010001;
   3236: result <= 12'b011110010010;
   3237: result <= 12'b011110010010;
   3238: result <= 12'b011110010010;
   3239: result <= 12'b011110010010;
   3240: result <= 12'b011110010011;
   3241: result <= 12'b011110010011;
   3242: result <= 12'b011110010011;
   3243: result <= 12'b011110010011;
   3244: result <= 12'b011110010100;
   3245: result <= 12'b011110010100;
   3246: result <= 12'b011110010100;
   3247: result <= 12'b011110010100;
   3248: result <= 12'b011110010101;
   3249: result <= 12'b011110010101;
   3250: result <= 12'b011110010101;
   3251: result <= 12'b011110010101;
   3252: result <= 12'b011110010110;
   3253: result <= 12'b011110010110;
   3254: result <= 12'b011110010110;
   3255: result <= 12'b011110010110;
   3256: result <= 12'b011110010111;
   3257: result <= 12'b011110010111;
   3258: result <= 12'b011110010111;
   3259: result <= 12'b011110010111;
   3260: result <= 12'b011110011000;
   3261: result <= 12'b011110011000;
   3262: result <= 12'b011110011000;
   3263: result <= 12'b011110011000;
   3264: result <= 12'b011110011001;
   3265: result <= 12'b011110011001;
   3266: result <= 12'b011110011001;
   3267: result <= 12'b011110011001;
   3268: result <= 12'b011110011010;
   3269: result <= 12'b011110011010;
   3270: result <= 12'b011110011010;
   3271: result <= 12'b011110011010;
   3272: result <= 12'b011110011011;
   3273: result <= 12'b011110011011;
   3274: result <= 12'b011110011011;
   3275: result <= 12'b011110011011;
   3276: result <= 12'b011110011100;
   3277: result <= 12'b011110011100;
   3278: result <= 12'b011110011100;
   3279: result <= 12'b011110011100;
   3280: result <= 12'b011110011101;
   3281: result <= 12'b011110011101;
   3282: result <= 12'b011110011101;
   3283: result <= 12'b011110011101;
   3284: result <= 12'b011110011110;
   3285: result <= 12'b011110011110;
   3286: result <= 12'b011110011110;
   3287: result <= 12'b011110011110;
   3288: result <= 12'b011110011110;
   3289: result <= 12'b011110011111;
   3290: result <= 12'b011110011111;
   3291: result <= 12'b011110011111;
   3292: result <= 12'b011110011111;
   3293: result <= 12'b011110100000;
   3294: result <= 12'b011110100000;
   3295: result <= 12'b011110100000;
   3296: result <= 12'b011110100000;
   3297: result <= 12'b011110100001;
   3298: result <= 12'b011110100001;
   3299: result <= 12'b011110100001;
   3300: result <= 12'b011110100001;
   3301: result <= 12'b011110100010;
   3302: result <= 12'b011110100010;
   3303: result <= 12'b011110100010;
   3304: result <= 12'b011110100010;
   3305: result <= 12'b011110100010;
   3306: result <= 12'b011110100011;
   3307: result <= 12'b011110100011;
   3308: result <= 12'b011110100011;
   3309: result <= 12'b011110100011;
   3310: result <= 12'b011110100100;
   3311: result <= 12'b011110100100;
   3312: result <= 12'b011110100100;
   3313: result <= 12'b011110100100;
   3314: result <= 12'b011110100101;
   3315: result <= 12'b011110100101;
   3316: result <= 12'b011110100101;
   3317: result <= 12'b011110100101;
   3318: result <= 12'b011110100110;
   3319: result <= 12'b011110100110;
   3320: result <= 12'b011110100110;
   3321: result <= 12'b011110100110;
   3322: result <= 12'b011110100110;
   3323: result <= 12'b011110100111;
   3324: result <= 12'b011110100111;
   3325: result <= 12'b011110100111;
   3326: result <= 12'b011110100111;
   3327: result <= 12'b011110101000;
   3328: result <= 12'b011110101000;
   3329: result <= 12'b011110101000;
   3330: result <= 12'b011110101000;
   3331: result <= 12'b011110101000;
   3332: result <= 12'b011110101001;
   3333: result <= 12'b011110101001;
   3334: result <= 12'b011110101001;
   3335: result <= 12'b011110101001;
   3336: result <= 12'b011110101010;
   3337: result <= 12'b011110101010;
   3338: result <= 12'b011110101010;
   3339: result <= 12'b011110101010;
   3340: result <= 12'b011110101011;
   3341: result <= 12'b011110101011;
   3342: result <= 12'b011110101011;
   3343: result <= 12'b011110101011;
   3344: result <= 12'b011110101011;
   3345: result <= 12'b011110101100;
   3346: result <= 12'b011110101100;
   3347: result <= 12'b011110101100;
   3348: result <= 12'b011110101100;
   3349: result <= 12'b011110101101;
   3350: result <= 12'b011110101101;
   3351: result <= 12'b011110101101;
   3352: result <= 12'b011110101101;
   3353: result <= 12'b011110101101;
   3354: result <= 12'b011110101110;
   3355: result <= 12'b011110101110;
   3356: result <= 12'b011110101110;
   3357: result <= 12'b011110101110;
   3358: result <= 12'b011110101111;
   3359: result <= 12'b011110101111;
   3360: result <= 12'b011110101111;
   3361: result <= 12'b011110101111;
   3362: result <= 12'b011110101111;
   3363: result <= 12'b011110110000;
   3364: result <= 12'b011110110000;
   3365: result <= 12'b011110110000;
   3366: result <= 12'b011110110000;
   3367: result <= 12'b011110110000;
   3368: result <= 12'b011110110001;
   3369: result <= 12'b011110110001;
   3370: result <= 12'b011110110001;
   3371: result <= 12'b011110110001;
   3372: result <= 12'b011110110010;
   3373: result <= 12'b011110110010;
   3374: result <= 12'b011110110010;
   3375: result <= 12'b011110110010;
   3376: result <= 12'b011110110010;
   3377: result <= 12'b011110110011;
   3378: result <= 12'b011110110011;
   3379: result <= 12'b011110110011;
   3380: result <= 12'b011110110011;
   3381: result <= 12'b011110110011;
   3382: result <= 12'b011110110100;
   3383: result <= 12'b011110110100;
   3384: result <= 12'b011110110100;
   3385: result <= 12'b011110110100;
   3386: result <= 12'b011110110101;
   3387: result <= 12'b011110110101;
   3388: result <= 12'b011110110101;
   3389: result <= 12'b011110110101;
   3390: result <= 12'b011110110101;
   3391: result <= 12'b011110110110;
   3392: result <= 12'b011110110110;
   3393: result <= 12'b011110110110;
   3394: result <= 12'b011110110110;
   3395: result <= 12'b011110110110;
   3396: result <= 12'b011110110111;
   3397: result <= 12'b011110110111;
   3398: result <= 12'b011110110111;
   3399: result <= 12'b011110110111;
   3400: result <= 12'b011110110111;
   3401: result <= 12'b011110111000;
   3402: result <= 12'b011110111000;
   3403: result <= 12'b011110111000;
   3404: result <= 12'b011110111000;
   3405: result <= 12'b011110111001;
   3406: result <= 12'b011110111001;
   3407: result <= 12'b011110111001;
   3408: result <= 12'b011110111001;
   3409: result <= 12'b011110111001;
   3410: result <= 12'b011110111010;
   3411: result <= 12'b011110111010;
   3412: result <= 12'b011110111010;
   3413: result <= 12'b011110111010;
   3414: result <= 12'b011110111010;
   3415: result <= 12'b011110111011;
   3416: result <= 12'b011110111011;
   3417: result <= 12'b011110111011;
   3418: result <= 12'b011110111011;
   3419: result <= 12'b011110111011;
   3420: result <= 12'b011110111100;
   3421: result <= 12'b011110111100;
   3422: result <= 12'b011110111100;
   3423: result <= 12'b011110111100;
   3424: result <= 12'b011110111100;
   3425: result <= 12'b011110111101;
   3426: result <= 12'b011110111101;
   3427: result <= 12'b011110111101;
   3428: result <= 12'b011110111101;
   3429: result <= 12'b011110111101;
   3430: result <= 12'b011110111110;
   3431: result <= 12'b011110111110;
   3432: result <= 12'b011110111110;
   3433: result <= 12'b011110111110;
   3434: result <= 12'b011110111110;
   3435: result <= 12'b011110111111;
   3436: result <= 12'b011110111111;
   3437: result <= 12'b011110111111;
   3438: result <= 12'b011110111111;
   3439: result <= 12'b011110111111;
   3440: result <= 12'b011111000000;
   3441: result <= 12'b011111000000;
   3442: result <= 12'b011111000000;
   3443: result <= 12'b011111000000;
   3444: result <= 12'b011111000000;
   3445: result <= 12'b011111000001;
   3446: result <= 12'b011111000001;
   3447: result <= 12'b011111000001;
   3448: result <= 12'b011111000001;
   3449: result <= 12'b011111000001;
   3450: result <= 12'b011111000001;
   3451: result <= 12'b011111000010;
   3452: result <= 12'b011111000010;
   3453: result <= 12'b011111000010;
   3454: result <= 12'b011111000010;
   3455: result <= 12'b011111000010;
   3456: result <= 12'b011111000011;
   3457: result <= 12'b011111000011;
   3458: result <= 12'b011111000011;
   3459: result <= 12'b011111000011;
   3460: result <= 12'b011111000011;
   3461: result <= 12'b011111000100;
   3462: result <= 12'b011111000100;
   3463: result <= 12'b011111000100;
   3464: result <= 12'b011111000100;
   3465: result <= 12'b011111000100;
   3466: result <= 12'b011111000101;
   3467: result <= 12'b011111000101;
   3468: result <= 12'b011111000101;
   3469: result <= 12'b011111000101;
   3470: result <= 12'b011111000101;
   3471: result <= 12'b011111000101;
   3472: result <= 12'b011111000110;
   3473: result <= 12'b011111000110;
   3474: result <= 12'b011111000110;
   3475: result <= 12'b011111000110;
   3476: result <= 12'b011111000110;
   3477: result <= 12'b011111000111;
   3478: result <= 12'b011111000111;
   3479: result <= 12'b011111000111;
   3480: result <= 12'b011111000111;
   3481: result <= 12'b011111000111;
   3482: result <= 12'b011111000111;
   3483: result <= 12'b011111001000;
   3484: result <= 12'b011111001000;
   3485: result <= 12'b011111001000;
   3486: result <= 12'b011111001000;
   3487: result <= 12'b011111001000;
   3488: result <= 12'b011111001001;
   3489: result <= 12'b011111001001;
   3490: result <= 12'b011111001001;
   3491: result <= 12'b011111001001;
   3492: result <= 12'b011111001001;
   3493: result <= 12'b011111001001;
   3494: result <= 12'b011111001010;
   3495: result <= 12'b011111001010;
   3496: result <= 12'b011111001010;
   3497: result <= 12'b011111001010;
   3498: result <= 12'b011111001010;
   3499: result <= 12'b011111001011;
   3500: result <= 12'b011111001011;
   3501: result <= 12'b011111001011;
   3502: result <= 12'b011111001011;
   3503: result <= 12'b011111001011;
   3504: result <= 12'b011111001011;
   3505: result <= 12'b011111001100;
   3506: result <= 12'b011111001100;
   3507: result <= 12'b011111001100;
   3508: result <= 12'b011111001100;
   3509: result <= 12'b011111001100;
   3510: result <= 12'b011111001101;
   3511: result <= 12'b011111001101;
   3512: result <= 12'b011111001101;
   3513: result <= 12'b011111001101;
   3514: result <= 12'b011111001101;
   3515: result <= 12'b011111001101;
   3516: result <= 12'b011111001110;
   3517: result <= 12'b011111001110;
   3518: result <= 12'b011111001110;
   3519: result <= 12'b011111001110;
   3520: result <= 12'b011111001110;
   3521: result <= 12'b011111001110;
   3522: result <= 12'b011111001111;
   3523: result <= 12'b011111001111;
   3524: result <= 12'b011111001111;
   3525: result <= 12'b011111001111;
   3526: result <= 12'b011111001111;
   3527: result <= 12'b011111001111;
   3528: result <= 12'b011111010000;
   3529: result <= 12'b011111010000;
   3530: result <= 12'b011111010000;
   3531: result <= 12'b011111010000;
   3532: result <= 12'b011111010000;
   3533: result <= 12'b011111010000;
   3534: result <= 12'b011111010001;
   3535: result <= 12'b011111010001;
   3536: result <= 12'b011111010001;
   3537: result <= 12'b011111010001;
   3538: result <= 12'b011111010001;
   3539: result <= 12'b011111010001;
   3540: result <= 12'b011111010010;
   3541: result <= 12'b011111010010;
   3542: result <= 12'b011111010010;
   3543: result <= 12'b011111010010;
   3544: result <= 12'b011111010010;
   3545: result <= 12'b011111010010;
   3546: result <= 12'b011111010011;
   3547: result <= 12'b011111010011;
   3548: result <= 12'b011111010011;
   3549: result <= 12'b011111010011;
   3550: result <= 12'b011111010011;
   3551: result <= 12'b011111010011;
   3552: result <= 12'b011111010100;
   3553: result <= 12'b011111010100;
   3554: result <= 12'b011111010100;
   3555: result <= 12'b011111010100;
   3556: result <= 12'b011111010100;
   3557: result <= 12'b011111010100;
   3558: result <= 12'b011111010101;
   3559: result <= 12'b011111010101;
   3560: result <= 12'b011111010101;
   3561: result <= 12'b011111010101;
   3562: result <= 12'b011111010101;
   3563: result <= 12'b011111010101;
   3564: result <= 12'b011111010110;
   3565: result <= 12'b011111010110;
   3566: result <= 12'b011111010110;
   3567: result <= 12'b011111010110;
   3568: result <= 12'b011111010110;
   3569: result <= 12'b011111010110;
   3570: result <= 12'b011111010110;
   3571: result <= 12'b011111010111;
   3572: result <= 12'b011111010111;
   3573: result <= 12'b011111010111;
   3574: result <= 12'b011111010111;
   3575: result <= 12'b011111010111;
   3576: result <= 12'b011111010111;
   3577: result <= 12'b011111011000;
   3578: result <= 12'b011111011000;
   3579: result <= 12'b011111011000;
   3580: result <= 12'b011111011000;
   3581: result <= 12'b011111011000;
   3582: result <= 12'b011111011000;
   3583: result <= 12'b011111011000;
   3584: result <= 12'b011111011001;
   3585: result <= 12'b011111011001;
   3586: result <= 12'b011111011001;
   3587: result <= 12'b011111011001;
   3588: result <= 12'b011111011001;
   3589: result <= 12'b011111011001;
   3590: result <= 12'b011111011010;
   3591: result <= 12'b011111011010;
   3592: result <= 12'b011111011010;
   3593: result <= 12'b011111011010;
   3594: result <= 12'b011111011010;
   3595: result <= 12'b011111011010;
   3596: result <= 12'b011111011010;
   3597: result <= 12'b011111011011;
   3598: result <= 12'b011111011011;
   3599: result <= 12'b011111011011;
   3600: result <= 12'b011111011011;
   3601: result <= 12'b011111011011;
   3602: result <= 12'b011111011011;
   3603: result <= 12'b011111011100;
   3604: result <= 12'b011111011100;
   3605: result <= 12'b011111011100;
   3606: result <= 12'b011111011100;
   3607: result <= 12'b011111011100;
   3608: result <= 12'b011111011100;
   3609: result <= 12'b011111011100;
   3610: result <= 12'b011111011101;
   3611: result <= 12'b011111011101;
   3612: result <= 12'b011111011101;
   3613: result <= 12'b011111011101;
   3614: result <= 12'b011111011101;
   3615: result <= 12'b011111011101;
   3616: result <= 12'b011111011101;
   3617: result <= 12'b011111011110;
   3618: result <= 12'b011111011110;
   3619: result <= 12'b011111011110;
   3620: result <= 12'b011111011110;
   3621: result <= 12'b011111011110;
   3622: result <= 12'b011111011110;
   3623: result <= 12'b011111011110;
   3624: result <= 12'b011111011111;
   3625: result <= 12'b011111011111;
   3626: result <= 12'b011111011111;
   3627: result <= 12'b011111011111;
   3628: result <= 12'b011111011111;
   3629: result <= 12'b011111011111;
   3630: result <= 12'b011111011111;
   3631: result <= 12'b011111100000;
   3632: result <= 12'b011111100000;
   3633: result <= 12'b011111100000;
   3634: result <= 12'b011111100000;
   3635: result <= 12'b011111100000;
   3636: result <= 12'b011111100000;
   3637: result <= 12'b011111100000;
   3638: result <= 12'b011111100000;
   3639: result <= 12'b011111100001;
   3640: result <= 12'b011111100001;
   3641: result <= 12'b011111100001;
   3642: result <= 12'b011111100001;
   3643: result <= 12'b011111100001;
   3644: result <= 12'b011111100001;
   3645: result <= 12'b011111100001;
   3646: result <= 12'b011111100010;
   3647: result <= 12'b011111100010;
   3648: result <= 12'b011111100010;
   3649: result <= 12'b011111100010;
   3650: result <= 12'b011111100010;
   3651: result <= 12'b011111100010;
   3652: result <= 12'b011111100010;
   3653: result <= 12'b011111100011;
   3654: result <= 12'b011111100011;
   3655: result <= 12'b011111100011;
   3656: result <= 12'b011111100011;
   3657: result <= 12'b011111100011;
   3658: result <= 12'b011111100011;
   3659: result <= 12'b011111100011;
   3660: result <= 12'b011111100011;
   3661: result <= 12'b011111100100;
   3662: result <= 12'b011111100100;
   3663: result <= 12'b011111100100;
   3664: result <= 12'b011111100100;
   3665: result <= 12'b011111100100;
   3666: result <= 12'b011111100100;
   3667: result <= 12'b011111100100;
   3668: result <= 12'b011111100100;
   3669: result <= 12'b011111100101;
   3670: result <= 12'b011111100101;
   3671: result <= 12'b011111100101;
   3672: result <= 12'b011111100101;
   3673: result <= 12'b011111100101;
   3674: result <= 12'b011111100101;
   3675: result <= 12'b011111100101;
   3676: result <= 12'b011111100101;
   3677: result <= 12'b011111100110;
   3678: result <= 12'b011111100110;
   3679: result <= 12'b011111100110;
   3680: result <= 12'b011111100110;
   3681: result <= 12'b011111100110;
   3682: result <= 12'b011111100110;
   3683: result <= 12'b011111100110;
   3684: result <= 12'b011111100110;
   3685: result <= 12'b011111100111;
   3686: result <= 12'b011111100111;
   3687: result <= 12'b011111100111;
   3688: result <= 12'b011111100111;
   3689: result <= 12'b011111100111;
   3690: result <= 12'b011111100111;
   3691: result <= 12'b011111100111;
   3692: result <= 12'b011111100111;
   3693: result <= 12'b011111101000;
   3694: result <= 12'b011111101000;
   3695: result <= 12'b011111101000;
   3696: result <= 12'b011111101000;
   3697: result <= 12'b011111101000;
   3698: result <= 12'b011111101000;
   3699: result <= 12'b011111101000;
   3700: result <= 12'b011111101000;
   3701: result <= 12'b011111101001;
   3702: result <= 12'b011111101001;
   3703: result <= 12'b011111101001;
   3704: result <= 12'b011111101001;
   3705: result <= 12'b011111101001;
   3706: result <= 12'b011111101001;
   3707: result <= 12'b011111101001;
   3708: result <= 12'b011111101001;
   3709: result <= 12'b011111101001;
   3710: result <= 12'b011111101010;
   3711: result <= 12'b011111101010;
   3712: result <= 12'b011111101010;
   3713: result <= 12'b011111101010;
   3714: result <= 12'b011111101010;
   3715: result <= 12'b011111101010;
   3716: result <= 12'b011111101010;
   3717: result <= 12'b011111101010;
   3718: result <= 12'b011111101011;
   3719: result <= 12'b011111101011;
   3720: result <= 12'b011111101011;
   3721: result <= 12'b011111101011;
   3722: result <= 12'b011111101011;
   3723: result <= 12'b011111101011;
   3724: result <= 12'b011111101011;
   3725: result <= 12'b011111101011;
   3726: result <= 12'b011111101011;
   3727: result <= 12'b011111101100;
   3728: result <= 12'b011111101100;
   3729: result <= 12'b011111101100;
   3730: result <= 12'b011111101100;
   3731: result <= 12'b011111101100;
   3732: result <= 12'b011111101100;
   3733: result <= 12'b011111101100;
   3734: result <= 12'b011111101100;
   3735: result <= 12'b011111101100;
   3736: result <= 12'b011111101101;
   3737: result <= 12'b011111101101;
   3738: result <= 12'b011111101101;
   3739: result <= 12'b011111101101;
   3740: result <= 12'b011111101101;
   3741: result <= 12'b011111101101;
   3742: result <= 12'b011111101101;
   3743: result <= 12'b011111101101;
   3744: result <= 12'b011111101101;
   3745: result <= 12'b011111101101;
   3746: result <= 12'b011111101110;
   3747: result <= 12'b011111101110;
   3748: result <= 12'b011111101110;
   3749: result <= 12'b011111101110;
   3750: result <= 12'b011111101110;
   3751: result <= 12'b011111101110;
   3752: result <= 12'b011111101110;
   3753: result <= 12'b011111101110;
   3754: result <= 12'b011111101110;
   3755: result <= 12'b011111101111;
   3756: result <= 12'b011111101111;
   3757: result <= 12'b011111101111;
   3758: result <= 12'b011111101111;
   3759: result <= 12'b011111101111;
   3760: result <= 12'b011111101111;
   3761: result <= 12'b011111101111;
   3762: result <= 12'b011111101111;
   3763: result <= 12'b011111101111;
   3764: result <= 12'b011111101111;
   3765: result <= 12'b011111110000;
   3766: result <= 12'b011111110000;
   3767: result <= 12'b011111110000;
   3768: result <= 12'b011111110000;
   3769: result <= 12'b011111110000;
   3770: result <= 12'b011111110000;
   3771: result <= 12'b011111110000;
   3772: result <= 12'b011111110000;
   3773: result <= 12'b011111110000;
   3774: result <= 12'b011111110000;
   3775: result <= 12'b011111110001;
   3776: result <= 12'b011111110001;
   3777: result <= 12'b011111110001;
   3778: result <= 12'b011111110001;
   3779: result <= 12'b011111110001;
   3780: result <= 12'b011111110001;
   3781: result <= 12'b011111110001;
   3782: result <= 12'b011111110001;
   3783: result <= 12'b011111110001;
   3784: result <= 12'b011111110001;
   3785: result <= 12'b011111110001;
   3786: result <= 12'b011111110010;
   3787: result <= 12'b011111110010;
   3788: result <= 12'b011111110010;
   3789: result <= 12'b011111110010;
   3790: result <= 12'b011111110010;
   3791: result <= 12'b011111110010;
   3792: result <= 12'b011111110010;
   3793: result <= 12'b011111110010;
   3794: result <= 12'b011111110010;
   3795: result <= 12'b011111110010;
   3796: result <= 12'b011111110010;
   3797: result <= 12'b011111110011;
   3798: result <= 12'b011111110011;
   3799: result <= 12'b011111110011;
   3800: result <= 12'b011111110011;
   3801: result <= 12'b011111110011;
   3802: result <= 12'b011111110011;
   3803: result <= 12'b011111110011;
   3804: result <= 12'b011111110011;
   3805: result <= 12'b011111110011;
   3806: result <= 12'b011111110011;
   3807: result <= 12'b011111110011;
   3808: result <= 12'b011111110100;
   3809: result <= 12'b011111110100;
   3810: result <= 12'b011111110100;
   3811: result <= 12'b011111110100;
   3812: result <= 12'b011111110100;
   3813: result <= 12'b011111110100;
   3814: result <= 12'b011111110100;
   3815: result <= 12'b011111110100;
   3816: result <= 12'b011111110100;
   3817: result <= 12'b011111110100;
   3818: result <= 12'b011111110100;
   3819: result <= 12'b011111110100;
   3820: result <= 12'b011111110101;
   3821: result <= 12'b011111110101;
   3822: result <= 12'b011111110101;
   3823: result <= 12'b011111110101;
   3824: result <= 12'b011111110101;
   3825: result <= 12'b011111110101;
   3826: result <= 12'b011111110101;
   3827: result <= 12'b011111110101;
   3828: result <= 12'b011111110101;
   3829: result <= 12'b011111110101;
   3830: result <= 12'b011111110101;
   3831: result <= 12'b011111110101;
   3832: result <= 12'b011111110110;
   3833: result <= 12'b011111110110;
   3834: result <= 12'b011111110110;
   3835: result <= 12'b011111110110;
   3836: result <= 12'b011111110110;
   3837: result <= 12'b011111110110;
   3838: result <= 12'b011111110110;
   3839: result <= 12'b011111110110;
   3840: result <= 12'b011111110110;
   3841: result <= 12'b011111110110;
   3842: result <= 12'b011111110110;
   3843: result <= 12'b011111110110;
   3844: result <= 12'b011111110110;
   3845: result <= 12'b011111110111;
   3846: result <= 12'b011111110111;
   3847: result <= 12'b011111110111;
   3848: result <= 12'b011111110111;
   3849: result <= 12'b011111110111;
   3850: result <= 12'b011111110111;
   3851: result <= 12'b011111110111;
   3852: result <= 12'b011111110111;
   3853: result <= 12'b011111110111;
   3854: result <= 12'b011111110111;
   3855: result <= 12'b011111110111;
   3856: result <= 12'b011111110111;
   3857: result <= 12'b011111110111;
   3858: result <= 12'b011111110111;
   3859: result <= 12'b011111111000;
   3860: result <= 12'b011111111000;
   3861: result <= 12'b011111111000;
   3862: result <= 12'b011111111000;
   3863: result <= 12'b011111111000;
   3864: result <= 12'b011111111000;
   3865: result <= 12'b011111111000;
   3866: result <= 12'b011111111000;
   3867: result <= 12'b011111111000;
   3868: result <= 12'b011111111000;
   3869: result <= 12'b011111111000;
   3870: result <= 12'b011111111000;
   3871: result <= 12'b011111111000;
   3872: result <= 12'b011111111000;
   3873: result <= 12'b011111111001;
   3874: result <= 12'b011111111001;
   3875: result <= 12'b011111111001;
   3876: result <= 12'b011111111001;
   3877: result <= 12'b011111111001;
   3878: result <= 12'b011111111001;
   3879: result <= 12'b011111111001;
   3880: result <= 12'b011111111001;
   3881: result <= 12'b011111111001;
   3882: result <= 12'b011111111001;
   3883: result <= 12'b011111111001;
   3884: result <= 12'b011111111001;
   3885: result <= 12'b011111111001;
   3886: result <= 12'b011111111001;
   3887: result <= 12'b011111111001;
   3888: result <= 12'b011111111001;
   3889: result <= 12'b011111111010;
   3890: result <= 12'b011111111010;
   3891: result <= 12'b011111111010;
   3892: result <= 12'b011111111010;
   3893: result <= 12'b011111111010;
   3894: result <= 12'b011111111010;
   3895: result <= 12'b011111111010;
   3896: result <= 12'b011111111010;
   3897: result <= 12'b011111111010;
   3898: result <= 12'b011111111010;
   3899: result <= 12'b011111111010;
   3900: result <= 12'b011111111010;
   3901: result <= 12'b011111111010;
   3902: result <= 12'b011111111010;
   3903: result <= 12'b011111111010;
   3904: result <= 12'b011111111010;
   3905: result <= 12'b011111111011;
   3906: result <= 12'b011111111011;
   3907: result <= 12'b011111111011;
   3908: result <= 12'b011111111011;
   3909: result <= 12'b011111111011;
   3910: result <= 12'b011111111011;
   3911: result <= 12'b011111111011;
   3912: result <= 12'b011111111011;
   3913: result <= 12'b011111111011;
   3914: result <= 12'b011111111011;
   3915: result <= 12'b011111111011;
   3916: result <= 12'b011111111011;
   3917: result <= 12'b011111111011;
   3918: result <= 12'b011111111011;
   3919: result <= 12'b011111111011;
   3920: result <= 12'b011111111011;
   3921: result <= 12'b011111111011;
   3922: result <= 12'b011111111011;
   3923: result <= 12'b011111111011;
   3924: result <= 12'b011111111100;
   3925: result <= 12'b011111111100;
   3926: result <= 12'b011111111100;
   3927: result <= 12'b011111111100;
   3928: result <= 12'b011111111100;
   3929: result <= 12'b011111111100;
   3930: result <= 12'b011111111100;
   3931: result <= 12'b011111111100;
   3932: result <= 12'b011111111100;
   3933: result <= 12'b011111111100;
   3934: result <= 12'b011111111100;
   3935: result <= 12'b011111111100;
   3936: result <= 12'b011111111100;
   3937: result <= 12'b011111111100;
   3938: result <= 12'b011111111100;
   3939: result <= 12'b011111111100;
   3940: result <= 12'b011111111100;
   3941: result <= 12'b011111111100;
   3942: result <= 12'b011111111100;
   3943: result <= 12'b011111111100;
   3944: result <= 12'b011111111101;
   3945: result <= 12'b011111111101;
   3946: result <= 12'b011111111101;
   3947: result <= 12'b011111111101;
   3948: result <= 12'b011111111101;
   3949: result <= 12'b011111111101;
   3950: result <= 12'b011111111101;
   3951: result <= 12'b011111111101;
   3952: result <= 12'b011111111101;
   3953: result <= 12'b011111111101;
   3954: result <= 12'b011111111101;
   3955: result <= 12'b011111111101;
   3956: result <= 12'b011111111101;
   3957: result <= 12'b011111111101;
   3958: result <= 12'b011111111101;
   3959: result <= 12'b011111111101;
   3960: result <= 12'b011111111101;
   3961: result <= 12'b011111111101;
   3962: result <= 12'b011111111101;
   3963: result <= 12'b011111111101;
   3964: result <= 12'b011111111101;
   3965: result <= 12'b011111111101;
   3966: result <= 12'b011111111101;
   3967: result <= 12'b011111111101;
   3968: result <= 12'b011111111110;
   3969: result <= 12'b011111111110;
   3970: result <= 12'b011111111110;
   3971: result <= 12'b011111111110;
   3972: result <= 12'b011111111110;
   3973: result <= 12'b011111111110;
   3974: result <= 12'b011111111110;
   3975: result <= 12'b011111111110;
   3976: result <= 12'b011111111110;
   3977: result <= 12'b011111111110;
   3978: result <= 12'b011111111110;
   3979: result <= 12'b011111111110;
   3980: result <= 12'b011111111110;
   3981: result <= 12'b011111111110;
   3982: result <= 12'b011111111110;
   3983: result <= 12'b011111111110;
   3984: result <= 12'b011111111110;
   3985: result <= 12'b011111111110;
   3986: result <= 12'b011111111110;
   3987: result <= 12'b011111111110;
   3988: result <= 12'b011111111110;
   3989: result <= 12'b011111111110;
   3990: result <= 12'b011111111110;
   3991: result <= 12'b011111111110;
   3992: result <= 12'b011111111110;
   3993: result <= 12'b011111111110;
   3994: result <= 12'b011111111110;
   3995: result <= 12'b011111111110;
   3996: result <= 12'b011111111110;
   3997: result <= 12'b011111111111;
   3998: result <= 12'b011111111111;
   3999: result <= 12'b011111111111;
   4000: result <= 12'b011111111111;
   4001: result <= 12'b011111111111;
   4002: result <= 12'b011111111111;
   4003: result <= 12'b011111111111;
   4004: result <= 12'b011111111111;
   4005: result <= 12'b011111111111;
   4006: result <= 12'b011111111111;
   4007: result <= 12'b011111111111;
   4008: result <= 12'b011111111111;
   4009: result <= 12'b011111111111;
   4010: result <= 12'b011111111111;
   4011: result <= 12'b011111111111;
   4012: result <= 12'b011111111111;
   4013: result <= 12'b011111111111;
   4014: result <= 12'b011111111111;
   4015: result <= 12'b011111111111;
   4016: result <= 12'b011111111111;
   4017: result <= 12'b011111111111;
   4018: result <= 12'b011111111111;
   4019: result <= 12'b011111111111;
   4020: result <= 12'b011111111111;
   4021: result <= 12'b011111111111;
   4022: result <= 12'b011111111111;
   4023: result <= 12'b011111111111;
   4024: result <= 12'b011111111111;
   4025: result <= 12'b011111111111;
   4026: result <= 12'b011111111111;
   4027: result <= 12'b011111111111;
   4028: result <= 12'b011111111111;
   4029: result <= 12'b011111111111;
   4030: result <= 12'b011111111111;
   4031: result <= 12'b011111111111;
   4032: result <= 12'b011111111111;
   4033: result <= 12'b011111111111;
   4034: result <= 12'b011111111111;
   4035: result <= 12'b011111111111;
   4036: result <= 12'b011111111111;
   4037: result <= 12'b011111111111;
   4038: result <= 12'b011111111111;
   4039: result <= 12'b011111111111;
   4040: result <= 12'b011111111111;
   4041: result <= 12'b011111111111;
   4042: result <= 12'b011111111111;
   4043: result <= 12'b011111111111;
   4044: result <= 12'b011111111111;
   4045: result <= 12'b011111111111;
   4046: result <= 12'b011111111111;
   4047: result <= 12'b011111111111;
   4048: result <= 12'b011111111111;
   4049: result <= 12'b011111111111;
   4050: result <= 12'b011111111111;
   4051: result <= 12'b011111111111;
   4052: result <= 12'b011111111111;
   4053: result <= 12'b011111111111;
   4054: result <= 12'b011111111111;
   4055: result <= 12'b011111111111;
   4056: result <= 12'b011111111111;
   4057: result <= 12'b011111111111;
   4058: result <= 12'b011111111111;
   4059: result <= 12'b011111111111;
   4060: result <= 12'b011111111111;
   4061: result <= 12'b011111111111;
   4062: result <= 12'b011111111111;
   4063: result <= 12'b011111111111;
   4064: result <= 12'b011111111111;
   4065: result <= 12'b011111111111;
   4066: result <= 12'b011111111111;
   4067: result <= 12'b011111111111;
   4068: result <= 12'b011111111111;
   4069: result <= 12'b011111111111;
   4070: result <= 12'b011111111111;
   4071: result <= 12'b011111111111;
   4072: result <= 12'b011111111111;
   4073: result <= 12'b011111111111;
   4074: result <= 12'b011111111111;
   4075: result <= 12'b011111111111;
   4076: result <= 12'b011111111111;
   4077: result <= 12'b011111111111;
   4078: result <= 12'b011111111111;
   4079: result <= 12'b011111111111;
   4080: result <= 12'b011111111111;
   4081: result <= 12'b011111111111;
   4082: result <= 12'b011111111111;
   4083: result <= 12'b011111111111;
   4084: result <= 12'b011111111111;
   4085: result <= 12'b011111111111;
   4086: result <= 12'b011111111111;
   4087: result <= 12'b011111111111;
   4088: result <= 12'b011111111111;
   4089: result <= 12'b011111111111;
   4090: result <= 12'b011111111111;
   4091: result <= 12'b011111111111;
   4092: result <= 12'b011111111111;
   4093: result <= 12'b011111111111;
   4094: result <= 12'b011111111111;
   4095: result <= 12'b011111111111;
   4096: result <= 12'b011111111111;
   4097: result <= 12'b011111111111;
   4098: result <= 12'b011111111111;
   4099: result <= 12'b011111111111;
   4100: result <= 12'b011111111111;
   4101: result <= 12'b011111111111;
   4102: result <= 12'b011111111111;
   4103: result <= 12'b011111111111;
   4104: result <= 12'b011111111111;
   4105: result <= 12'b011111111111;
   4106: result <= 12'b011111111111;
   4107: result <= 12'b011111111111;
   4108: result <= 12'b011111111111;
   4109: result <= 12'b011111111111;
   4110: result <= 12'b011111111111;
   4111: result <= 12'b011111111111;
   4112: result <= 12'b011111111111;
   4113: result <= 12'b011111111111;
   4114: result <= 12'b011111111111;
   4115: result <= 12'b011111111111;
   4116: result <= 12'b011111111111;
   4117: result <= 12'b011111111111;
   4118: result <= 12'b011111111111;
   4119: result <= 12'b011111111111;
   4120: result <= 12'b011111111111;
   4121: result <= 12'b011111111111;
   4122: result <= 12'b011111111111;
   4123: result <= 12'b011111111111;
   4124: result <= 12'b011111111111;
   4125: result <= 12'b011111111111;
   4126: result <= 12'b011111111111;
   4127: result <= 12'b011111111111;
   4128: result <= 12'b011111111111;
   4129: result <= 12'b011111111111;
   4130: result <= 12'b011111111111;
   4131: result <= 12'b011111111111;
   4132: result <= 12'b011111111111;
   4133: result <= 12'b011111111111;
   4134: result <= 12'b011111111111;
   4135: result <= 12'b011111111111;
   4136: result <= 12'b011111111111;
   4137: result <= 12'b011111111111;
   4138: result <= 12'b011111111111;
   4139: result <= 12'b011111111111;
   4140: result <= 12'b011111111111;
   4141: result <= 12'b011111111111;
   4142: result <= 12'b011111111111;
   4143: result <= 12'b011111111111;
   4144: result <= 12'b011111111111;
   4145: result <= 12'b011111111111;
   4146: result <= 12'b011111111111;
   4147: result <= 12'b011111111111;
   4148: result <= 12'b011111111111;
   4149: result <= 12'b011111111111;
   4150: result <= 12'b011111111111;
   4151: result <= 12'b011111111111;
   4152: result <= 12'b011111111111;
   4153: result <= 12'b011111111111;
   4154: result <= 12'b011111111111;
   4155: result <= 12'b011111111111;
   4156: result <= 12'b011111111111;
   4157: result <= 12'b011111111111;
   4158: result <= 12'b011111111111;
   4159: result <= 12'b011111111111;
   4160: result <= 12'b011111111111;
   4161: result <= 12'b011111111111;
   4162: result <= 12'b011111111111;
   4163: result <= 12'b011111111111;
   4164: result <= 12'b011111111111;
   4165: result <= 12'b011111111111;
   4166: result <= 12'b011111111111;
   4167: result <= 12'b011111111111;
   4168: result <= 12'b011111111111;
   4169: result <= 12'b011111111111;
   4170: result <= 12'b011111111111;
   4171: result <= 12'b011111111111;
   4172: result <= 12'b011111111111;
   4173: result <= 12'b011111111111;
   4174: result <= 12'b011111111111;
   4175: result <= 12'b011111111111;
   4176: result <= 12'b011111111111;
   4177: result <= 12'b011111111111;
   4178: result <= 12'b011111111111;
   4179: result <= 12'b011111111111;
   4180: result <= 12'b011111111111;
   4181: result <= 12'b011111111111;
   4182: result <= 12'b011111111111;
   4183: result <= 12'b011111111111;
   4184: result <= 12'b011111111111;
   4185: result <= 12'b011111111111;
   4186: result <= 12'b011111111111;
   4187: result <= 12'b011111111111;
   4188: result <= 12'b011111111111;
   4189: result <= 12'b011111111111;
   4190: result <= 12'b011111111111;
   4191: result <= 12'b011111111111;
   4192: result <= 12'b011111111111;
   4193: result <= 12'b011111111111;
   4194: result <= 12'b011111111111;
   4195: result <= 12'b011111111111;
   4196: result <= 12'b011111111110;
   4197: result <= 12'b011111111110;
   4198: result <= 12'b011111111110;
   4199: result <= 12'b011111111110;
   4200: result <= 12'b011111111110;
   4201: result <= 12'b011111111110;
   4202: result <= 12'b011111111110;
   4203: result <= 12'b011111111110;
   4204: result <= 12'b011111111110;
   4205: result <= 12'b011111111110;
   4206: result <= 12'b011111111110;
   4207: result <= 12'b011111111110;
   4208: result <= 12'b011111111110;
   4209: result <= 12'b011111111110;
   4210: result <= 12'b011111111110;
   4211: result <= 12'b011111111110;
   4212: result <= 12'b011111111110;
   4213: result <= 12'b011111111110;
   4214: result <= 12'b011111111110;
   4215: result <= 12'b011111111110;
   4216: result <= 12'b011111111110;
   4217: result <= 12'b011111111110;
   4218: result <= 12'b011111111110;
   4219: result <= 12'b011111111110;
   4220: result <= 12'b011111111110;
   4221: result <= 12'b011111111110;
   4222: result <= 12'b011111111110;
   4223: result <= 12'b011111111110;
   4224: result <= 12'b011111111110;
   4225: result <= 12'b011111111101;
   4226: result <= 12'b011111111101;
   4227: result <= 12'b011111111101;
   4228: result <= 12'b011111111101;
   4229: result <= 12'b011111111101;
   4230: result <= 12'b011111111101;
   4231: result <= 12'b011111111101;
   4232: result <= 12'b011111111101;
   4233: result <= 12'b011111111101;
   4234: result <= 12'b011111111101;
   4235: result <= 12'b011111111101;
   4236: result <= 12'b011111111101;
   4237: result <= 12'b011111111101;
   4238: result <= 12'b011111111101;
   4239: result <= 12'b011111111101;
   4240: result <= 12'b011111111101;
   4241: result <= 12'b011111111101;
   4242: result <= 12'b011111111101;
   4243: result <= 12'b011111111101;
   4244: result <= 12'b011111111101;
   4245: result <= 12'b011111111101;
   4246: result <= 12'b011111111101;
   4247: result <= 12'b011111111101;
   4248: result <= 12'b011111111101;
   4249: result <= 12'b011111111100;
   4250: result <= 12'b011111111100;
   4251: result <= 12'b011111111100;
   4252: result <= 12'b011111111100;
   4253: result <= 12'b011111111100;
   4254: result <= 12'b011111111100;
   4255: result <= 12'b011111111100;
   4256: result <= 12'b011111111100;
   4257: result <= 12'b011111111100;
   4258: result <= 12'b011111111100;
   4259: result <= 12'b011111111100;
   4260: result <= 12'b011111111100;
   4261: result <= 12'b011111111100;
   4262: result <= 12'b011111111100;
   4263: result <= 12'b011111111100;
   4264: result <= 12'b011111111100;
   4265: result <= 12'b011111111100;
   4266: result <= 12'b011111111100;
   4267: result <= 12'b011111111100;
   4268: result <= 12'b011111111100;
   4269: result <= 12'b011111111011;
   4270: result <= 12'b011111111011;
   4271: result <= 12'b011111111011;
   4272: result <= 12'b011111111011;
   4273: result <= 12'b011111111011;
   4274: result <= 12'b011111111011;
   4275: result <= 12'b011111111011;
   4276: result <= 12'b011111111011;
   4277: result <= 12'b011111111011;
   4278: result <= 12'b011111111011;
   4279: result <= 12'b011111111011;
   4280: result <= 12'b011111111011;
   4281: result <= 12'b011111111011;
   4282: result <= 12'b011111111011;
   4283: result <= 12'b011111111011;
   4284: result <= 12'b011111111011;
   4285: result <= 12'b011111111011;
   4286: result <= 12'b011111111011;
   4287: result <= 12'b011111111011;
   4288: result <= 12'b011111111010;
   4289: result <= 12'b011111111010;
   4290: result <= 12'b011111111010;
   4291: result <= 12'b011111111010;
   4292: result <= 12'b011111111010;
   4293: result <= 12'b011111111010;
   4294: result <= 12'b011111111010;
   4295: result <= 12'b011111111010;
   4296: result <= 12'b011111111010;
   4297: result <= 12'b011111111010;
   4298: result <= 12'b011111111010;
   4299: result <= 12'b011111111010;
   4300: result <= 12'b011111111010;
   4301: result <= 12'b011111111010;
   4302: result <= 12'b011111111010;
   4303: result <= 12'b011111111010;
   4304: result <= 12'b011111111001;
   4305: result <= 12'b011111111001;
   4306: result <= 12'b011111111001;
   4307: result <= 12'b011111111001;
   4308: result <= 12'b011111111001;
   4309: result <= 12'b011111111001;
   4310: result <= 12'b011111111001;
   4311: result <= 12'b011111111001;
   4312: result <= 12'b011111111001;
   4313: result <= 12'b011111111001;
   4314: result <= 12'b011111111001;
   4315: result <= 12'b011111111001;
   4316: result <= 12'b011111111001;
   4317: result <= 12'b011111111001;
   4318: result <= 12'b011111111001;
   4319: result <= 12'b011111111001;
   4320: result <= 12'b011111111000;
   4321: result <= 12'b011111111000;
   4322: result <= 12'b011111111000;
   4323: result <= 12'b011111111000;
   4324: result <= 12'b011111111000;
   4325: result <= 12'b011111111000;
   4326: result <= 12'b011111111000;
   4327: result <= 12'b011111111000;
   4328: result <= 12'b011111111000;
   4329: result <= 12'b011111111000;
   4330: result <= 12'b011111111000;
   4331: result <= 12'b011111111000;
   4332: result <= 12'b011111111000;
   4333: result <= 12'b011111111000;
   4334: result <= 12'b011111110111;
   4335: result <= 12'b011111110111;
   4336: result <= 12'b011111110111;
   4337: result <= 12'b011111110111;
   4338: result <= 12'b011111110111;
   4339: result <= 12'b011111110111;
   4340: result <= 12'b011111110111;
   4341: result <= 12'b011111110111;
   4342: result <= 12'b011111110111;
   4343: result <= 12'b011111110111;
   4344: result <= 12'b011111110111;
   4345: result <= 12'b011111110111;
   4346: result <= 12'b011111110111;
   4347: result <= 12'b011111110111;
   4348: result <= 12'b011111110110;
   4349: result <= 12'b011111110110;
   4350: result <= 12'b011111110110;
   4351: result <= 12'b011111110110;
   4352: result <= 12'b011111110110;
   4353: result <= 12'b011111110110;
   4354: result <= 12'b011111110110;
   4355: result <= 12'b011111110110;
   4356: result <= 12'b011111110110;
   4357: result <= 12'b011111110110;
   4358: result <= 12'b011111110110;
   4359: result <= 12'b011111110110;
   4360: result <= 12'b011111110110;
   4361: result <= 12'b011111110101;
   4362: result <= 12'b011111110101;
   4363: result <= 12'b011111110101;
   4364: result <= 12'b011111110101;
   4365: result <= 12'b011111110101;
   4366: result <= 12'b011111110101;
   4367: result <= 12'b011111110101;
   4368: result <= 12'b011111110101;
   4369: result <= 12'b011111110101;
   4370: result <= 12'b011111110101;
   4371: result <= 12'b011111110101;
   4372: result <= 12'b011111110101;
   4373: result <= 12'b011111110100;
   4374: result <= 12'b011111110100;
   4375: result <= 12'b011111110100;
   4376: result <= 12'b011111110100;
   4377: result <= 12'b011111110100;
   4378: result <= 12'b011111110100;
   4379: result <= 12'b011111110100;
   4380: result <= 12'b011111110100;
   4381: result <= 12'b011111110100;
   4382: result <= 12'b011111110100;
   4383: result <= 12'b011111110100;
   4384: result <= 12'b011111110100;
   4385: result <= 12'b011111110011;
   4386: result <= 12'b011111110011;
   4387: result <= 12'b011111110011;
   4388: result <= 12'b011111110011;
   4389: result <= 12'b011111110011;
   4390: result <= 12'b011111110011;
   4391: result <= 12'b011111110011;
   4392: result <= 12'b011111110011;
   4393: result <= 12'b011111110011;
   4394: result <= 12'b011111110011;
   4395: result <= 12'b011111110011;
   4396: result <= 12'b011111110010;
   4397: result <= 12'b011111110010;
   4398: result <= 12'b011111110010;
   4399: result <= 12'b011111110010;
   4400: result <= 12'b011111110010;
   4401: result <= 12'b011111110010;
   4402: result <= 12'b011111110010;
   4403: result <= 12'b011111110010;
   4404: result <= 12'b011111110010;
   4405: result <= 12'b011111110010;
   4406: result <= 12'b011111110010;
   4407: result <= 12'b011111110001;
   4408: result <= 12'b011111110001;
   4409: result <= 12'b011111110001;
   4410: result <= 12'b011111110001;
   4411: result <= 12'b011111110001;
   4412: result <= 12'b011111110001;
   4413: result <= 12'b011111110001;
   4414: result <= 12'b011111110001;
   4415: result <= 12'b011111110001;
   4416: result <= 12'b011111110001;
   4417: result <= 12'b011111110001;
   4418: result <= 12'b011111110000;
   4419: result <= 12'b011111110000;
   4420: result <= 12'b011111110000;
   4421: result <= 12'b011111110000;
   4422: result <= 12'b011111110000;
   4423: result <= 12'b011111110000;
   4424: result <= 12'b011111110000;
   4425: result <= 12'b011111110000;
   4426: result <= 12'b011111110000;
   4427: result <= 12'b011111110000;
   4428: result <= 12'b011111101111;
   4429: result <= 12'b011111101111;
   4430: result <= 12'b011111101111;
   4431: result <= 12'b011111101111;
   4432: result <= 12'b011111101111;
   4433: result <= 12'b011111101111;
   4434: result <= 12'b011111101111;
   4435: result <= 12'b011111101111;
   4436: result <= 12'b011111101111;
   4437: result <= 12'b011111101111;
   4438: result <= 12'b011111101110;
   4439: result <= 12'b011111101110;
   4440: result <= 12'b011111101110;
   4441: result <= 12'b011111101110;
   4442: result <= 12'b011111101110;
   4443: result <= 12'b011111101110;
   4444: result <= 12'b011111101110;
   4445: result <= 12'b011111101110;
   4446: result <= 12'b011111101110;
   4447: result <= 12'b011111101101;
   4448: result <= 12'b011111101101;
   4449: result <= 12'b011111101101;
   4450: result <= 12'b011111101101;
   4451: result <= 12'b011111101101;
   4452: result <= 12'b011111101101;
   4453: result <= 12'b011111101101;
   4454: result <= 12'b011111101101;
   4455: result <= 12'b011111101101;
   4456: result <= 12'b011111101101;
   4457: result <= 12'b011111101100;
   4458: result <= 12'b011111101100;
   4459: result <= 12'b011111101100;
   4460: result <= 12'b011111101100;
   4461: result <= 12'b011111101100;
   4462: result <= 12'b011111101100;
   4463: result <= 12'b011111101100;
   4464: result <= 12'b011111101100;
   4465: result <= 12'b011111101100;
   4466: result <= 12'b011111101011;
   4467: result <= 12'b011111101011;
   4468: result <= 12'b011111101011;
   4469: result <= 12'b011111101011;
   4470: result <= 12'b011111101011;
   4471: result <= 12'b011111101011;
   4472: result <= 12'b011111101011;
   4473: result <= 12'b011111101011;
   4474: result <= 12'b011111101011;
   4475: result <= 12'b011111101010;
   4476: result <= 12'b011111101010;
   4477: result <= 12'b011111101010;
   4478: result <= 12'b011111101010;
   4479: result <= 12'b011111101010;
   4480: result <= 12'b011111101010;
   4481: result <= 12'b011111101010;
   4482: result <= 12'b011111101010;
   4483: result <= 12'b011111101001;
   4484: result <= 12'b011111101001;
   4485: result <= 12'b011111101001;
   4486: result <= 12'b011111101001;
   4487: result <= 12'b011111101001;
   4488: result <= 12'b011111101001;
   4489: result <= 12'b011111101001;
   4490: result <= 12'b011111101001;
   4491: result <= 12'b011111101001;
   4492: result <= 12'b011111101000;
   4493: result <= 12'b011111101000;
   4494: result <= 12'b011111101000;
   4495: result <= 12'b011111101000;
   4496: result <= 12'b011111101000;
   4497: result <= 12'b011111101000;
   4498: result <= 12'b011111101000;
   4499: result <= 12'b011111101000;
   4500: result <= 12'b011111100111;
   4501: result <= 12'b011111100111;
   4502: result <= 12'b011111100111;
   4503: result <= 12'b011111100111;
   4504: result <= 12'b011111100111;
   4505: result <= 12'b011111100111;
   4506: result <= 12'b011111100111;
   4507: result <= 12'b011111100111;
   4508: result <= 12'b011111100110;
   4509: result <= 12'b011111100110;
   4510: result <= 12'b011111100110;
   4511: result <= 12'b011111100110;
   4512: result <= 12'b011111100110;
   4513: result <= 12'b011111100110;
   4514: result <= 12'b011111100110;
   4515: result <= 12'b011111100110;
   4516: result <= 12'b011111100101;
   4517: result <= 12'b011111100101;
   4518: result <= 12'b011111100101;
   4519: result <= 12'b011111100101;
   4520: result <= 12'b011111100101;
   4521: result <= 12'b011111100101;
   4522: result <= 12'b011111100101;
   4523: result <= 12'b011111100101;
   4524: result <= 12'b011111100100;
   4525: result <= 12'b011111100100;
   4526: result <= 12'b011111100100;
   4527: result <= 12'b011111100100;
   4528: result <= 12'b011111100100;
   4529: result <= 12'b011111100100;
   4530: result <= 12'b011111100100;
   4531: result <= 12'b011111100100;
   4532: result <= 12'b011111100011;
   4533: result <= 12'b011111100011;
   4534: result <= 12'b011111100011;
   4535: result <= 12'b011111100011;
   4536: result <= 12'b011111100011;
   4537: result <= 12'b011111100011;
   4538: result <= 12'b011111100011;
   4539: result <= 12'b011111100011;
   4540: result <= 12'b011111100010;
   4541: result <= 12'b011111100010;
   4542: result <= 12'b011111100010;
   4543: result <= 12'b011111100010;
   4544: result <= 12'b011111100010;
   4545: result <= 12'b011111100010;
   4546: result <= 12'b011111100010;
   4547: result <= 12'b011111100001;
   4548: result <= 12'b011111100001;
   4549: result <= 12'b011111100001;
   4550: result <= 12'b011111100001;
   4551: result <= 12'b011111100001;
   4552: result <= 12'b011111100001;
   4553: result <= 12'b011111100001;
   4554: result <= 12'b011111100000;
   4555: result <= 12'b011111100000;
   4556: result <= 12'b011111100000;
   4557: result <= 12'b011111100000;
   4558: result <= 12'b011111100000;
   4559: result <= 12'b011111100000;
   4560: result <= 12'b011111100000;
   4561: result <= 12'b011111100000;
   4562: result <= 12'b011111011111;
   4563: result <= 12'b011111011111;
   4564: result <= 12'b011111011111;
   4565: result <= 12'b011111011111;
   4566: result <= 12'b011111011111;
   4567: result <= 12'b011111011111;
   4568: result <= 12'b011111011111;
   4569: result <= 12'b011111011110;
   4570: result <= 12'b011111011110;
   4571: result <= 12'b011111011110;
   4572: result <= 12'b011111011110;
   4573: result <= 12'b011111011110;
   4574: result <= 12'b011111011110;
   4575: result <= 12'b011111011110;
   4576: result <= 12'b011111011101;
   4577: result <= 12'b011111011101;
   4578: result <= 12'b011111011101;
   4579: result <= 12'b011111011101;
   4580: result <= 12'b011111011101;
   4581: result <= 12'b011111011101;
   4582: result <= 12'b011111011101;
   4583: result <= 12'b011111011100;
   4584: result <= 12'b011111011100;
   4585: result <= 12'b011111011100;
   4586: result <= 12'b011111011100;
   4587: result <= 12'b011111011100;
   4588: result <= 12'b011111011100;
   4589: result <= 12'b011111011100;
   4590: result <= 12'b011111011011;
   4591: result <= 12'b011111011011;
   4592: result <= 12'b011111011011;
   4593: result <= 12'b011111011011;
   4594: result <= 12'b011111011011;
   4595: result <= 12'b011111011011;
   4596: result <= 12'b011111011010;
   4597: result <= 12'b011111011010;
   4598: result <= 12'b011111011010;
   4599: result <= 12'b011111011010;
   4600: result <= 12'b011111011010;
   4601: result <= 12'b011111011010;
   4602: result <= 12'b011111011010;
   4603: result <= 12'b011111011001;
   4604: result <= 12'b011111011001;
   4605: result <= 12'b011111011001;
   4606: result <= 12'b011111011001;
   4607: result <= 12'b011111011001;
   4608: result <= 12'b011111011001;
   4609: result <= 12'b011111011000;
   4610: result <= 12'b011111011000;
   4611: result <= 12'b011111011000;
   4612: result <= 12'b011111011000;
   4613: result <= 12'b011111011000;
   4614: result <= 12'b011111011000;
   4615: result <= 12'b011111011000;
   4616: result <= 12'b011111010111;
   4617: result <= 12'b011111010111;
   4618: result <= 12'b011111010111;
   4619: result <= 12'b011111010111;
   4620: result <= 12'b011111010111;
   4621: result <= 12'b011111010111;
   4622: result <= 12'b011111010110;
   4623: result <= 12'b011111010110;
   4624: result <= 12'b011111010110;
   4625: result <= 12'b011111010110;
   4626: result <= 12'b011111010110;
   4627: result <= 12'b011111010110;
   4628: result <= 12'b011111010110;
   4629: result <= 12'b011111010101;
   4630: result <= 12'b011111010101;
   4631: result <= 12'b011111010101;
   4632: result <= 12'b011111010101;
   4633: result <= 12'b011111010101;
   4634: result <= 12'b011111010101;
   4635: result <= 12'b011111010100;
   4636: result <= 12'b011111010100;
   4637: result <= 12'b011111010100;
   4638: result <= 12'b011111010100;
   4639: result <= 12'b011111010100;
   4640: result <= 12'b011111010100;
   4641: result <= 12'b011111010011;
   4642: result <= 12'b011111010011;
   4643: result <= 12'b011111010011;
   4644: result <= 12'b011111010011;
   4645: result <= 12'b011111010011;
   4646: result <= 12'b011111010011;
   4647: result <= 12'b011111010010;
   4648: result <= 12'b011111010010;
   4649: result <= 12'b011111010010;
   4650: result <= 12'b011111010010;
   4651: result <= 12'b011111010010;
   4652: result <= 12'b011111010010;
   4653: result <= 12'b011111010001;
   4654: result <= 12'b011111010001;
   4655: result <= 12'b011111010001;
   4656: result <= 12'b011111010001;
   4657: result <= 12'b011111010001;
   4658: result <= 12'b011111010001;
   4659: result <= 12'b011111010000;
   4660: result <= 12'b011111010000;
   4661: result <= 12'b011111010000;
   4662: result <= 12'b011111010000;
   4663: result <= 12'b011111010000;
   4664: result <= 12'b011111010000;
   4665: result <= 12'b011111001111;
   4666: result <= 12'b011111001111;
   4667: result <= 12'b011111001111;
   4668: result <= 12'b011111001111;
   4669: result <= 12'b011111001111;
   4670: result <= 12'b011111001111;
   4671: result <= 12'b011111001110;
   4672: result <= 12'b011111001110;
   4673: result <= 12'b011111001110;
   4674: result <= 12'b011111001110;
   4675: result <= 12'b011111001110;
   4676: result <= 12'b011111001110;
   4677: result <= 12'b011111001101;
   4678: result <= 12'b011111001101;
   4679: result <= 12'b011111001101;
   4680: result <= 12'b011111001101;
   4681: result <= 12'b011111001101;
   4682: result <= 12'b011111001101;
   4683: result <= 12'b011111001100;
   4684: result <= 12'b011111001100;
   4685: result <= 12'b011111001100;
   4686: result <= 12'b011111001100;
   4687: result <= 12'b011111001100;
   4688: result <= 12'b011111001011;
   4689: result <= 12'b011111001011;
   4690: result <= 12'b011111001011;
   4691: result <= 12'b011111001011;
   4692: result <= 12'b011111001011;
   4693: result <= 12'b011111001011;
   4694: result <= 12'b011111001010;
   4695: result <= 12'b011111001010;
   4696: result <= 12'b011111001010;
   4697: result <= 12'b011111001010;
   4698: result <= 12'b011111001010;
   4699: result <= 12'b011111001001;
   4700: result <= 12'b011111001001;
   4701: result <= 12'b011111001001;
   4702: result <= 12'b011111001001;
   4703: result <= 12'b011111001001;
   4704: result <= 12'b011111001001;
   4705: result <= 12'b011111001000;
   4706: result <= 12'b011111001000;
   4707: result <= 12'b011111001000;
   4708: result <= 12'b011111001000;
   4709: result <= 12'b011111001000;
   4710: result <= 12'b011111000111;
   4711: result <= 12'b011111000111;
   4712: result <= 12'b011111000111;
   4713: result <= 12'b011111000111;
   4714: result <= 12'b011111000111;
   4715: result <= 12'b011111000111;
   4716: result <= 12'b011111000110;
   4717: result <= 12'b011111000110;
   4718: result <= 12'b011111000110;
   4719: result <= 12'b011111000110;
   4720: result <= 12'b011111000110;
   4721: result <= 12'b011111000101;
   4722: result <= 12'b011111000101;
   4723: result <= 12'b011111000101;
   4724: result <= 12'b011111000101;
   4725: result <= 12'b011111000101;
   4726: result <= 12'b011111000101;
   4727: result <= 12'b011111000100;
   4728: result <= 12'b011111000100;
   4729: result <= 12'b011111000100;
   4730: result <= 12'b011111000100;
   4731: result <= 12'b011111000100;
   4732: result <= 12'b011111000011;
   4733: result <= 12'b011111000011;
   4734: result <= 12'b011111000011;
   4735: result <= 12'b011111000011;
   4736: result <= 12'b011111000011;
   4737: result <= 12'b011111000010;
   4738: result <= 12'b011111000010;
   4739: result <= 12'b011111000010;
   4740: result <= 12'b011111000010;
   4741: result <= 12'b011111000010;
   4742: result <= 12'b011111000001;
   4743: result <= 12'b011111000001;
   4744: result <= 12'b011111000001;
   4745: result <= 12'b011111000001;
   4746: result <= 12'b011111000001;
   4747: result <= 12'b011111000001;
   4748: result <= 12'b011111000000;
   4749: result <= 12'b011111000000;
   4750: result <= 12'b011111000000;
   4751: result <= 12'b011111000000;
   4752: result <= 12'b011111000000;
   4753: result <= 12'b011110111111;
   4754: result <= 12'b011110111111;
   4755: result <= 12'b011110111111;
   4756: result <= 12'b011110111111;
   4757: result <= 12'b011110111111;
   4758: result <= 12'b011110111110;
   4759: result <= 12'b011110111110;
   4760: result <= 12'b011110111110;
   4761: result <= 12'b011110111110;
   4762: result <= 12'b011110111110;
   4763: result <= 12'b011110111101;
   4764: result <= 12'b011110111101;
   4765: result <= 12'b011110111101;
   4766: result <= 12'b011110111101;
   4767: result <= 12'b011110111101;
   4768: result <= 12'b011110111100;
   4769: result <= 12'b011110111100;
   4770: result <= 12'b011110111100;
   4771: result <= 12'b011110111100;
   4772: result <= 12'b011110111100;
   4773: result <= 12'b011110111011;
   4774: result <= 12'b011110111011;
   4775: result <= 12'b011110111011;
   4776: result <= 12'b011110111011;
   4777: result <= 12'b011110111011;
   4778: result <= 12'b011110111010;
   4779: result <= 12'b011110111010;
   4780: result <= 12'b011110111010;
   4781: result <= 12'b011110111010;
   4782: result <= 12'b011110111010;
   4783: result <= 12'b011110111001;
   4784: result <= 12'b011110111001;
   4785: result <= 12'b011110111001;
   4786: result <= 12'b011110111001;
   4787: result <= 12'b011110111001;
   4788: result <= 12'b011110111000;
   4789: result <= 12'b011110111000;
   4790: result <= 12'b011110111000;
   4791: result <= 12'b011110111000;
   4792: result <= 12'b011110110111;
   4793: result <= 12'b011110110111;
   4794: result <= 12'b011110110111;
   4795: result <= 12'b011110110111;
   4796: result <= 12'b011110110111;
   4797: result <= 12'b011110110110;
   4798: result <= 12'b011110110110;
   4799: result <= 12'b011110110110;
   4800: result <= 12'b011110110110;
   4801: result <= 12'b011110110110;
   4802: result <= 12'b011110110101;
   4803: result <= 12'b011110110101;
   4804: result <= 12'b011110110101;
   4805: result <= 12'b011110110101;
   4806: result <= 12'b011110110101;
   4807: result <= 12'b011110110100;
   4808: result <= 12'b011110110100;
   4809: result <= 12'b011110110100;
   4810: result <= 12'b011110110100;
   4811: result <= 12'b011110110011;
   4812: result <= 12'b011110110011;
   4813: result <= 12'b011110110011;
   4814: result <= 12'b011110110011;
   4815: result <= 12'b011110110011;
   4816: result <= 12'b011110110010;
   4817: result <= 12'b011110110010;
   4818: result <= 12'b011110110010;
   4819: result <= 12'b011110110010;
   4820: result <= 12'b011110110010;
   4821: result <= 12'b011110110001;
   4822: result <= 12'b011110110001;
   4823: result <= 12'b011110110001;
   4824: result <= 12'b011110110001;
   4825: result <= 12'b011110110000;
   4826: result <= 12'b011110110000;
   4827: result <= 12'b011110110000;
   4828: result <= 12'b011110110000;
   4829: result <= 12'b011110110000;
   4830: result <= 12'b011110101111;
   4831: result <= 12'b011110101111;
   4832: result <= 12'b011110101111;
   4833: result <= 12'b011110101111;
   4834: result <= 12'b011110101111;
   4835: result <= 12'b011110101110;
   4836: result <= 12'b011110101110;
   4837: result <= 12'b011110101110;
   4838: result <= 12'b011110101110;
   4839: result <= 12'b011110101101;
   4840: result <= 12'b011110101101;
   4841: result <= 12'b011110101101;
   4842: result <= 12'b011110101101;
   4843: result <= 12'b011110101101;
   4844: result <= 12'b011110101100;
   4845: result <= 12'b011110101100;
   4846: result <= 12'b011110101100;
   4847: result <= 12'b011110101100;
   4848: result <= 12'b011110101011;
   4849: result <= 12'b011110101011;
   4850: result <= 12'b011110101011;
   4851: result <= 12'b011110101011;
   4852: result <= 12'b011110101011;
   4853: result <= 12'b011110101010;
   4854: result <= 12'b011110101010;
   4855: result <= 12'b011110101010;
   4856: result <= 12'b011110101010;
   4857: result <= 12'b011110101001;
   4858: result <= 12'b011110101001;
   4859: result <= 12'b011110101001;
   4860: result <= 12'b011110101001;
   4861: result <= 12'b011110101000;
   4862: result <= 12'b011110101000;
   4863: result <= 12'b011110101000;
   4864: result <= 12'b011110101000;
   4865: result <= 12'b011110101000;
   4866: result <= 12'b011110100111;
   4867: result <= 12'b011110100111;
   4868: result <= 12'b011110100111;
   4869: result <= 12'b011110100111;
   4870: result <= 12'b011110100110;
   4871: result <= 12'b011110100110;
   4872: result <= 12'b011110100110;
   4873: result <= 12'b011110100110;
   4874: result <= 12'b011110100110;
   4875: result <= 12'b011110100101;
   4876: result <= 12'b011110100101;
   4877: result <= 12'b011110100101;
   4878: result <= 12'b011110100101;
   4879: result <= 12'b011110100100;
   4880: result <= 12'b011110100100;
   4881: result <= 12'b011110100100;
   4882: result <= 12'b011110100100;
   4883: result <= 12'b011110100011;
   4884: result <= 12'b011110100011;
   4885: result <= 12'b011110100011;
   4886: result <= 12'b011110100011;
   4887: result <= 12'b011110100010;
   4888: result <= 12'b011110100010;
   4889: result <= 12'b011110100010;
   4890: result <= 12'b011110100010;
   4891: result <= 12'b011110100010;
   4892: result <= 12'b011110100001;
   4893: result <= 12'b011110100001;
   4894: result <= 12'b011110100001;
   4895: result <= 12'b011110100001;
   4896: result <= 12'b011110100000;
   4897: result <= 12'b011110100000;
   4898: result <= 12'b011110100000;
   4899: result <= 12'b011110100000;
   4900: result <= 12'b011110011111;
   4901: result <= 12'b011110011111;
   4902: result <= 12'b011110011111;
   4903: result <= 12'b011110011111;
   4904: result <= 12'b011110011110;
   4905: result <= 12'b011110011110;
   4906: result <= 12'b011110011110;
   4907: result <= 12'b011110011110;
   4908: result <= 12'b011110011110;
   4909: result <= 12'b011110011101;
   4910: result <= 12'b011110011101;
   4911: result <= 12'b011110011101;
   4912: result <= 12'b011110011101;
   4913: result <= 12'b011110011100;
   4914: result <= 12'b011110011100;
   4915: result <= 12'b011110011100;
   4916: result <= 12'b011110011100;
   4917: result <= 12'b011110011011;
   4918: result <= 12'b011110011011;
   4919: result <= 12'b011110011011;
   4920: result <= 12'b011110011011;
   4921: result <= 12'b011110011010;
   4922: result <= 12'b011110011010;
   4923: result <= 12'b011110011010;
   4924: result <= 12'b011110011010;
   4925: result <= 12'b011110011001;
   4926: result <= 12'b011110011001;
   4927: result <= 12'b011110011001;
   4928: result <= 12'b011110011001;
   4929: result <= 12'b011110011000;
   4930: result <= 12'b011110011000;
   4931: result <= 12'b011110011000;
   4932: result <= 12'b011110011000;
   4933: result <= 12'b011110010111;
   4934: result <= 12'b011110010111;
   4935: result <= 12'b011110010111;
   4936: result <= 12'b011110010111;
   4937: result <= 12'b011110010110;
   4938: result <= 12'b011110010110;
   4939: result <= 12'b011110010110;
   4940: result <= 12'b011110010110;
   4941: result <= 12'b011110010101;
   4942: result <= 12'b011110010101;
   4943: result <= 12'b011110010101;
   4944: result <= 12'b011110010101;
   4945: result <= 12'b011110010100;
   4946: result <= 12'b011110010100;
   4947: result <= 12'b011110010100;
   4948: result <= 12'b011110010100;
   4949: result <= 12'b011110010011;
   4950: result <= 12'b011110010011;
   4951: result <= 12'b011110010011;
   4952: result <= 12'b011110010011;
   4953: result <= 12'b011110010010;
   4954: result <= 12'b011110010010;
   4955: result <= 12'b011110010010;
   4956: result <= 12'b011110010010;
   4957: result <= 12'b011110010001;
   4958: result <= 12'b011110010001;
   4959: result <= 12'b011110010001;
   4960: result <= 12'b011110010001;
   4961: result <= 12'b011110010000;
   4962: result <= 12'b011110010000;
   4963: result <= 12'b011110010000;
   4964: result <= 12'b011110010000;
   4965: result <= 12'b011110001111;
   4966: result <= 12'b011110001111;
   4967: result <= 12'b011110001111;
   4968: result <= 12'b011110001111;
   4969: result <= 12'b011110001110;
   4970: result <= 12'b011110001110;
   4971: result <= 12'b011110001110;
   4972: result <= 12'b011110001110;
   4973: result <= 12'b011110001101;
   4974: result <= 12'b011110001101;
   4975: result <= 12'b011110001101;
   4976: result <= 12'b011110001100;
   4977: result <= 12'b011110001100;
   4978: result <= 12'b011110001100;
   4979: result <= 12'b011110001100;
   4980: result <= 12'b011110001011;
   4981: result <= 12'b011110001011;
   4982: result <= 12'b011110001011;
   4983: result <= 12'b011110001011;
   4984: result <= 12'b011110001010;
   4985: result <= 12'b011110001010;
   4986: result <= 12'b011110001010;
   4987: result <= 12'b011110001010;
   4988: result <= 12'b011110001001;
   4989: result <= 12'b011110001001;
   4990: result <= 12'b011110001001;
   4991: result <= 12'b011110001001;
   4992: result <= 12'b011110001000;
   4993: result <= 12'b011110001000;
   4994: result <= 12'b011110001000;
   4995: result <= 12'b011110000111;
   4996: result <= 12'b011110000111;
   4997: result <= 12'b011110000111;
   4998: result <= 12'b011110000111;
   4999: result <= 12'b011110000110;
   5000: result <= 12'b011110000110;
   5001: result <= 12'b011110000110;
   5002: result <= 12'b011110000110;
   5003: result <= 12'b011110000101;
   5004: result <= 12'b011110000101;
   5005: result <= 12'b011110000101;
   5006: result <= 12'b011110000101;
   5007: result <= 12'b011110000100;
   5008: result <= 12'b011110000100;
   5009: result <= 12'b011110000100;
   5010: result <= 12'b011110000011;
   5011: result <= 12'b011110000011;
   5012: result <= 12'b011110000011;
   5013: result <= 12'b011110000011;
   5014: result <= 12'b011110000010;
   5015: result <= 12'b011110000010;
   5016: result <= 12'b011110000010;
   5017: result <= 12'b011110000010;
   5018: result <= 12'b011110000001;
   5019: result <= 12'b011110000001;
   5020: result <= 12'b011110000001;
   5021: result <= 12'b011110000000;
   5022: result <= 12'b011110000000;
   5023: result <= 12'b011110000000;
   5024: result <= 12'b011110000000;
   5025: result <= 12'b011101111111;
   5026: result <= 12'b011101111111;
   5027: result <= 12'b011101111111;
   5028: result <= 12'b011101111111;
   5029: result <= 12'b011101111110;
   5030: result <= 12'b011101111110;
   5031: result <= 12'b011101111110;
   5032: result <= 12'b011101111101;
   5033: result <= 12'b011101111101;
   5034: result <= 12'b011101111101;
   5035: result <= 12'b011101111101;
   5036: result <= 12'b011101111100;
   5037: result <= 12'b011101111100;
   5038: result <= 12'b011101111100;
   5039: result <= 12'b011101111100;
   5040: result <= 12'b011101111011;
   5041: result <= 12'b011101111011;
   5042: result <= 12'b011101111011;
   5043: result <= 12'b011101111010;
   5044: result <= 12'b011101111010;
   5045: result <= 12'b011101111010;
   5046: result <= 12'b011101111010;
   5047: result <= 12'b011101111001;
   5048: result <= 12'b011101111001;
   5049: result <= 12'b011101111001;
   5050: result <= 12'b011101111000;
   5051: result <= 12'b011101111000;
   5052: result <= 12'b011101111000;
   5053: result <= 12'b011101111000;
   5054: result <= 12'b011101110111;
   5055: result <= 12'b011101110111;
   5056: result <= 12'b011101110111;
   5057: result <= 12'b011101110110;
   5058: result <= 12'b011101110110;
   5059: result <= 12'b011101110110;
   5060: result <= 12'b011101110110;
   5061: result <= 12'b011101110101;
   5062: result <= 12'b011101110101;
   5063: result <= 12'b011101110101;
   5064: result <= 12'b011101110100;
   5065: result <= 12'b011101110100;
   5066: result <= 12'b011101110100;
   5067: result <= 12'b011101110100;
   5068: result <= 12'b011101110011;
   5069: result <= 12'b011101110011;
   5070: result <= 12'b011101110011;
   5071: result <= 12'b011101110010;
   5072: result <= 12'b011101110010;
   5073: result <= 12'b011101110010;
   5074: result <= 12'b011101110010;
   5075: result <= 12'b011101110001;
   5076: result <= 12'b011101110001;
   5077: result <= 12'b011101110001;
   5078: result <= 12'b011101110000;
   5079: result <= 12'b011101110000;
   5080: result <= 12'b011101110000;
   5081: result <= 12'b011101110000;
   5082: result <= 12'b011101101111;
   5083: result <= 12'b011101101111;
   5084: result <= 12'b011101101111;
   5085: result <= 12'b011101101110;
   5086: result <= 12'b011101101110;
   5087: result <= 12'b011101101110;
   5088: result <= 12'b011101101110;
   5089: result <= 12'b011101101101;
   5090: result <= 12'b011101101101;
   5091: result <= 12'b011101101101;
   5092: result <= 12'b011101101100;
   5093: result <= 12'b011101101100;
   5094: result <= 12'b011101101100;
   5095: result <= 12'b011101101100;
   5096: result <= 12'b011101101011;
   5097: result <= 12'b011101101011;
   5098: result <= 12'b011101101011;
   5099: result <= 12'b011101101010;
   5100: result <= 12'b011101101010;
   5101: result <= 12'b011101101010;
   5102: result <= 12'b011101101001;
   5103: result <= 12'b011101101001;
   5104: result <= 12'b011101101001;
   5105: result <= 12'b011101101001;
   5106: result <= 12'b011101101000;
   5107: result <= 12'b011101101000;
   5108: result <= 12'b011101101000;
   5109: result <= 12'b011101100111;
   5110: result <= 12'b011101100111;
   5111: result <= 12'b011101100111;
   5112: result <= 12'b011101100111;
   5113: result <= 12'b011101100110;
   5114: result <= 12'b011101100110;
   5115: result <= 12'b011101100110;
   5116: result <= 12'b011101100101;
   5117: result <= 12'b011101100101;
   5118: result <= 12'b011101100101;
   5119: result <= 12'b011101100100;
   5120: result <= 12'b011101100100;
   5121: result <= 12'b011101100100;
   5122: result <= 12'b011101100100;
   5123: result <= 12'b011101100011;
   5124: result <= 12'b011101100011;
   5125: result <= 12'b011101100011;
   5126: result <= 12'b011101100010;
   5127: result <= 12'b011101100010;
   5128: result <= 12'b011101100010;
   5129: result <= 12'b011101100001;
   5130: result <= 12'b011101100001;
   5131: result <= 12'b011101100001;
   5132: result <= 12'b011101100000;
   5133: result <= 12'b011101100000;
   5134: result <= 12'b011101100000;
   5135: result <= 12'b011101100000;
   5136: result <= 12'b011101011111;
   5137: result <= 12'b011101011111;
   5138: result <= 12'b011101011111;
   5139: result <= 12'b011101011110;
   5140: result <= 12'b011101011110;
   5141: result <= 12'b011101011110;
   5142: result <= 12'b011101011101;
   5143: result <= 12'b011101011101;
   5144: result <= 12'b011101011101;
   5145: result <= 12'b011101011101;
   5146: result <= 12'b011101011100;
   5147: result <= 12'b011101011100;
   5148: result <= 12'b011101011100;
   5149: result <= 12'b011101011011;
   5150: result <= 12'b011101011011;
   5151: result <= 12'b011101011011;
   5152: result <= 12'b011101011010;
   5153: result <= 12'b011101011010;
   5154: result <= 12'b011101011010;
   5155: result <= 12'b011101011001;
   5156: result <= 12'b011101011001;
   5157: result <= 12'b011101011001;
   5158: result <= 12'b011101011000;
   5159: result <= 12'b011101011000;
   5160: result <= 12'b011101011000;
   5161: result <= 12'b011101011000;
   5162: result <= 12'b011101010111;
   5163: result <= 12'b011101010111;
   5164: result <= 12'b011101010111;
   5165: result <= 12'b011101010110;
   5166: result <= 12'b011101010110;
   5167: result <= 12'b011101010110;
   5168: result <= 12'b011101010101;
   5169: result <= 12'b011101010101;
   5170: result <= 12'b011101010101;
   5171: result <= 12'b011101010100;
   5172: result <= 12'b011101010100;
   5173: result <= 12'b011101010100;
   5174: result <= 12'b011101010011;
   5175: result <= 12'b011101010011;
   5176: result <= 12'b011101010011;
   5177: result <= 12'b011101010011;
   5178: result <= 12'b011101010010;
   5179: result <= 12'b011101010010;
   5180: result <= 12'b011101010010;
   5181: result <= 12'b011101010001;
   5182: result <= 12'b011101010001;
   5183: result <= 12'b011101010001;
   5184: result <= 12'b011101010000;
   5185: result <= 12'b011101010000;
   5186: result <= 12'b011101010000;
   5187: result <= 12'b011101001111;
   5188: result <= 12'b011101001111;
   5189: result <= 12'b011101001111;
   5190: result <= 12'b011101001110;
   5191: result <= 12'b011101001110;
   5192: result <= 12'b011101001110;
   5193: result <= 12'b011101001101;
   5194: result <= 12'b011101001101;
   5195: result <= 12'b011101001101;
   5196: result <= 12'b011101001100;
   5197: result <= 12'b011101001100;
   5198: result <= 12'b011101001100;
   5199: result <= 12'b011101001011;
   5200: result <= 12'b011101001011;
   5201: result <= 12'b011101001011;
   5202: result <= 12'b011101001011;
   5203: result <= 12'b011101001010;
   5204: result <= 12'b011101001010;
   5205: result <= 12'b011101001010;
   5206: result <= 12'b011101001001;
   5207: result <= 12'b011101001001;
   5208: result <= 12'b011101001001;
   5209: result <= 12'b011101001000;
   5210: result <= 12'b011101001000;
   5211: result <= 12'b011101001000;
   5212: result <= 12'b011101000111;
   5213: result <= 12'b011101000111;
   5214: result <= 12'b011101000111;
   5215: result <= 12'b011101000110;
   5216: result <= 12'b011101000110;
   5217: result <= 12'b011101000110;
   5218: result <= 12'b011101000101;
   5219: result <= 12'b011101000101;
   5220: result <= 12'b011101000101;
   5221: result <= 12'b011101000100;
   5222: result <= 12'b011101000100;
   5223: result <= 12'b011101000100;
   5224: result <= 12'b011101000011;
   5225: result <= 12'b011101000011;
   5226: result <= 12'b011101000011;
   5227: result <= 12'b011101000010;
   5228: result <= 12'b011101000010;
   5229: result <= 12'b011101000010;
   5230: result <= 12'b011101000001;
   5231: result <= 12'b011101000001;
   5232: result <= 12'b011101000001;
   5233: result <= 12'b011101000000;
   5234: result <= 12'b011101000000;
   5235: result <= 12'b011101000000;
   5236: result <= 12'b011100111111;
   5237: result <= 12'b011100111111;
   5238: result <= 12'b011100111111;
   5239: result <= 12'b011100111110;
   5240: result <= 12'b011100111110;
   5241: result <= 12'b011100111110;
   5242: result <= 12'b011100111101;
   5243: result <= 12'b011100111101;
   5244: result <= 12'b011100111101;
   5245: result <= 12'b011100111100;
   5246: result <= 12'b011100111100;
   5247: result <= 12'b011100111100;
   5248: result <= 12'b011100111011;
   5249: result <= 12'b011100111011;
   5250: result <= 12'b011100111011;
   5251: result <= 12'b011100111010;
   5252: result <= 12'b011100111010;
   5253: result <= 12'b011100111010;
   5254: result <= 12'b011100111001;
   5255: result <= 12'b011100111001;
   5256: result <= 12'b011100111001;
   5257: result <= 12'b011100111000;
   5258: result <= 12'b011100111000;
   5259: result <= 12'b011100111000;
   5260: result <= 12'b011100110111;
   5261: result <= 12'b011100110111;
   5262: result <= 12'b011100110111;
   5263: result <= 12'b011100110110;
   5264: result <= 12'b011100110110;
   5265: result <= 12'b011100110110;
   5266: result <= 12'b011100110101;
   5267: result <= 12'b011100110101;
   5268: result <= 12'b011100110101;
   5269: result <= 12'b011100110100;
   5270: result <= 12'b011100110100;
   5271: result <= 12'b011100110100;
   5272: result <= 12'b011100110011;
   5273: result <= 12'b011100110011;
   5274: result <= 12'b011100110011;
   5275: result <= 12'b011100110010;
   5276: result <= 12'b011100110010;
   5277: result <= 12'b011100110010;
   5278: result <= 12'b011100110001;
   5279: result <= 12'b011100110001;
   5280: result <= 12'b011100110000;
   5281: result <= 12'b011100110000;
   5282: result <= 12'b011100110000;
   5283: result <= 12'b011100101111;
   5284: result <= 12'b011100101111;
   5285: result <= 12'b011100101111;
   5286: result <= 12'b011100101110;
   5287: result <= 12'b011100101110;
   5288: result <= 12'b011100101110;
   5289: result <= 12'b011100101101;
   5290: result <= 12'b011100101101;
   5291: result <= 12'b011100101101;
   5292: result <= 12'b011100101100;
   5293: result <= 12'b011100101100;
   5294: result <= 12'b011100101100;
   5295: result <= 12'b011100101011;
   5296: result <= 12'b011100101011;
   5297: result <= 12'b011100101011;
   5298: result <= 12'b011100101010;
   5299: result <= 12'b011100101010;
   5300: result <= 12'b011100101010;
   5301: result <= 12'b011100101001;
   5302: result <= 12'b011100101001;
   5303: result <= 12'b011100101000;
   5304: result <= 12'b011100101000;
   5305: result <= 12'b011100101000;
   5306: result <= 12'b011100100111;
   5307: result <= 12'b011100100111;
   5308: result <= 12'b011100100111;
   5309: result <= 12'b011100100110;
   5310: result <= 12'b011100100110;
   5311: result <= 12'b011100100110;
   5312: result <= 12'b011100100101;
   5313: result <= 12'b011100100101;
   5314: result <= 12'b011100100101;
   5315: result <= 12'b011100100100;
   5316: result <= 12'b011100100100;
   5317: result <= 12'b011100100100;
   5318: result <= 12'b011100100011;
   5319: result <= 12'b011100100011;
   5320: result <= 12'b011100100010;
   5321: result <= 12'b011100100010;
   5322: result <= 12'b011100100010;
   5323: result <= 12'b011100100001;
   5324: result <= 12'b011100100001;
   5325: result <= 12'b011100100001;
   5326: result <= 12'b011100100000;
   5327: result <= 12'b011100100000;
   5328: result <= 12'b011100100000;
   5329: result <= 12'b011100011111;
   5330: result <= 12'b011100011111;
   5331: result <= 12'b011100011111;
   5332: result <= 12'b011100011110;
   5333: result <= 12'b011100011110;
   5334: result <= 12'b011100011101;
   5335: result <= 12'b011100011101;
   5336: result <= 12'b011100011101;
   5337: result <= 12'b011100011100;
   5338: result <= 12'b011100011100;
   5339: result <= 12'b011100011100;
   5340: result <= 12'b011100011011;
   5341: result <= 12'b011100011011;
   5342: result <= 12'b011100011011;
   5343: result <= 12'b011100011010;
   5344: result <= 12'b011100011010;
   5345: result <= 12'b011100011010;
   5346: result <= 12'b011100011001;
   5347: result <= 12'b011100011001;
   5348: result <= 12'b011100011000;
   5349: result <= 12'b011100011000;
   5350: result <= 12'b011100011000;
   5351: result <= 12'b011100010111;
   5352: result <= 12'b011100010111;
   5353: result <= 12'b011100010111;
   5354: result <= 12'b011100010110;
   5355: result <= 12'b011100010110;
   5356: result <= 12'b011100010110;
   5357: result <= 12'b011100010101;
   5358: result <= 12'b011100010101;
   5359: result <= 12'b011100010100;
   5360: result <= 12'b011100010100;
   5361: result <= 12'b011100010100;
   5362: result <= 12'b011100010011;
   5363: result <= 12'b011100010011;
   5364: result <= 12'b011100010011;
   5365: result <= 12'b011100010010;
   5366: result <= 12'b011100010010;
   5367: result <= 12'b011100010001;
   5368: result <= 12'b011100010001;
   5369: result <= 12'b011100010001;
   5370: result <= 12'b011100010000;
   5371: result <= 12'b011100010000;
   5372: result <= 12'b011100010000;
   5373: result <= 12'b011100001111;
   5374: result <= 12'b011100001111;
   5375: result <= 12'b011100001111;
   5376: result <= 12'b011100001110;
   5377: result <= 12'b011100001110;
   5378: result <= 12'b011100001101;
   5379: result <= 12'b011100001101;
   5380: result <= 12'b011100001101;
   5381: result <= 12'b011100001100;
   5382: result <= 12'b011100001100;
   5383: result <= 12'b011100001100;
   5384: result <= 12'b011100001011;
   5385: result <= 12'b011100001011;
   5386: result <= 12'b011100001010;
   5387: result <= 12'b011100001010;
   5388: result <= 12'b011100001010;
   5389: result <= 12'b011100001001;
   5390: result <= 12'b011100001001;
   5391: result <= 12'b011100001001;
   5392: result <= 12'b011100001000;
   5393: result <= 12'b011100001000;
   5394: result <= 12'b011100000111;
   5395: result <= 12'b011100000111;
   5396: result <= 12'b011100000111;
   5397: result <= 12'b011100000110;
   5398: result <= 12'b011100000110;
   5399: result <= 12'b011100000110;
   5400: result <= 12'b011100000101;
   5401: result <= 12'b011100000101;
   5402: result <= 12'b011100000100;
   5403: result <= 12'b011100000100;
   5404: result <= 12'b011100000100;
   5405: result <= 12'b011100000011;
   5406: result <= 12'b011100000011;
   5407: result <= 12'b011100000011;
   5408: result <= 12'b011100000010;
   5409: result <= 12'b011100000010;
   5410: result <= 12'b011100000001;
   5411: result <= 12'b011100000001;
   5412: result <= 12'b011100000001;
   5413: result <= 12'b011100000000;
   5414: result <= 12'b011100000000;
   5415: result <= 12'b011100000000;
   5416: result <= 12'b011011111111;
   5417: result <= 12'b011011111111;
   5418: result <= 12'b011011111110;
   5419: result <= 12'b011011111110;
   5420: result <= 12'b011011111110;
   5421: result <= 12'b011011111101;
   5422: result <= 12'b011011111101;
   5423: result <= 12'b011011111100;
   5424: result <= 12'b011011111100;
   5425: result <= 12'b011011111100;
   5426: result <= 12'b011011111011;
   5427: result <= 12'b011011111011;
   5428: result <= 12'b011011111011;
   5429: result <= 12'b011011111010;
   5430: result <= 12'b011011111010;
   5431: result <= 12'b011011111001;
   5432: result <= 12'b011011111001;
   5433: result <= 12'b011011111001;
   5434: result <= 12'b011011111000;
   5435: result <= 12'b011011111000;
   5436: result <= 12'b011011110111;
   5437: result <= 12'b011011110111;
   5438: result <= 12'b011011110111;
   5439: result <= 12'b011011110110;
   5440: result <= 12'b011011110110;
   5441: result <= 12'b011011110110;
   5442: result <= 12'b011011110101;
   5443: result <= 12'b011011110101;
   5444: result <= 12'b011011110100;
   5445: result <= 12'b011011110100;
   5446: result <= 12'b011011110100;
   5447: result <= 12'b011011110011;
   5448: result <= 12'b011011110011;
   5449: result <= 12'b011011110010;
   5450: result <= 12'b011011110010;
   5451: result <= 12'b011011110010;
   5452: result <= 12'b011011110001;
   5453: result <= 12'b011011110001;
   5454: result <= 12'b011011110000;
   5455: result <= 12'b011011110000;
   5456: result <= 12'b011011110000;
   5457: result <= 12'b011011101111;
   5458: result <= 12'b011011101111;
   5459: result <= 12'b011011101111;
   5460: result <= 12'b011011101110;
   5461: result <= 12'b011011101110;
   5462: result <= 12'b011011101101;
   5463: result <= 12'b011011101101;
   5464: result <= 12'b011011101101;
   5465: result <= 12'b011011101100;
   5466: result <= 12'b011011101100;
   5467: result <= 12'b011011101011;
   5468: result <= 12'b011011101011;
   5469: result <= 12'b011011101011;
   5470: result <= 12'b011011101010;
   5471: result <= 12'b011011101010;
   5472: result <= 12'b011011101001;
   5473: result <= 12'b011011101001;
   5474: result <= 12'b011011101001;
   5475: result <= 12'b011011101000;
   5476: result <= 12'b011011101000;
   5477: result <= 12'b011011100111;
   5478: result <= 12'b011011100111;
   5479: result <= 12'b011011100111;
   5480: result <= 12'b011011100110;
   5481: result <= 12'b011011100110;
   5482: result <= 12'b011011100101;
   5483: result <= 12'b011011100101;
   5484: result <= 12'b011011100101;
   5485: result <= 12'b011011100100;
   5486: result <= 12'b011011100100;
   5487: result <= 12'b011011100011;
   5488: result <= 12'b011011100011;
   5489: result <= 12'b011011100011;
   5490: result <= 12'b011011100010;
   5491: result <= 12'b011011100010;
   5492: result <= 12'b011011100001;
   5493: result <= 12'b011011100001;
   5494: result <= 12'b011011100001;
   5495: result <= 12'b011011100000;
   5496: result <= 12'b011011100000;
   5497: result <= 12'b011011011111;
   5498: result <= 12'b011011011111;
   5499: result <= 12'b011011011111;
   5500: result <= 12'b011011011110;
   5501: result <= 12'b011011011110;
   5502: result <= 12'b011011011101;
   5503: result <= 12'b011011011101;
   5504: result <= 12'b011011011101;
   5505: result <= 12'b011011011100;
   5506: result <= 12'b011011011100;
   5507: result <= 12'b011011011011;
   5508: result <= 12'b011011011011;
   5509: result <= 12'b011011011011;
   5510: result <= 12'b011011011010;
   5511: result <= 12'b011011011010;
   5512: result <= 12'b011011011001;
   5513: result <= 12'b011011011001;
   5514: result <= 12'b011011011001;
   5515: result <= 12'b011011011000;
   5516: result <= 12'b011011011000;
   5517: result <= 12'b011011010111;
   5518: result <= 12'b011011010111;
   5519: result <= 12'b011011010111;
   5520: result <= 12'b011011010110;
   5521: result <= 12'b011011010110;
   5522: result <= 12'b011011010101;
   5523: result <= 12'b011011010101;
   5524: result <= 12'b011011010101;
   5525: result <= 12'b011011010100;
   5526: result <= 12'b011011010100;
   5527: result <= 12'b011011010011;
   5528: result <= 12'b011011010011;
   5529: result <= 12'b011011010010;
   5530: result <= 12'b011011010010;
   5531: result <= 12'b011011010010;
   5532: result <= 12'b011011010001;
   5533: result <= 12'b011011010001;
   5534: result <= 12'b011011010000;
   5535: result <= 12'b011011010000;
   5536: result <= 12'b011011010000;
   5537: result <= 12'b011011001111;
   5538: result <= 12'b011011001111;
   5539: result <= 12'b011011001110;
   5540: result <= 12'b011011001110;
   5541: result <= 12'b011011001110;
   5542: result <= 12'b011011001101;
   5543: result <= 12'b011011001101;
   5544: result <= 12'b011011001100;
   5545: result <= 12'b011011001100;
   5546: result <= 12'b011011001011;
   5547: result <= 12'b011011001011;
   5548: result <= 12'b011011001011;
   5549: result <= 12'b011011001010;
   5550: result <= 12'b011011001010;
   5551: result <= 12'b011011001001;
   5552: result <= 12'b011011001001;
   5553: result <= 12'b011011001001;
   5554: result <= 12'b011011001000;
   5555: result <= 12'b011011001000;
   5556: result <= 12'b011011000111;
   5557: result <= 12'b011011000111;
   5558: result <= 12'b011011000110;
   5559: result <= 12'b011011000110;
   5560: result <= 12'b011011000110;
   5561: result <= 12'b011011000101;
   5562: result <= 12'b011011000101;
   5563: result <= 12'b011011000100;
   5564: result <= 12'b011011000100;
   5565: result <= 12'b011011000100;
   5566: result <= 12'b011011000011;
   5567: result <= 12'b011011000011;
   5568: result <= 12'b011011000010;
   5569: result <= 12'b011011000010;
   5570: result <= 12'b011011000001;
   5571: result <= 12'b011011000001;
   5572: result <= 12'b011011000001;
   5573: result <= 12'b011011000000;
   5574: result <= 12'b011011000000;
   5575: result <= 12'b011010111111;
   5576: result <= 12'b011010111111;
   5577: result <= 12'b011010111110;
   5578: result <= 12'b011010111110;
   5579: result <= 12'b011010111110;
   5580: result <= 12'b011010111101;
   5581: result <= 12'b011010111101;
   5582: result <= 12'b011010111100;
   5583: result <= 12'b011010111100;
   5584: result <= 12'b011010111100;
   5585: result <= 12'b011010111011;
   5586: result <= 12'b011010111011;
   5587: result <= 12'b011010111010;
   5588: result <= 12'b011010111010;
   5589: result <= 12'b011010111001;
   5590: result <= 12'b011010111001;
   5591: result <= 12'b011010111001;
   5592: result <= 12'b011010111000;
   5593: result <= 12'b011010111000;
   5594: result <= 12'b011010110111;
   5595: result <= 12'b011010110111;
   5596: result <= 12'b011010110110;
   5597: result <= 12'b011010110110;
   5598: result <= 12'b011010110110;
   5599: result <= 12'b011010110101;
   5600: result <= 12'b011010110101;
   5601: result <= 12'b011010110100;
   5602: result <= 12'b011010110100;
   5603: result <= 12'b011010110011;
   5604: result <= 12'b011010110011;
   5605: result <= 12'b011010110011;
   5606: result <= 12'b011010110010;
   5607: result <= 12'b011010110010;
   5608: result <= 12'b011010110001;
   5609: result <= 12'b011010110001;
   5610: result <= 12'b011010110000;
   5611: result <= 12'b011010110000;
   5612: result <= 12'b011010110000;
   5613: result <= 12'b011010101111;
   5614: result <= 12'b011010101111;
   5615: result <= 12'b011010101110;
   5616: result <= 12'b011010101110;
   5617: result <= 12'b011010101101;
   5618: result <= 12'b011010101101;
   5619: result <= 12'b011010101101;
   5620: result <= 12'b011010101100;
   5621: result <= 12'b011010101100;
   5622: result <= 12'b011010101011;
   5623: result <= 12'b011010101011;
   5624: result <= 12'b011010101010;
   5625: result <= 12'b011010101010;
   5626: result <= 12'b011010101001;
   5627: result <= 12'b011010101001;
   5628: result <= 12'b011010101001;
   5629: result <= 12'b011010101000;
   5630: result <= 12'b011010101000;
   5631: result <= 12'b011010100111;
   5632: result <= 12'b011010100111;
   5633: result <= 12'b011010100110;
   5634: result <= 12'b011010100110;
   5635: result <= 12'b011010100110;
   5636: result <= 12'b011010100101;
   5637: result <= 12'b011010100101;
   5638: result <= 12'b011010100100;
   5639: result <= 12'b011010100100;
   5640: result <= 12'b011010100011;
   5641: result <= 12'b011010100011;
   5642: result <= 12'b011010100010;
   5643: result <= 12'b011010100010;
   5644: result <= 12'b011010100010;
   5645: result <= 12'b011010100001;
   5646: result <= 12'b011010100001;
   5647: result <= 12'b011010100000;
   5648: result <= 12'b011010100000;
   5649: result <= 12'b011010011111;
   5650: result <= 12'b011010011111;
   5651: result <= 12'b011010011111;
   5652: result <= 12'b011010011110;
   5653: result <= 12'b011010011110;
   5654: result <= 12'b011010011101;
   5655: result <= 12'b011010011101;
   5656: result <= 12'b011010011100;
   5657: result <= 12'b011010011100;
   5658: result <= 12'b011010011011;
   5659: result <= 12'b011010011011;
   5660: result <= 12'b011010011011;
   5661: result <= 12'b011010011010;
   5662: result <= 12'b011010011010;
   5663: result <= 12'b011010011001;
   5664: result <= 12'b011010011001;
   5665: result <= 12'b011010011000;
   5666: result <= 12'b011010011000;
   5667: result <= 12'b011010010111;
   5668: result <= 12'b011010010111;
   5669: result <= 12'b011010010111;
   5670: result <= 12'b011010010110;
   5671: result <= 12'b011010010110;
   5672: result <= 12'b011010010101;
   5673: result <= 12'b011010010101;
   5674: result <= 12'b011010010100;
   5675: result <= 12'b011010010100;
   5676: result <= 12'b011010010011;
   5677: result <= 12'b011010010011;
   5678: result <= 12'b011010010011;
   5679: result <= 12'b011010010010;
   5680: result <= 12'b011010010010;
   5681: result <= 12'b011010010001;
   5682: result <= 12'b011010010001;
   5683: result <= 12'b011010010000;
   5684: result <= 12'b011010010000;
   5685: result <= 12'b011010001111;
   5686: result <= 12'b011010001111;
   5687: result <= 12'b011010001110;
   5688: result <= 12'b011010001110;
   5689: result <= 12'b011010001110;
   5690: result <= 12'b011010001101;
   5691: result <= 12'b011010001101;
   5692: result <= 12'b011010001100;
   5693: result <= 12'b011010001100;
   5694: result <= 12'b011010001011;
   5695: result <= 12'b011010001011;
   5696: result <= 12'b011010001010;
   5697: result <= 12'b011010001010;
   5698: result <= 12'b011010001010;
   5699: result <= 12'b011010001001;
   5700: result <= 12'b011010001001;
   5701: result <= 12'b011010001000;
   5702: result <= 12'b011010001000;
   5703: result <= 12'b011010000111;
   5704: result <= 12'b011010000111;
   5705: result <= 12'b011010000110;
   5706: result <= 12'b011010000110;
   5707: result <= 12'b011010000101;
   5708: result <= 12'b011010000101;
   5709: result <= 12'b011010000101;
   5710: result <= 12'b011010000100;
   5711: result <= 12'b011010000100;
   5712: result <= 12'b011010000011;
   5713: result <= 12'b011010000011;
   5714: result <= 12'b011010000010;
   5715: result <= 12'b011010000010;
   5716: result <= 12'b011010000001;
   5717: result <= 12'b011010000001;
   5718: result <= 12'b011010000000;
   5719: result <= 12'b011010000000;
   5720: result <= 12'b011001111111;
   5721: result <= 12'b011001111111;
   5722: result <= 12'b011001111111;
   5723: result <= 12'b011001111110;
   5724: result <= 12'b011001111110;
   5725: result <= 12'b011001111101;
   5726: result <= 12'b011001111101;
   5727: result <= 12'b011001111100;
   5728: result <= 12'b011001111100;
   5729: result <= 12'b011001111011;
   5730: result <= 12'b011001111011;
   5731: result <= 12'b011001111010;
   5732: result <= 12'b011001111010;
   5733: result <= 12'b011001111010;
   5734: result <= 12'b011001111001;
   5735: result <= 12'b011001111001;
   5736: result <= 12'b011001111000;
   5737: result <= 12'b011001111000;
   5738: result <= 12'b011001110111;
   5739: result <= 12'b011001110111;
   5740: result <= 12'b011001110110;
   5741: result <= 12'b011001110110;
   5742: result <= 12'b011001110101;
   5743: result <= 12'b011001110101;
   5744: result <= 12'b011001110100;
   5745: result <= 12'b011001110100;
   5746: result <= 12'b011001110011;
   5747: result <= 12'b011001110011;
   5748: result <= 12'b011001110011;
   5749: result <= 12'b011001110010;
   5750: result <= 12'b011001110010;
   5751: result <= 12'b011001110001;
   5752: result <= 12'b011001110001;
   5753: result <= 12'b011001110000;
   5754: result <= 12'b011001110000;
   5755: result <= 12'b011001101111;
   5756: result <= 12'b011001101111;
   5757: result <= 12'b011001101110;
   5758: result <= 12'b011001101110;
   5759: result <= 12'b011001101101;
   5760: result <= 12'b011001101101;
   5761: result <= 12'b011001101101;
   5762: result <= 12'b011001101100;
   5763: result <= 12'b011001101100;
   5764: result <= 12'b011001101011;
   5765: result <= 12'b011001101011;
   5766: result <= 12'b011001101010;
   5767: result <= 12'b011001101010;
   5768: result <= 12'b011001101001;
   5769: result <= 12'b011001101001;
   5770: result <= 12'b011001101000;
   5771: result <= 12'b011001101000;
   5772: result <= 12'b011001100111;
   5773: result <= 12'b011001100111;
   5774: result <= 12'b011001100110;
   5775: result <= 12'b011001100110;
   5776: result <= 12'b011001100101;
   5777: result <= 12'b011001100101;
   5778: result <= 12'b011001100101;
   5779: result <= 12'b011001100100;
   5780: result <= 12'b011001100100;
   5781: result <= 12'b011001100011;
   5782: result <= 12'b011001100011;
   5783: result <= 12'b011001100010;
   5784: result <= 12'b011001100010;
   5785: result <= 12'b011001100001;
   5786: result <= 12'b011001100001;
   5787: result <= 12'b011001100000;
   5788: result <= 12'b011001100000;
   5789: result <= 12'b011001011111;
   5790: result <= 12'b011001011111;
   5791: result <= 12'b011001011110;
   5792: result <= 12'b011001011110;
   5793: result <= 12'b011001011101;
   5794: result <= 12'b011001011101;
   5795: result <= 12'b011001011100;
   5796: result <= 12'b011001011100;
   5797: result <= 12'b011001011011;
   5798: result <= 12'b011001011011;
   5799: result <= 12'b011001011011;
   5800: result <= 12'b011001011010;
   5801: result <= 12'b011001011010;
   5802: result <= 12'b011001011001;
   5803: result <= 12'b011001011001;
   5804: result <= 12'b011001011000;
   5805: result <= 12'b011001011000;
   5806: result <= 12'b011001010111;
   5807: result <= 12'b011001010111;
   5808: result <= 12'b011001010110;
   5809: result <= 12'b011001010110;
   5810: result <= 12'b011001010101;
   5811: result <= 12'b011001010101;
   5812: result <= 12'b011001010100;
   5813: result <= 12'b011001010100;
   5814: result <= 12'b011001010011;
   5815: result <= 12'b011001010011;
   5816: result <= 12'b011001010010;
   5817: result <= 12'b011001010010;
   5818: result <= 12'b011001010001;
   5819: result <= 12'b011001010001;
   5820: result <= 12'b011001010000;
   5821: result <= 12'b011001010000;
   5822: result <= 12'b011001001111;
   5823: result <= 12'b011001001111;
   5824: result <= 12'b011001001111;
   5825: result <= 12'b011001001110;
   5826: result <= 12'b011001001110;
   5827: result <= 12'b011001001101;
   5828: result <= 12'b011001001101;
   5829: result <= 12'b011001001100;
   5830: result <= 12'b011001001100;
   5831: result <= 12'b011001001011;
   5832: result <= 12'b011001001011;
   5833: result <= 12'b011001001010;
   5834: result <= 12'b011001001010;
   5835: result <= 12'b011001001001;
   5836: result <= 12'b011001001001;
   5837: result <= 12'b011001001000;
   5838: result <= 12'b011001001000;
   5839: result <= 12'b011001000111;
   5840: result <= 12'b011001000111;
   5841: result <= 12'b011001000110;
   5842: result <= 12'b011001000110;
   5843: result <= 12'b011001000101;
   5844: result <= 12'b011001000101;
   5845: result <= 12'b011001000100;
   5846: result <= 12'b011001000100;
   5847: result <= 12'b011001000011;
   5848: result <= 12'b011001000011;
   5849: result <= 12'b011001000010;
   5850: result <= 12'b011001000010;
   5851: result <= 12'b011001000001;
   5852: result <= 12'b011001000001;
   5853: result <= 12'b011001000000;
   5854: result <= 12'b011001000000;
   5855: result <= 12'b011000111111;
   5856: result <= 12'b011000111111;
   5857: result <= 12'b011000111110;
   5858: result <= 12'b011000111110;
   5859: result <= 12'b011000111101;
   5860: result <= 12'b011000111101;
   5861: result <= 12'b011000111100;
   5862: result <= 12'b011000111100;
   5863: result <= 12'b011000111100;
   5864: result <= 12'b011000111011;
   5865: result <= 12'b011000111011;
   5866: result <= 12'b011000111010;
   5867: result <= 12'b011000111010;
   5868: result <= 12'b011000111001;
   5869: result <= 12'b011000111001;
   5870: result <= 12'b011000111000;
   5871: result <= 12'b011000111000;
   5872: result <= 12'b011000110111;
   5873: result <= 12'b011000110111;
   5874: result <= 12'b011000110110;
   5875: result <= 12'b011000110110;
   5876: result <= 12'b011000110101;
   5877: result <= 12'b011000110101;
   5878: result <= 12'b011000110100;
   5879: result <= 12'b011000110100;
   5880: result <= 12'b011000110011;
   5881: result <= 12'b011000110011;
   5882: result <= 12'b011000110010;
   5883: result <= 12'b011000110010;
   5884: result <= 12'b011000110001;
   5885: result <= 12'b011000110001;
   5886: result <= 12'b011000110000;
   5887: result <= 12'b011000110000;
   5888: result <= 12'b011000101111;
   5889: result <= 12'b011000101111;
   5890: result <= 12'b011000101110;
   5891: result <= 12'b011000101110;
   5892: result <= 12'b011000101101;
   5893: result <= 12'b011000101101;
   5894: result <= 12'b011000101100;
   5895: result <= 12'b011000101100;
   5896: result <= 12'b011000101011;
   5897: result <= 12'b011000101011;
   5898: result <= 12'b011000101010;
   5899: result <= 12'b011000101010;
   5900: result <= 12'b011000101001;
   5901: result <= 12'b011000101001;
   5902: result <= 12'b011000101000;
   5903: result <= 12'b011000101000;
   5904: result <= 12'b011000100111;
   5905: result <= 12'b011000100111;
   5906: result <= 12'b011000100110;
   5907: result <= 12'b011000100110;
   5908: result <= 12'b011000100101;
   5909: result <= 12'b011000100101;
   5910: result <= 12'b011000100100;
   5911: result <= 12'b011000100100;
   5912: result <= 12'b011000100011;
   5913: result <= 12'b011000100011;
   5914: result <= 12'b011000100010;
   5915: result <= 12'b011000100010;
   5916: result <= 12'b011000100001;
   5917: result <= 12'b011000100001;
   5918: result <= 12'b011000100000;
   5919: result <= 12'b011000100000;
   5920: result <= 12'b011000011111;
   5921: result <= 12'b011000011111;
   5922: result <= 12'b011000011110;
   5923: result <= 12'b011000011110;
   5924: result <= 12'b011000011101;
   5925: result <= 12'b011000011101;
   5926: result <= 12'b011000011100;
   5927: result <= 12'b011000011100;
   5928: result <= 12'b011000011011;
   5929: result <= 12'b011000011011;
   5930: result <= 12'b011000011010;
   5931: result <= 12'b011000011001;
   5932: result <= 12'b011000011001;
   5933: result <= 12'b011000011000;
   5934: result <= 12'b011000011000;
   5935: result <= 12'b011000010111;
   5936: result <= 12'b011000010111;
   5937: result <= 12'b011000010110;
   5938: result <= 12'b011000010110;
   5939: result <= 12'b011000010101;
   5940: result <= 12'b011000010101;
   5941: result <= 12'b011000010100;
   5942: result <= 12'b011000010100;
   5943: result <= 12'b011000010011;
   5944: result <= 12'b011000010011;
   5945: result <= 12'b011000010010;
   5946: result <= 12'b011000010010;
   5947: result <= 12'b011000010001;
   5948: result <= 12'b011000010001;
   5949: result <= 12'b011000010000;
   5950: result <= 12'b011000010000;
   5951: result <= 12'b011000001111;
   5952: result <= 12'b011000001111;
   5953: result <= 12'b011000001110;
   5954: result <= 12'b011000001110;
   5955: result <= 12'b011000001101;
   5956: result <= 12'b011000001101;
   5957: result <= 12'b011000001100;
   5958: result <= 12'b011000001100;
   5959: result <= 12'b011000001011;
   5960: result <= 12'b011000001011;
   5961: result <= 12'b011000001010;
   5962: result <= 12'b011000001010;
   5963: result <= 12'b011000001001;
   5964: result <= 12'b011000001001;
   5965: result <= 12'b011000001000;
   5966: result <= 12'b011000001000;
   5967: result <= 12'b011000000111;
   5968: result <= 12'b011000000111;
   5969: result <= 12'b011000000110;
   5970: result <= 12'b011000000101;
   5971: result <= 12'b011000000101;
   5972: result <= 12'b011000000100;
   5973: result <= 12'b011000000100;
   5974: result <= 12'b011000000011;
   5975: result <= 12'b011000000011;
   5976: result <= 12'b011000000010;
   5977: result <= 12'b011000000010;
   5978: result <= 12'b011000000001;
   5979: result <= 12'b011000000001;
   5980: result <= 12'b011000000000;
   5981: result <= 12'b011000000000;
   5982: result <= 12'b010111111111;
   5983: result <= 12'b010111111111;
   5984: result <= 12'b010111111110;
   5985: result <= 12'b010111111110;
   5986: result <= 12'b010111111101;
   5987: result <= 12'b010111111101;
   5988: result <= 12'b010111111100;
   5989: result <= 12'b010111111100;
   5990: result <= 12'b010111111011;
   5991: result <= 12'b010111111011;
   5992: result <= 12'b010111111010;
   5993: result <= 12'b010111111010;
   5994: result <= 12'b010111111001;
   5995: result <= 12'b010111111000;
   5996: result <= 12'b010111111000;
   5997: result <= 12'b010111110111;
   5998: result <= 12'b010111110111;
   5999: result <= 12'b010111110110;
   6000: result <= 12'b010111110110;
   6001: result <= 12'b010111110101;
   6002: result <= 12'b010111110101;
   6003: result <= 12'b010111110100;
   6004: result <= 12'b010111110100;
   6005: result <= 12'b010111110011;
   6006: result <= 12'b010111110011;
   6007: result <= 12'b010111110010;
   6008: result <= 12'b010111110010;
   6009: result <= 12'b010111110001;
   6010: result <= 12'b010111110001;
   6011: result <= 12'b010111110000;
   6012: result <= 12'b010111110000;
   6013: result <= 12'b010111101111;
   6014: result <= 12'b010111101111;
   6015: result <= 12'b010111101110;
   6016: result <= 12'b010111101101;
   6017: result <= 12'b010111101101;
   6018: result <= 12'b010111101100;
   6019: result <= 12'b010111101100;
   6020: result <= 12'b010111101011;
   6021: result <= 12'b010111101011;
   6022: result <= 12'b010111101010;
   6023: result <= 12'b010111101010;
   6024: result <= 12'b010111101001;
   6025: result <= 12'b010111101001;
   6026: result <= 12'b010111101000;
   6027: result <= 12'b010111101000;
   6028: result <= 12'b010111100111;
   6029: result <= 12'b010111100111;
   6030: result <= 12'b010111100110;
   6031: result <= 12'b010111100110;
   6032: result <= 12'b010111100101;
   6033: result <= 12'b010111100100;
   6034: result <= 12'b010111100100;
   6035: result <= 12'b010111100011;
   6036: result <= 12'b010111100011;
   6037: result <= 12'b010111100010;
   6038: result <= 12'b010111100010;
   6039: result <= 12'b010111100001;
   6040: result <= 12'b010111100001;
   6041: result <= 12'b010111100000;
   6042: result <= 12'b010111100000;
   6043: result <= 12'b010111011111;
   6044: result <= 12'b010111011111;
   6045: result <= 12'b010111011110;
   6046: result <= 12'b010111011110;
   6047: result <= 12'b010111011101;
   6048: result <= 12'b010111011100;
   6049: result <= 12'b010111011100;
   6050: result <= 12'b010111011011;
   6051: result <= 12'b010111011011;
   6052: result <= 12'b010111011010;
   6053: result <= 12'b010111011010;
   6054: result <= 12'b010111011001;
   6055: result <= 12'b010111011001;
   6056: result <= 12'b010111011000;
   6057: result <= 12'b010111011000;
   6058: result <= 12'b010111010111;
   6059: result <= 12'b010111010111;
   6060: result <= 12'b010111010110;
   6061: result <= 12'b010111010110;
   6062: result <= 12'b010111010101;
   6063: result <= 12'b010111010100;
   6064: result <= 12'b010111010100;
   6065: result <= 12'b010111010011;
   6066: result <= 12'b010111010011;
   6067: result <= 12'b010111010010;
   6068: result <= 12'b010111010010;
   6069: result <= 12'b010111010001;
   6070: result <= 12'b010111010001;
   6071: result <= 12'b010111010000;
   6072: result <= 12'b010111010000;
   6073: result <= 12'b010111001111;
   6074: result <= 12'b010111001111;
   6075: result <= 12'b010111001110;
   6076: result <= 12'b010111001101;
   6077: result <= 12'b010111001101;
   6078: result <= 12'b010111001100;
   6079: result <= 12'b010111001100;
   6080: result <= 12'b010111001011;
   6081: result <= 12'b010111001011;
   6082: result <= 12'b010111001010;
   6083: result <= 12'b010111001010;
   6084: result <= 12'b010111001001;
   6085: result <= 12'b010111001001;
   6086: result <= 12'b010111001000;
   6087: result <= 12'b010111000111;
   6088: result <= 12'b010111000111;
   6089: result <= 12'b010111000110;
   6090: result <= 12'b010111000110;
   6091: result <= 12'b010111000101;
   6092: result <= 12'b010111000101;
   6093: result <= 12'b010111000100;
   6094: result <= 12'b010111000100;
   6095: result <= 12'b010111000011;
   6096: result <= 12'b010111000011;
   6097: result <= 12'b010111000010;
   6098: result <= 12'b010111000001;
   6099: result <= 12'b010111000001;
   6100: result <= 12'b010111000000;
   6101: result <= 12'b010111000000;
   6102: result <= 12'b010110111111;
   6103: result <= 12'b010110111111;
   6104: result <= 12'b010110111110;
   6105: result <= 12'b010110111110;
   6106: result <= 12'b010110111101;
   6107: result <= 12'b010110111101;
   6108: result <= 12'b010110111100;
   6109: result <= 12'b010110111011;
   6110: result <= 12'b010110111011;
   6111: result <= 12'b010110111010;
   6112: result <= 12'b010110111010;
   6113: result <= 12'b010110111001;
   6114: result <= 12'b010110111001;
   6115: result <= 12'b010110111000;
   6116: result <= 12'b010110111000;
   6117: result <= 12'b010110110111;
   6118: result <= 12'b010110110111;
   6119: result <= 12'b010110110110;
   6120: result <= 12'b010110110101;
   6121: result <= 12'b010110110101;
   6122: result <= 12'b010110110100;
   6123: result <= 12'b010110110100;
   6124: result <= 12'b010110110011;
   6125: result <= 12'b010110110011;
   6126: result <= 12'b010110110010;
   6127: result <= 12'b010110110010;
   6128: result <= 12'b010110110001;
   6129: result <= 12'b010110110000;
   6130: result <= 12'b010110110000;
   6131: result <= 12'b010110101111;
   6132: result <= 12'b010110101111;
   6133: result <= 12'b010110101110;
   6134: result <= 12'b010110101110;
   6135: result <= 12'b010110101101;
   6136: result <= 12'b010110101101;
   6137: result <= 12'b010110101100;
   6138: result <= 12'b010110101011;
   6139: result <= 12'b010110101011;
   6140: result <= 12'b010110101010;
   6141: result <= 12'b010110101010;
   6142: result <= 12'b010110101001;
   6143: result <= 12'b010110101001;
   6144: result <= 12'b010110101000;
   6145: result <= 12'b010110101000;
   6146: result <= 12'b010110100111;
   6147: result <= 12'b010110100110;
   6148: result <= 12'b010110100110;
   6149: result <= 12'b010110100101;
   6150: result <= 12'b010110100101;
   6151: result <= 12'b010110100100;
   6152: result <= 12'b010110100100;
   6153: result <= 12'b010110100011;
   6154: result <= 12'b010110100011;
   6155: result <= 12'b010110100010;
   6156: result <= 12'b010110100001;
   6157: result <= 12'b010110100001;
   6158: result <= 12'b010110100000;
   6159: result <= 12'b010110100000;
   6160: result <= 12'b010110011111;
   6161: result <= 12'b010110011111;
   6162: result <= 12'b010110011110;
   6163: result <= 12'b010110011110;
   6164: result <= 12'b010110011101;
   6165: result <= 12'b010110011100;
   6166: result <= 12'b010110011100;
   6167: result <= 12'b010110011011;
   6168: result <= 12'b010110011011;
   6169: result <= 12'b010110011010;
   6170: result <= 12'b010110011010;
   6171: result <= 12'b010110011001;
   6172: result <= 12'b010110011001;
   6173: result <= 12'b010110011000;
   6174: result <= 12'b010110010111;
   6175: result <= 12'b010110010111;
   6176: result <= 12'b010110010110;
   6177: result <= 12'b010110010110;
   6178: result <= 12'b010110010101;
   6179: result <= 12'b010110010101;
   6180: result <= 12'b010110010100;
   6181: result <= 12'b010110010011;
   6182: result <= 12'b010110010011;
   6183: result <= 12'b010110010010;
   6184: result <= 12'b010110010010;
   6185: result <= 12'b010110010001;
   6186: result <= 12'b010110010001;
   6187: result <= 12'b010110010000;
   6188: result <= 12'b010110010000;
   6189: result <= 12'b010110001111;
   6190: result <= 12'b010110001110;
   6191: result <= 12'b010110001110;
   6192: result <= 12'b010110001101;
   6193: result <= 12'b010110001101;
   6194: result <= 12'b010110001100;
   6195: result <= 12'b010110001100;
   6196: result <= 12'b010110001011;
   6197: result <= 12'b010110001010;
   6198: result <= 12'b010110001010;
   6199: result <= 12'b010110001001;
   6200: result <= 12'b010110001001;
   6201: result <= 12'b010110001000;
   6202: result <= 12'b010110001000;
   6203: result <= 12'b010110000111;
   6204: result <= 12'b010110000110;
   6205: result <= 12'b010110000110;
   6206: result <= 12'b010110000101;
   6207: result <= 12'b010110000101;
   6208: result <= 12'b010110000100;
   6209: result <= 12'b010110000100;
   6210: result <= 12'b010110000011;
   6211: result <= 12'b010110000010;
   6212: result <= 12'b010110000010;
   6213: result <= 12'b010110000001;
   6214: result <= 12'b010110000001;
   6215: result <= 12'b010110000000;
   6216: result <= 12'b010110000000;
   6217: result <= 12'b010101111111;
   6218: result <= 12'b010101111110;
   6219: result <= 12'b010101111110;
   6220: result <= 12'b010101111101;
   6221: result <= 12'b010101111101;
   6222: result <= 12'b010101111100;
   6223: result <= 12'b010101111100;
   6224: result <= 12'b010101111011;
   6225: result <= 12'b010101111010;
   6226: result <= 12'b010101111010;
   6227: result <= 12'b010101111001;
   6228: result <= 12'b010101111001;
   6229: result <= 12'b010101111000;
   6230: result <= 12'b010101111000;
   6231: result <= 12'b010101110111;
   6232: result <= 12'b010101110110;
   6233: result <= 12'b010101110110;
   6234: result <= 12'b010101110101;
   6235: result <= 12'b010101110101;
   6236: result <= 12'b010101110100;
   6237: result <= 12'b010101110100;
   6238: result <= 12'b010101110011;
   6239: result <= 12'b010101110010;
   6240: result <= 12'b010101110010;
   6241: result <= 12'b010101110001;
   6242: result <= 12'b010101110001;
   6243: result <= 12'b010101110000;
   6244: result <= 12'b010101110000;
   6245: result <= 12'b010101101111;
   6246: result <= 12'b010101101110;
   6247: result <= 12'b010101101110;
   6248: result <= 12'b010101101101;
   6249: result <= 12'b010101101101;
   6250: result <= 12'b010101101100;
   6251: result <= 12'b010101101100;
   6252: result <= 12'b010101101011;
   6253: result <= 12'b010101101010;
   6254: result <= 12'b010101101010;
   6255: result <= 12'b010101101001;
   6256: result <= 12'b010101101001;
   6257: result <= 12'b010101101000;
   6258: result <= 12'b010101100111;
   6259: result <= 12'b010101100111;
   6260: result <= 12'b010101100110;
   6261: result <= 12'b010101100110;
   6262: result <= 12'b010101100101;
   6263: result <= 12'b010101100101;
   6264: result <= 12'b010101100100;
   6265: result <= 12'b010101100011;
   6266: result <= 12'b010101100011;
   6267: result <= 12'b010101100010;
   6268: result <= 12'b010101100010;
   6269: result <= 12'b010101100001;
   6270: result <= 12'b010101100001;
   6271: result <= 12'b010101100000;
   6272: result <= 12'b010101011111;
   6273: result <= 12'b010101011111;
   6274: result <= 12'b010101011110;
   6275: result <= 12'b010101011110;
   6276: result <= 12'b010101011101;
   6277: result <= 12'b010101011100;
   6278: result <= 12'b010101011100;
   6279: result <= 12'b010101011011;
   6280: result <= 12'b010101011011;
   6281: result <= 12'b010101011010;
   6282: result <= 12'b010101011010;
   6283: result <= 12'b010101011001;
   6284: result <= 12'b010101011000;
   6285: result <= 12'b010101011000;
   6286: result <= 12'b010101010111;
   6287: result <= 12'b010101010111;
   6288: result <= 12'b010101010110;
   6289: result <= 12'b010101010101;
   6290: result <= 12'b010101010101;
   6291: result <= 12'b010101010100;
   6292: result <= 12'b010101010100;
   6293: result <= 12'b010101010011;
   6294: result <= 12'b010101010011;
   6295: result <= 12'b010101010010;
   6296: result <= 12'b010101010001;
   6297: result <= 12'b010101010001;
   6298: result <= 12'b010101010000;
   6299: result <= 12'b010101010000;
   6300: result <= 12'b010101001111;
   6301: result <= 12'b010101001110;
   6302: result <= 12'b010101001110;
   6303: result <= 12'b010101001101;
   6304: result <= 12'b010101001101;
   6305: result <= 12'b010101001100;
   6306: result <= 12'b010101001011;
   6307: result <= 12'b010101001011;
   6308: result <= 12'b010101001010;
   6309: result <= 12'b010101001010;
   6310: result <= 12'b010101001001;
   6311: result <= 12'b010101001001;
   6312: result <= 12'b010101001000;
   6313: result <= 12'b010101000111;
   6314: result <= 12'b010101000111;
   6315: result <= 12'b010101000110;
   6316: result <= 12'b010101000110;
   6317: result <= 12'b010101000101;
   6318: result <= 12'b010101000100;
   6319: result <= 12'b010101000100;
   6320: result <= 12'b010101000011;
   6321: result <= 12'b010101000011;
   6322: result <= 12'b010101000010;
   6323: result <= 12'b010101000001;
   6324: result <= 12'b010101000001;
   6325: result <= 12'b010101000000;
   6326: result <= 12'b010101000000;
   6327: result <= 12'b010100111111;
   6328: result <= 12'b010100111110;
   6329: result <= 12'b010100111110;
   6330: result <= 12'b010100111101;
   6331: result <= 12'b010100111101;
   6332: result <= 12'b010100111100;
   6333: result <= 12'b010100111011;
   6334: result <= 12'b010100111011;
   6335: result <= 12'b010100111010;
   6336: result <= 12'b010100111010;
   6337: result <= 12'b010100111001;
   6338: result <= 12'b010100111001;
   6339: result <= 12'b010100111000;
   6340: result <= 12'b010100110111;
   6341: result <= 12'b010100110111;
   6342: result <= 12'b010100110110;
   6343: result <= 12'b010100110110;
   6344: result <= 12'b010100110101;
   6345: result <= 12'b010100110100;
   6346: result <= 12'b010100110100;
   6347: result <= 12'b010100110011;
   6348: result <= 12'b010100110011;
   6349: result <= 12'b010100110010;
   6350: result <= 12'b010100110001;
   6351: result <= 12'b010100110001;
   6352: result <= 12'b010100110000;
   6353: result <= 12'b010100110000;
   6354: result <= 12'b010100101111;
   6355: result <= 12'b010100101110;
   6356: result <= 12'b010100101110;
   6357: result <= 12'b010100101101;
   6358: result <= 12'b010100101101;
   6359: result <= 12'b010100101100;
   6360: result <= 12'b010100101011;
   6361: result <= 12'b010100101011;
   6362: result <= 12'b010100101010;
   6363: result <= 12'b010100101010;
   6364: result <= 12'b010100101001;
   6365: result <= 12'b010100101000;
   6366: result <= 12'b010100101000;
   6367: result <= 12'b010100100111;
   6368: result <= 12'b010100100111;
   6369: result <= 12'b010100100110;
   6370: result <= 12'b010100100101;
   6371: result <= 12'b010100100101;
   6372: result <= 12'b010100100100;
   6373: result <= 12'b010100100100;
   6374: result <= 12'b010100100011;
   6375: result <= 12'b010100100010;
   6376: result <= 12'b010100100010;
   6377: result <= 12'b010100100001;
   6378: result <= 12'b010100100001;
   6379: result <= 12'b010100100000;
   6380: result <= 12'b010100011111;
   6381: result <= 12'b010100011111;
   6382: result <= 12'b010100011110;
   6383: result <= 12'b010100011110;
   6384: result <= 12'b010100011101;
   6385: result <= 12'b010100011100;
   6386: result <= 12'b010100011100;
   6387: result <= 12'b010100011011;
   6388: result <= 12'b010100011011;
   6389: result <= 12'b010100011010;
   6390: result <= 12'b010100011001;
   6391: result <= 12'b010100011001;
   6392: result <= 12'b010100011000;
   6393: result <= 12'b010100010111;
   6394: result <= 12'b010100010111;
   6395: result <= 12'b010100010110;
   6396: result <= 12'b010100010110;
   6397: result <= 12'b010100010101;
   6398: result <= 12'b010100010100;
   6399: result <= 12'b010100010100;
   6400: result <= 12'b010100010011;
   6401: result <= 12'b010100010011;
   6402: result <= 12'b010100010010;
   6403: result <= 12'b010100010001;
   6404: result <= 12'b010100010001;
   6405: result <= 12'b010100010000;
   6406: result <= 12'b010100010000;
   6407: result <= 12'b010100001111;
   6408: result <= 12'b010100001110;
   6409: result <= 12'b010100001110;
   6410: result <= 12'b010100001101;
   6411: result <= 12'b010100001101;
   6412: result <= 12'b010100001100;
   6413: result <= 12'b010100001011;
   6414: result <= 12'b010100001011;
   6415: result <= 12'b010100001010;
   6416: result <= 12'b010100001001;
   6417: result <= 12'b010100001001;
   6418: result <= 12'b010100001000;
   6419: result <= 12'b010100001000;
   6420: result <= 12'b010100000111;
   6421: result <= 12'b010100000110;
   6422: result <= 12'b010100000110;
   6423: result <= 12'b010100000101;
   6424: result <= 12'b010100000101;
   6425: result <= 12'b010100000100;
   6426: result <= 12'b010100000011;
   6427: result <= 12'b010100000011;
   6428: result <= 12'b010100000010;
   6429: result <= 12'b010100000010;
   6430: result <= 12'b010100000001;
   6431: result <= 12'b010100000000;
   6432: result <= 12'b010100000000;
   6433: result <= 12'b010011111111;
   6434: result <= 12'b010011111110;
   6435: result <= 12'b010011111110;
   6436: result <= 12'b010011111101;
   6437: result <= 12'b010011111101;
   6438: result <= 12'b010011111100;
   6439: result <= 12'b010011111011;
   6440: result <= 12'b010011111011;
   6441: result <= 12'b010011111010;
   6442: result <= 12'b010011111010;
   6443: result <= 12'b010011111001;
   6444: result <= 12'b010011111000;
   6445: result <= 12'b010011111000;
   6446: result <= 12'b010011110111;
   6447: result <= 12'b010011110110;
   6448: result <= 12'b010011110110;
   6449: result <= 12'b010011110101;
   6450: result <= 12'b010011110101;
   6451: result <= 12'b010011110100;
   6452: result <= 12'b010011110011;
   6453: result <= 12'b010011110011;
   6454: result <= 12'b010011110010;
   6455: result <= 12'b010011110010;
   6456: result <= 12'b010011110001;
   6457: result <= 12'b010011110000;
   6458: result <= 12'b010011110000;
   6459: result <= 12'b010011101111;
   6460: result <= 12'b010011101110;
   6461: result <= 12'b010011101110;
   6462: result <= 12'b010011101101;
   6463: result <= 12'b010011101101;
   6464: result <= 12'b010011101100;
   6465: result <= 12'b010011101011;
   6466: result <= 12'b010011101011;
   6467: result <= 12'b010011101010;
   6468: result <= 12'b010011101010;
   6469: result <= 12'b010011101001;
   6470: result <= 12'b010011101000;
   6471: result <= 12'b010011101000;
   6472: result <= 12'b010011100111;
   6473: result <= 12'b010011100110;
   6474: result <= 12'b010011100110;
   6475: result <= 12'b010011100101;
   6476: result <= 12'b010011100101;
   6477: result <= 12'b010011100100;
   6478: result <= 12'b010011100011;
   6479: result <= 12'b010011100011;
   6480: result <= 12'b010011100010;
   6481: result <= 12'b010011100001;
   6482: result <= 12'b010011100001;
   6483: result <= 12'b010011100000;
   6484: result <= 12'b010011100000;
   6485: result <= 12'b010011011111;
   6486: result <= 12'b010011011110;
   6487: result <= 12'b010011011110;
   6488: result <= 12'b010011011101;
   6489: result <= 12'b010011011100;
   6490: result <= 12'b010011011100;
   6491: result <= 12'b010011011011;
   6492: result <= 12'b010011011011;
   6493: result <= 12'b010011011010;
   6494: result <= 12'b010011011001;
   6495: result <= 12'b010011011001;
   6496: result <= 12'b010011011000;
   6497: result <= 12'b010011010111;
   6498: result <= 12'b010011010111;
   6499: result <= 12'b010011010110;
   6500: result <= 12'b010011010110;
   6501: result <= 12'b010011010101;
   6502: result <= 12'b010011010100;
   6503: result <= 12'b010011010100;
   6504: result <= 12'b010011010011;
   6505: result <= 12'b010011010010;
   6506: result <= 12'b010011010010;
   6507: result <= 12'b010011010001;
   6508: result <= 12'b010011010001;
   6509: result <= 12'b010011010000;
   6510: result <= 12'b010011001111;
   6511: result <= 12'b010011001111;
   6512: result <= 12'b010011001110;
   6513: result <= 12'b010011001101;
   6514: result <= 12'b010011001101;
   6515: result <= 12'b010011001100;
   6516: result <= 12'b010011001100;
   6517: result <= 12'b010011001011;
   6518: result <= 12'b010011001010;
   6519: result <= 12'b010011001010;
   6520: result <= 12'b010011001001;
   6521: result <= 12'b010011001000;
   6522: result <= 12'b010011001000;
   6523: result <= 12'b010011000111;
   6524: result <= 12'b010011000111;
   6525: result <= 12'b010011000110;
   6526: result <= 12'b010011000101;
   6527: result <= 12'b010011000101;
   6528: result <= 12'b010011000100;
   6529: result <= 12'b010011000011;
   6530: result <= 12'b010011000011;
   6531: result <= 12'b010011000010;
   6532: result <= 12'b010011000001;
   6533: result <= 12'b010011000001;
   6534: result <= 12'b010011000000;
   6535: result <= 12'b010011000000;
   6536: result <= 12'b010010111111;
   6537: result <= 12'b010010111110;
   6538: result <= 12'b010010111110;
   6539: result <= 12'b010010111101;
   6540: result <= 12'b010010111100;
   6541: result <= 12'b010010111100;
   6542: result <= 12'b010010111011;
   6543: result <= 12'b010010111011;
   6544: result <= 12'b010010111010;
   6545: result <= 12'b010010111001;
   6546: result <= 12'b010010111001;
   6547: result <= 12'b010010111000;
   6548: result <= 12'b010010110111;
   6549: result <= 12'b010010110111;
   6550: result <= 12'b010010110110;
   6551: result <= 12'b010010110101;
   6552: result <= 12'b010010110101;
   6553: result <= 12'b010010110100;
   6554: result <= 12'b010010110100;
   6555: result <= 12'b010010110011;
   6556: result <= 12'b010010110010;
   6557: result <= 12'b010010110010;
   6558: result <= 12'b010010110001;
   6559: result <= 12'b010010110000;
   6560: result <= 12'b010010110000;
   6561: result <= 12'b010010101111;
   6562: result <= 12'b010010101110;
   6563: result <= 12'b010010101110;
   6564: result <= 12'b010010101101;
   6565: result <= 12'b010010101101;
   6566: result <= 12'b010010101100;
   6567: result <= 12'b010010101011;
   6568: result <= 12'b010010101011;
   6569: result <= 12'b010010101010;
   6570: result <= 12'b010010101001;
   6571: result <= 12'b010010101001;
   6572: result <= 12'b010010101000;
   6573: result <= 12'b010010100111;
   6574: result <= 12'b010010100111;
   6575: result <= 12'b010010100110;
   6576: result <= 12'b010010100110;
   6577: result <= 12'b010010100101;
   6578: result <= 12'b010010100100;
   6579: result <= 12'b010010100100;
   6580: result <= 12'b010010100011;
   6581: result <= 12'b010010100010;
   6582: result <= 12'b010010100010;
   6583: result <= 12'b010010100001;
   6584: result <= 12'b010010100000;
   6585: result <= 12'b010010100000;
   6586: result <= 12'b010010011111;
   6587: result <= 12'b010010011110;
   6588: result <= 12'b010010011110;
   6589: result <= 12'b010010011101;
   6590: result <= 12'b010010011101;
   6591: result <= 12'b010010011100;
   6592: result <= 12'b010010011011;
   6593: result <= 12'b010010011011;
   6594: result <= 12'b010010011010;
   6595: result <= 12'b010010011001;
   6596: result <= 12'b010010011001;
   6597: result <= 12'b010010011000;
   6598: result <= 12'b010010010111;
   6599: result <= 12'b010010010111;
   6600: result <= 12'b010010010110;
   6601: result <= 12'b010010010101;
   6602: result <= 12'b010010010101;
   6603: result <= 12'b010010010100;
   6604: result <= 12'b010010010100;
   6605: result <= 12'b010010010011;
   6606: result <= 12'b010010010010;
   6607: result <= 12'b010010010010;
   6608: result <= 12'b010010010001;
   6609: result <= 12'b010010010000;
   6610: result <= 12'b010010010000;
   6611: result <= 12'b010010001111;
   6612: result <= 12'b010010001110;
   6613: result <= 12'b010010001110;
   6614: result <= 12'b010010001101;
   6615: result <= 12'b010010001100;
   6616: result <= 12'b010010001100;
   6617: result <= 12'b010010001011;
   6618: result <= 12'b010010001011;
   6619: result <= 12'b010010001010;
   6620: result <= 12'b010010001001;
   6621: result <= 12'b010010001001;
   6622: result <= 12'b010010001000;
   6623: result <= 12'b010010000111;
   6624: result <= 12'b010010000111;
   6625: result <= 12'b010010000110;
   6626: result <= 12'b010010000101;
   6627: result <= 12'b010010000101;
   6628: result <= 12'b010010000100;
   6629: result <= 12'b010010000011;
   6630: result <= 12'b010010000011;
   6631: result <= 12'b010010000010;
   6632: result <= 12'b010010000001;
   6633: result <= 12'b010010000001;
   6634: result <= 12'b010010000000;
   6635: result <= 12'b010001111111;
   6636: result <= 12'b010001111111;
   6637: result <= 12'b010001111110;
   6638: result <= 12'b010001111110;
   6639: result <= 12'b010001111101;
   6640: result <= 12'b010001111100;
   6641: result <= 12'b010001111100;
   6642: result <= 12'b010001111011;
   6643: result <= 12'b010001111010;
   6644: result <= 12'b010001111010;
   6645: result <= 12'b010001111001;
   6646: result <= 12'b010001111000;
   6647: result <= 12'b010001111000;
   6648: result <= 12'b010001110111;
   6649: result <= 12'b010001110110;
   6650: result <= 12'b010001110110;
   6651: result <= 12'b010001110101;
   6652: result <= 12'b010001110100;
   6653: result <= 12'b010001110100;
   6654: result <= 12'b010001110011;
   6655: result <= 12'b010001110010;
   6656: result <= 12'b010001110010;
   6657: result <= 12'b010001110001;
   6658: result <= 12'b010001110001;
   6659: result <= 12'b010001110000;
   6660: result <= 12'b010001101111;
   6661: result <= 12'b010001101111;
   6662: result <= 12'b010001101110;
   6663: result <= 12'b010001101101;
   6664: result <= 12'b010001101101;
   6665: result <= 12'b010001101100;
   6666: result <= 12'b010001101011;
   6667: result <= 12'b010001101011;
   6668: result <= 12'b010001101010;
   6669: result <= 12'b010001101001;
   6670: result <= 12'b010001101001;
   6671: result <= 12'b010001101000;
   6672: result <= 12'b010001100111;
   6673: result <= 12'b010001100111;
   6674: result <= 12'b010001100110;
   6675: result <= 12'b010001100101;
   6676: result <= 12'b010001100101;
   6677: result <= 12'b010001100100;
   6678: result <= 12'b010001100011;
   6679: result <= 12'b010001100011;
   6680: result <= 12'b010001100010;
   6681: result <= 12'b010001100001;
   6682: result <= 12'b010001100001;
   6683: result <= 12'b010001100000;
   6684: result <= 12'b010001011111;
   6685: result <= 12'b010001011111;
   6686: result <= 12'b010001011110;
   6687: result <= 12'b010001011101;
   6688: result <= 12'b010001011101;
   6689: result <= 12'b010001011100;
   6690: result <= 12'b010001011100;
   6691: result <= 12'b010001011011;
   6692: result <= 12'b010001011010;
   6693: result <= 12'b010001011010;
   6694: result <= 12'b010001011001;
   6695: result <= 12'b010001011000;
   6696: result <= 12'b010001011000;
   6697: result <= 12'b010001010111;
   6698: result <= 12'b010001010110;
   6699: result <= 12'b010001010110;
   6700: result <= 12'b010001010101;
   6701: result <= 12'b010001010100;
   6702: result <= 12'b010001010100;
   6703: result <= 12'b010001010011;
   6704: result <= 12'b010001010010;
   6705: result <= 12'b010001010010;
   6706: result <= 12'b010001010001;
   6707: result <= 12'b010001010000;
   6708: result <= 12'b010001010000;
   6709: result <= 12'b010001001111;
   6710: result <= 12'b010001001110;
   6711: result <= 12'b010001001110;
   6712: result <= 12'b010001001101;
   6713: result <= 12'b010001001100;
   6714: result <= 12'b010001001100;
   6715: result <= 12'b010001001011;
   6716: result <= 12'b010001001010;
   6717: result <= 12'b010001001010;
   6718: result <= 12'b010001001001;
   6719: result <= 12'b010001001000;
   6720: result <= 12'b010001001000;
   6721: result <= 12'b010001000111;
   6722: result <= 12'b010001000110;
   6723: result <= 12'b010001000110;
   6724: result <= 12'b010001000101;
   6725: result <= 12'b010001000100;
   6726: result <= 12'b010001000100;
   6727: result <= 12'b010001000011;
   6728: result <= 12'b010001000010;
   6729: result <= 12'b010001000010;
   6730: result <= 12'b010001000001;
   6731: result <= 12'b010001000000;
   6732: result <= 12'b010001000000;
   6733: result <= 12'b010000111111;
   6734: result <= 12'b010000111110;
   6735: result <= 12'b010000111110;
   6736: result <= 12'b010000111101;
   6737: result <= 12'b010000111100;
   6738: result <= 12'b010000111100;
   6739: result <= 12'b010000111011;
   6740: result <= 12'b010000111010;
   6741: result <= 12'b010000111010;
   6742: result <= 12'b010000111001;
   6743: result <= 12'b010000111000;
   6744: result <= 12'b010000111000;
   6745: result <= 12'b010000110111;
   6746: result <= 12'b010000110110;
   6747: result <= 12'b010000110110;
   6748: result <= 12'b010000110101;
   6749: result <= 12'b010000110100;
   6750: result <= 12'b010000110100;
   6751: result <= 12'b010000110011;
   6752: result <= 12'b010000110010;
   6753: result <= 12'b010000110010;
   6754: result <= 12'b010000110001;
   6755: result <= 12'b010000110000;
   6756: result <= 12'b010000110000;
   6757: result <= 12'b010000101111;
   6758: result <= 12'b010000101110;
   6759: result <= 12'b010000101110;
   6760: result <= 12'b010000101101;
   6761: result <= 12'b010000101100;
   6762: result <= 12'b010000101100;
   6763: result <= 12'b010000101011;
   6764: result <= 12'b010000101010;
   6765: result <= 12'b010000101010;
   6766: result <= 12'b010000101001;
   6767: result <= 12'b010000101000;
   6768: result <= 12'b010000101000;
   6769: result <= 12'b010000100111;
   6770: result <= 12'b010000100110;
   6771: result <= 12'b010000100110;
   6772: result <= 12'b010000100101;
   6773: result <= 12'b010000100100;
   6774: result <= 12'b010000100100;
   6775: result <= 12'b010000100011;
   6776: result <= 12'b010000100010;
   6777: result <= 12'b010000100010;
   6778: result <= 12'b010000100001;
   6779: result <= 12'b010000100000;
   6780: result <= 12'b010000100000;
   6781: result <= 12'b010000011111;
   6782: result <= 12'b010000011110;
   6783: result <= 12'b010000011110;
   6784: result <= 12'b010000011101;
   6785: result <= 12'b010000011100;
   6786: result <= 12'b010000011100;
   6787: result <= 12'b010000011011;
   6788: result <= 12'b010000011010;
   6789: result <= 12'b010000011010;
   6790: result <= 12'b010000011001;
   6791: result <= 12'b010000011000;
   6792: result <= 12'b010000010111;
   6793: result <= 12'b010000010111;
   6794: result <= 12'b010000010110;
   6795: result <= 12'b010000010101;
   6796: result <= 12'b010000010101;
   6797: result <= 12'b010000010100;
   6798: result <= 12'b010000010011;
   6799: result <= 12'b010000010011;
   6800: result <= 12'b010000010010;
   6801: result <= 12'b010000010001;
   6802: result <= 12'b010000010001;
   6803: result <= 12'b010000010000;
   6804: result <= 12'b010000001111;
   6805: result <= 12'b010000001111;
   6806: result <= 12'b010000001110;
   6807: result <= 12'b010000001101;
   6808: result <= 12'b010000001101;
   6809: result <= 12'b010000001100;
   6810: result <= 12'b010000001011;
   6811: result <= 12'b010000001011;
   6812: result <= 12'b010000001010;
   6813: result <= 12'b010000001001;
   6814: result <= 12'b010000001001;
   6815: result <= 12'b010000001000;
   6816: result <= 12'b010000000111;
   6817: result <= 12'b010000000111;
   6818: result <= 12'b010000000110;
   6819: result <= 12'b010000000101;
   6820: result <= 12'b010000000101;
   6821: result <= 12'b010000000100;
   6822: result <= 12'b010000000011;
   6823: result <= 12'b010000000010;
   6824: result <= 12'b010000000010;
   6825: result <= 12'b010000000001;
   6826: result <= 12'b010000000000;
   6827: result <= 12'b010000000000;
   6828: result <= 12'b001111111111;
   6829: result <= 12'b001111111110;
   6830: result <= 12'b001111111110;
   6831: result <= 12'b001111111101;
   6832: result <= 12'b001111111100;
   6833: result <= 12'b001111111100;
   6834: result <= 12'b001111111011;
   6835: result <= 12'b001111111010;
   6836: result <= 12'b001111111010;
   6837: result <= 12'b001111111001;
   6838: result <= 12'b001111111000;
   6839: result <= 12'b001111111000;
   6840: result <= 12'b001111110111;
   6841: result <= 12'b001111110110;
   6842: result <= 12'b001111110110;
   6843: result <= 12'b001111110101;
   6844: result <= 12'b001111110100;
   6845: result <= 12'b001111110100;
   6846: result <= 12'b001111110011;
   6847: result <= 12'b001111110010;
   6848: result <= 12'b001111110001;
   6849: result <= 12'b001111110001;
   6850: result <= 12'b001111110000;
   6851: result <= 12'b001111101111;
   6852: result <= 12'b001111101111;
   6853: result <= 12'b001111101110;
   6854: result <= 12'b001111101101;
   6855: result <= 12'b001111101101;
   6856: result <= 12'b001111101100;
   6857: result <= 12'b001111101011;
   6858: result <= 12'b001111101011;
   6859: result <= 12'b001111101010;
   6860: result <= 12'b001111101001;
   6861: result <= 12'b001111101001;
   6862: result <= 12'b001111101000;
   6863: result <= 12'b001111100111;
   6864: result <= 12'b001111100111;
   6865: result <= 12'b001111100110;
   6866: result <= 12'b001111100101;
   6867: result <= 12'b001111100100;
   6868: result <= 12'b001111100100;
   6869: result <= 12'b001111100011;
   6870: result <= 12'b001111100010;
   6871: result <= 12'b001111100010;
   6872: result <= 12'b001111100001;
   6873: result <= 12'b001111100000;
   6874: result <= 12'b001111100000;
   6875: result <= 12'b001111011111;
   6876: result <= 12'b001111011110;
   6877: result <= 12'b001111011110;
   6878: result <= 12'b001111011101;
   6879: result <= 12'b001111011100;
   6880: result <= 12'b001111011100;
   6881: result <= 12'b001111011011;
   6882: result <= 12'b001111011010;
   6883: result <= 12'b001111011001;
   6884: result <= 12'b001111011001;
   6885: result <= 12'b001111011000;
   6886: result <= 12'b001111010111;
   6887: result <= 12'b001111010111;
   6888: result <= 12'b001111010110;
   6889: result <= 12'b001111010101;
   6890: result <= 12'b001111010101;
   6891: result <= 12'b001111010100;
   6892: result <= 12'b001111010011;
   6893: result <= 12'b001111010011;
   6894: result <= 12'b001111010010;
   6895: result <= 12'b001111010001;
   6896: result <= 12'b001111010000;
   6897: result <= 12'b001111010000;
   6898: result <= 12'b001111001111;
   6899: result <= 12'b001111001110;
   6900: result <= 12'b001111001110;
   6901: result <= 12'b001111001101;
   6902: result <= 12'b001111001100;
   6903: result <= 12'b001111001100;
   6904: result <= 12'b001111001011;
   6905: result <= 12'b001111001010;
   6906: result <= 12'b001111001010;
   6907: result <= 12'b001111001001;
   6908: result <= 12'b001111001000;
   6909: result <= 12'b001111000111;
   6910: result <= 12'b001111000111;
   6911: result <= 12'b001111000110;
   6912: result <= 12'b001111000101;
   6913: result <= 12'b001111000101;
   6914: result <= 12'b001111000100;
   6915: result <= 12'b001111000011;
   6916: result <= 12'b001111000011;
   6917: result <= 12'b001111000010;
   6918: result <= 12'b001111000001;
   6919: result <= 12'b001111000001;
   6920: result <= 12'b001111000000;
   6921: result <= 12'b001110111111;
   6922: result <= 12'b001110111110;
   6923: result <= 12'b001110111110;
   6924: result <= 12'b001110111101;
   6925: result <= 12'b001110111100;
   6926: result <= 12'b001110111100;
   6927: result <= 12'b001110111011;
   6928: result <= 12'b001110111010;
   6929: result <= 12'b001110111010;
   6930: result <= 12'b001110111001;
   6931: result <= 12'b001110111000;
   6932: result <= 12'b001110111000;
   6933: result <= 12'b001110110111;
   6934: result <= 12'b001110110110;
   6935: result <= 12'b001110110101;
   6936: result <= 12'b001110110101;
   6937: result <= 12'b001110110100;
   6938: result <= 12'b001110110011;
   6939: result <= 12'b001110110011;
   6940: result <= 12'b001110110010;
   6941: result <= 12'b001110110001;
   6942: result <= 12'b001110110001;
   6943: result <= 12'b001110110000;
   6944: result <= 12'b001110101111;
   6945: result <= 12'b001110101110;
   6946: result <= 12'b001110101110;
   6947: result <= 12'b001110101101;
   6948: result <= 12'b001110101100;
   6949: result <= 12'b001110101100;
   6950: result <= 12'b001110101011;
   6951: result <= 12'b001110101010;
   6952: result <= 12'b001110101010;
   6953: result <= 12'b001110101001;
   6954: result <= 12'b001110101000;
   6955: result <= 12'b001110101000;
   6956: result <= 12'b001110100111;
   6957: result <= 12'b001110100110;
   6958: result <= 12'b001110100101;
   6959: result <= 12'b001110100101;
   6960: result <= 12'b001110100100;
   6961: result <= 12'b001110100011;
   6962: result <= 12'b001110100011;
   6963: result <= 12'b001110100010;
   6964: result <= 12'b001110100001;
   6965: result <= 12'b001110100001;
   6966: result <= 12'b001110100000;
   6967: result <= 12'b001110011111;
   6968: result <= 12'b001110011110;
   6969: result <= 12'b001110011110;
   6970: result <= 12'b001110011101;
   6971: result <= 12'b001110011100;
   6972: result <= 12'b001110011100;
   6973: result <= 12'b001110011011;
   6974: result <= 12'b001110011010;
   6975: result <= 12'b001110011010;
   6976: result <= 12'b001110011001;
   6977: result <= 12'b001110011000;
   6978: result <= 12'b001110010111;
   6979: result <= 12'b001110010111;
   6980: result <= 12'b001110010110;
   6981: result <= 12'b001110010101;
   6982: result <= 12'b001110010101;
   6983: result <= 12'b001110010100;
   6984: result <= 12'b001110010011;
   6985: result <= 12'b001110010010;
   6986: result <= 12'b001110010010;
   6987: result <= 12'b001110010001;
   6988: result <= 12'b001110010000;
   6989: result <= 12'b001110010000;
   6990: result <= 12'b001110001111;
   6991: result <= 12'b001110001110;
   6992: result <= 12'b001110001110;
   6993: result <= 12'b001110001101;
   6994: result <= 12'b001110001100;
   6995: result <= 12'b001110001011;
   6996: result <= 12'b001110001011;
   6997: result <= 12'b001110001010;
   6998: result <= 12'b001110001001;
   6999: result <= 12'b001110001001;
   7000: result <= 12'b001110001000;
   7001: result <= 12'b001110000111;
   7002: result <= 12'b001110000111;
   7003: result <= 12'b001110000110;
   7004: result <= 12'b001110000101;
   7005: result <= 12'b001110000100;
   7006: result <= 12'b001110000100;
   7007: result <= 12'b001110000011;
   7008: result <= 12'b001110000010;
   7009: result <= 12'b001110000010;
   7010: result <= 12'b001110000001;
   7011: result <= 12'b001110000000;
   7012: result <= 12'b001101111111;
   7013: result <= 12'b001101111111;
   7014: result <= 12'b001101111110;
   7015: result <= 12'b001101111101;
   7016: result <= 12'b001101111101;
   7017: result <= 12'b001101111100;
   7018: result <= 12'b001101111011;
   7019: result <= 12'b001101111011;
   7020: result <= 12'b001101111010;
   7021: result <= 12'b001101111001;
   7022: result <= 12'b001101111000;
   7023: result <= 12'b001101111000;
   7024: result <= 12'b001101110111;
   7025: result <= 12'b001101110110;
   7026: result <= 12'b001101110110;
   7027: result <= 12'b001101110101;
   7028: result <= 12'b001101110100;
   7029: result <= 12'b001101110011;
   7030: result <= 12'b001101110011;
   7031: result <= 12'b001101110010;
   7032: result <= 12'b001101110001;
   7033: result <= 12'b001101110001;
   7034: result <= 12'b001101110000;
   7035: result <= 12'b001101101111;
   7036: result <= 12'b001101101110;
   7037: result <= 12'b001101101110;
   7038: result <= 12'b001101101101;
   7039: result <= 12'b001101101100;
   7040: result <= 12'b001101101100;
   7041: result <= 12'b001101101011;
   7042: result <= 12'b001101101010;
   7043: result <= 12'b001101101010;
   7044: result <= 12'b001101101001;
   7045: result <= 12'b001101101000;
   7046: result <= 12'b001101100111;
   7047: result <= 12'b001101100111;
   7048: result <= 12'b001101100110;
   7049: result <= 12'b001101100101;
   7050: result <= 12'b001101100101;
   7051: result <= 12'b001101100100;
   7052: result <= 12'b001101100011;
   7053: result <= 12'b001101100010;
   7054: result <= 12'b001101100010;
   7055: result <= 12'b001101100001;
   7056: result <= 12'b001101100000;
   7057: result <= 12'b001101100000;
   7058: result <= 12'b001101011111;
   7059: result <= 12'b001101011110;
   7060: result <= 12'b001101011101;
   7061: result <= 12'b001101011101;
   7062: result <= 12'b001101011100;
   7063: result <= 12'b001101011011;
   7064: result <= 12'b001101011011;
   7065: result <= 12'b001101011010;
   7066: result <= 12'b001101011001;
   7067: result <= 12'b001101011000;
   7068: result <= 12'b001101011000;
   7069: result <= 12'b001101010111;
   7070: result <= 12'b001101010110;
   7071: result <= 12'b001101010110;
   7072: result <= 12'b001101010101;
   7073: result <= 12'b001101010100;
   7074: result <= 12'b001101010011;
   7075: result <= 12'b001101010011;
   7076: result <= 12'b001101010010;
   7077: result <= 12'b001101010001;
   7078: result <= 12'b001101010001;
   7079: result <= 12'b001101010000;
   7080: result <= 12'b001101001111;
   7081: result <= 12'b001101001110;
   7082: result <= 12'b001101001110;
   7083: result <= 12'b001101001101;
   7084: result <= 12'b001101001100;
   7085: result <= 12'b001101001100;
   7086: result <= 12'b001101001011;
   7087: result <= 12'b001101001010;
   7088: result <= 12'b001101001001;
   7089: result <= 12'b001101001001;
   7090: result <= 12'b001101001000;
   7091: result <= 12'b001101000111;
   7092: result <= 12'b001101000111;
   7093: result <= 12'b001101000110;
   7094: result <= 12'b001101000101;
   7095: result <= 12'b001101000100;
   7096: result <= 12'b001101000100;
   7097: result <= 12'b001101000011;
   7098: result <= 12'b001101000010;
   7099: result <= 12'b001101000010;
   7100: result <= 12'b001101000001;
   7101: result <= 12'b001101000000;
   7102: result <= 12'b001100111111;
   7103: result <= 12'b001100111111;
   7104: result <= 12'b001100111110;
   7105: result <= 12'b001100111101;
   7106: result <= 12'b001100111100;
   7107: result <= 12'b001100111100;
   7108: result <= 12'b001100111011;
   7109: result <= 12'b001100111010;
   7110: result <= 12'b001100111010;
   7111: result <= 12'b001100111001;
   7112: result <= 12'b001100111000;
   7113: result <= 12'b001100110111;
   7114: result <= 12'b001100110111;
   7115: result <= 12'b001100110110;
   7116: result <= 12'b001100110101;
   7117: result <= 12'b001100110101;
   7118: result <= 12'b001100110100;
   7119: result <= 12'b001100110011;
   7120: result <= 12'b001100110010;
   7121: result <= 12'b001100110010;
   7122: result <= 12'b001100110001;
   7123: result <= 12'b001100110000;
   7124: result <= 12'b001100110000;
   7125: result <= 12'b001100101111;
   7126: result <= 12'b001100101110;
   7127: result <= 12'b001100101101;
   7128: result <= 12'b001100101101;
   7129: result <= 12'b001100101100;
   7130: result <= 12'b001100101011;
   7131: result <= 12'b001100101011;
   7132: result <= 12'b001100101010;
   7133: result <= 12'b001100101001;
   7134: result <= 12'b001100101000;
   7135: result <= 12'b001100101000;
   7136: result <= 12'b001100100111;
   7137: result <= 12'b001100100110;
   7138: result <= 12'b001100100101;
   7139: result <= 12'b001100100101;
   7140: result <= 12'b001100100100;
   7141: result <= 12'b001100100011;
   7142: result <= 12'b001100100011;
   7143: result <= 12'b001100100010;
   7144: result <= 12'b001100100001;
   7145: result <= 12'b001100100000;
   7146: result <= 12'b001100100000;
   7147: result <= 12'b001100011111;
   7148: result <= 12'b001100011110;
   7149: result <= 12'b001100011110;
   7150: result <= 12'b001100011101;
   7151: result <= 12'b001100011100;
   7152: result <= 12'b001100011011;
   7153: result <= 12'b001100011011;
   7154: result <= 12'b001100011010;
   7155: result <= 12'b001100011001;
   7156: result <= 12'b001100011000;
   7157: result <= 12'b001100011000;
   7158: result <= 12'b001100010111;
   7159: result <= 12'b001100010110;
   7160: result <= 12'b001100010110;
   7161: result <= 12'b001100010101;
   7162: result <= 12'b001100010100;
   7163: result <= 12'b001100010011;
   7164: result <= 12'b001100010011;
   7165: result <= 12'b001100010010;
   7166: result <= 12'b001100010001;
   7167: result <= 12'b001100010000;
   7168: result <= 12'b001100010000;
   7169: result <= 12'b001100001111;
   7170: result <= 12'b001100001110;
   7171: result <= 12'b001100001110;
   7172: result <= 12'b001100001101;
   7173: result <= 12'b001100001100;
   7174: result <= 12'b001100001011;
   7175: result <= 12'b001100001011;
   7176: result <= 12'b001100001010;
   7177: result <= 12'b001100001001;
   7178: result <= 12'b001100001000;
   7179: result <= 12'b001100001000;
   7180: result <= 12'b001100000111;
   7181: result <= 12'b001100000110;
   7182: result <= 12'b001100000110;
   7183: result <= 12'b001100000101;
   7184: result <= 12'b001100000100;
   7185: result <= 12'b001100000011;
   7186: result <= 12'b001100000011;
   7187: result <= 12'b001100000010;
   7188: result <= 12'b001100000001;
   7189: result <= 12'b001100000000;
   7190: result <= 12'b001100000000;
   7191: result <= 12'b001011111111;
   7192: result <= 12'b001011111110;
   7193: result <= 12'b001011111110;
   7194: result <= 12'b001011111101;
   7195: result <= 12'b001011111100;
   7196: result <= 12'b001011111011;
   7197: result <= 12'b001011111011;
   7198: result <= 12'b001011111010;
   7199: result <= 12'b001011111001;
   7200: result <= 12'b001011111000;
   7201: result <= 12'b001011111000;
   7202: result <= 12'b001011110111;
   7203: result <= 12'b001011110110;
   7204: result <= 12'b001011110110;
   7205: result <= 12'b001011110101;
   7206: result <= 12'b001011110100;
   7207: result <= 12'b001011110011;
   7208: result <= 12'b001011110011;
   7209: result <= 12'b001011110010;
   7210: result <= 12'b001011110001;
   7211: result <= 12'b001011110000;
   7212: result <= 12'b001011110000;
   7213: result <= 12'b001011101111;
   7214: result <= 12'b001011101110;
   7215: result <= 12'b001011101110;
   7216: result <= 12'b001011101101;
   7217: result <= 12'b001011101100;
   7218: result <= 12'b001011101011;
   7219: result <= 12'b001011101011;
   7220: result <= 12'b001011101010;
   7221: result <= 12'b001011101001;
   7222: result <= 12'b001011101000;
   7223: result <= 12'b001011101000;
   7224: result <= 12'b001011100111;
   7225: result <= 12'b001011100110;
   7226: result <= 12'b001011100101;
   7227: result <= 12'b001011100101;
   7228: result <= 12'b001011100100;
   7229: result <= 12'b001011100011;
   7230: result <= 12'b001011100011;
   7231: result <= 12'b001011100010;
   7232: result <= 12'b001011100001;
   7233: result <= 12'b001011100000;
   7234: result <= 12'b001011100000;
   7235: result <= 12'b001011011111;
   7236: result <= 12'b001011011110;
   7237: result <= 12'b001011011101;
   7238: result <= 12'b001011011101;
   7239: result <= 12'b001011011100;
   7240: result <= 12'b001011011011;
   7241: result <= 12'b001011011010;
   7242: result <= 12'b001011011010;
   7243: result <= 12'b001011011001;
   7244: result <= 12'b001011011000;
   7245: result <= 12'b001011011000;
   7246: result <= 12'b001011010111;
   7247: result <= 12'b001011010110;
   7248: result <= 12'b001011010101;
   7249: result <= 12'b001011010101;
   7250: result <= 12'b001011010100;
   7251: result <= 12'b001011010011;
   7252: result <= 12'b001011010010;
   7253: result <= 12'b001011010010;
   7254: result <= 12'b001011010001;
   7255: result <= 12'b001011010000;
   7256: result <= 12'b001011001111;
   7257: result <= 12'b001011001111;
   7258: result <= 12'b001011001110;
   7259: result <= 12'b001011001101;
   7260: result <= 12'b001011001101;
   7261: result <= 12'b001011001100;
   7262: result <= 12'b001011001011;
   7263: result <= 12'b001011001010;
   7264: result <= 12'b001011001010;
   7265: result <= 12'b001011001001;
   7266: result <= 12'b001011001000;
   7267: result <= 12'b001011000111;
   7268: result <= 12'b001011000111;
   7269: result <= 12'b001011000110;
   7270: result <= 12'b001011000101;
   7271: result <= 12'b001011000100;
   7272: result <= 12'b001011000100;
   7273: result <= 12'b001011000011;
   7274: result <= 12'b001011000010;
   7275: result <= 12'b001011000001;
   7276: result <= 12'b001011000001;
   7277: result <= 12'b001011000000;
   7278: result <= 12'b001010111111;
   7279: result <= 12'b001010111111;
   7280: result <= 12'b001010111110;
   7281: result <= 12'b001010111101;
   7282: result <= 12'b001010111100;
   7283: result <= 12'b001010111100;
   7284: result <= 12'b001010111011;
   7285: result <= 12'b001010111010;
   7286: result <= 12'b001010111001;
   7287: result <= 12'b001010111001;
   7288: result <= 12'b001010111000;
   7289: result <= 12'b001010110111;
   7290: result <= 12'b001010110110;
   7291: result <= 12'b001010110110;
   7292: result <= 12'b001010110101;
   7293: result <= 12'b001010110100;
   7294: result <= 12'b001010110011;
   7295: result <= 12'b001010110011;
   7296: result <= 12'b001010110010;
   7297: result <= 12'b001010110001;
   7298: result <= 12'b001010110000;
   7299: result <= 12'b001010110000;
   7300: result <= 12'b001010101111;
   7301: result <= 12'b001010101110;
   7302: result <= 12'b001010101110;
   7303: result <= 12'b001010101101;
   7304: result <= 12'b001010101100;
   7305: result <= 12'b001010101011;
   7306: result <= 12'b001010101011;
   7307: result <= 12'b001010101010;
   7308: result <= 12'b001010101001;
   7309: result <= 12'b001010101000;
   7310: result <= 12'b001010101000;
   7311: result <= 12'b001010100111;
   7312: result <= 12'b001010100110;
   7313: result <= 12'b001010100101;
   7314: result <= 12'b001010100101;
   7315: result <= 12'b001010100100;
   7316: result <= 12'b001010100011;
   7317: result <= 12'b001010100010;
   7318: result <= 12'b001010100010;
   7319: result <= 12'b001010100001;
   7320: result <= 12'b001010100000;
   7321: result <= 12'b001010011111;
   7322: result <= 12'b001010011111;
   7323: result <= 12'b001010011110;
   7324: result <= 12'b001010011101;
   7325: result <= 12'b001010011100;
   7326: result <= 12'b001010011100;
   7327: result <= 12'b001010011011;
   7328: result <= 12'b001010011010;
   7329: result <= 12'b001010011001;
   7330: result <= 12'b001010011001;
   7331: result <= 12'b001010011000;
   7332: result <= 12'b001010010111;
   7333: result <= 12'b001010010111;
   7334: result <= 12'b001010010110;
   7335: result <= 12'b001010010101;
   7336: result <= 12'b001010010100;
   7337: result <= 12'b001010010100;
   7338: result <= 12'b001010010011;
   7339: result <= 12'b001010010010;
   7340: result <= 12'b001010010001;
   7341: result <= 12'b001010010001;
   7342: result <= 12'b001010010000;
   7343: result <= 12'b001010001111;
   7344: result <= 12'b001010001110;
   7345: result <= 12'b001010001110;
   7346: result <= 12'b001010001101;
   7347: result <= 12'b001010001100;
   7348: result <= 12'b001010001011;
   7349: result <= 12'b001010001011;
   7350: result <= 12'b001010001010;
   7351: result <= 12'b001010001001;
   7352: result <= 12'b001010001000;
   7353: result <= 12'b001010001000;
   7354: result <= 12'b001010000111;
   7355: result <= 12'b001010000110;
   7356: result <= 12'b001010000101;
   7357: result <= 12'b001010000101;
   7358: result <= 12'b001010000100;
   7359: result <= 12'b001010000011;
   7360: result <= 12'b001010000010;
   7361: result <= 12'b001010000010;
   7362: result <= 12'b001010000001;
   7363: result <= 12'b001010000000;
   7364: result <= 12'b001001111111;
   7365: result <= 12'b001001111111;
   7366: result <= 12'b001001111110;
   7367: result <= 12'b001001111101;
   7368: result <= 12'b001001111100;
   7369: result <= 12'b001001111100;
   7370: result <= 12'b001001111011;
   7371: result <= 12'b001001111010;
   7372: result <= 12'b001001111001;
   7373: result <= 12'b001001111001;
   7374: result <= 12'b001001111000;
   7375: result <= 12'b001001110111;
   7376: result <= 12'b001001110110;
   7377: result <= 12'b001001110110;
   7378: result <= 12'b001001110101;
   7379: result <= 12'b001001110100;
   7380: result <= 12'b001001110011;
   7381: result <= 12'b001001110011;
   7382: result <= 12'b001001110010;
   7383: result <= 12'b001001110001;
   7384: result <= 12'b001001110000;
   7385: result <= 12'b001001110000;
   7386: result <= 12'b001001101111;
   7387: result <= 12'b001001101110;
   7388: result <= 12'b001001101110;
   7389: result <= 12'b001001101101;
   7390: result <= 12'b001001101100;
   7391: result <= 12'b001001101011;
   7392: result <= 12'b001001101011;
   7393: result <= 12'b001001101010;
   7394: result <= 12'b001001101001;
   7395: result <= 12'b001001101000;
   7396: result <= 12'b001001101000;
   7397: result <= 12'b001001100111;
   7398: result <= 12'b001001100110;
   7399: result <= 12'b001001100101;
   7400: result <= 12'b001001100101;
   7401: result <= 12'b001001100100;
   7402: result <= 12'b001001100011;
   7403: result <= 12'b001001100010;
   7404: result <= 12'b001001100010;
   7405: result <= 12'b001001100001;
   7406: result <= 12'b001001100000;
   7407: result <= 12'b001001011111;
   7408: result <= 12'b001001011111;
   7409: result <= 12'b001001011110;
   7410: result <= 12'b001001011101;
   7411: result <= 12'b001001011100;
   7412: result <= 12'b001001011100;
   7413: result <= 12'b001001011011;
   7414: result <= 12'b001001011010;
   7415: result <= 12'b001001011001;
   7416: result <= 12'b001001011001;
   7417: result <= 12'b001001011000;
   7418: result <= 12'b001001010111;
   7419: result <= 12'b001001010110;
   7420: result <= 12'b001001010110;
   7421: result <= 12'b001001010101;
   7422: result <= 12'b001001010100;
   7423: result <= 12'b001001010011;
   7424: result <= 12'b001001010011;
   7425: result <= 12'b001001010010;
   7426: result <= 12'b001001010001;
   7427: result <= 12'b001001010000;
   7428: result <= 12'b001001001111;
   7429: result <= 12'b001001001111;
   7430: result <= 12'b001001001110;
   7431: result <= 12'b001001001101;
   7432: result <= 12'b001001001100;
   7433: result <= 12'b001001001100;
   7434: result <= 12'b001001001011;
   7435: result <= 12'b001001001010;
   7436: result <= 12'b001001001001;
   7437: result <= 12'b001001001001;
   7438: result <= 12'b001001001000;
   7439: result <= 12'b001001000111;
   7440: result <= 12'b001001000110;
   7441: result <= 12'b001001000110;
   7442: result <= 12'b001001000101;
   7443: result <= 12'b001001000100;
   7444: result <= 12'b001001000011;
   7445: result <= 12'b001001000011;
   7446: result <= 12'b001001000010;
   7447: result <= 12'b001001000001;
   7448: result <= 12'b001001000000;
   7449: result <= 12'b001001000000;
   7450: result <= 12'b001000111111;
   7451: result <= 12'b001000111110;
   7452: result <= 12'b001000111101;
   7453: result <= 12'b001000111101;
   7454: result <= 12'b001000111100;
   7455: result <= 12'b001000111011;
   7456: result <= 12'b001000111010;
   7457: result <= 12'b001000111010;
   7458: result <= 12'b001000111001;
   7459: result <= 12'b001000111000;
   7460: result <= 12'b001000110111;
   7461: result <= 12'b001000110111;
   7462: result <= 12'b001000110110;
   7463: result <= 12'b001000110101;
   7464: result <= 12'b001000110100;
   7465: result <= 12'b001000110100;
   7466: result <= 12'b001000110011;
   7467: result <= 12'b001000110010;
   7468: result <= 12'b001000110001;
   7469: result <= 12'b001000110001;
   7470: result <= 12'b001000110000;
   7471: result <= 12'b001000101111;
   7472: result <= 12'b001000101110;
   7473: result <= 12'b001000101110;
   7474: result <= 12'b001000101101;
   7475: result <= 12'b001000101100;
   7476: result <= 12'b001000101011;
   7477: result <= 12'b001000101011;
   7478: result <= 12'b001000101010;
   7479: result <= 12'b001000101001;
   7480: result <= 12'b001000101000;
   7481: result <= 12'b001000101000;
   7482: result <= 12'b001000100111;
   7483: result <= 12'b001000100110;
   7484: result <= 12'b001000100101;
   7485: result <= 12'b001000100100;
   7486: result <= 12'b001000100100;
   7487: result <= 12'b001000100011;
   7488: result <= 12'b001000100010;
   7489: result <= 12'b001000100001;
   7490: result <= 12'b001000100001;
   7491: result <= 12'b001000100000;
   7492: result <= 12'b001000011111;
   7493: result <= 12'b001000011110;
   7494: result <= 12'b001000011110;
   7495: result <= 12'b001000011101;
   7496: result <= 12'b001000011100;
   7497: result <= 12'b001000011011;
   7498: result <= 12'b001000011011;
   7499: result <= 12'b001000011010;
   7500: result <= 12'b001000011001;
   7501: result <= 12'b001000011000;
   7502: result <= 12'b001000011000;
   7503: result <= 12'b001000010111;
   7504: result <= 12'b001000010110;
   7505: result <= 12'b001000010101;
   7506: result <= 12'b001000010101;
   7507: result <= 12'b001000010100;
   7508: result <= 12'b001000010011;
   7509: result <= 12'b001000010010;
   7510: result <= 12'b001000010010;
   7511: result <= 12'b001000010001;
   7512: result <= 12'b001000010000;
   7513: result <= 12'b001000001111;
   7514: result <= 12'b001000001111;
   7515: result <= 12'b001000001110;
   7516: result <= 12'b001000001101;
   7517: result <= 12'b001000001100;
   7518: result <= 12'b001000001011;
   7519: result <= 12'b001000001011;
   7520: result <= 12'b001000001010;
   7521: result <= 12'b001000001001;
   7522: result <= 12'b001000001000;
   7523: result <= 12'b001000001000;
   7524: result <= 12'b001000000111;
   7525: result <= 12'b001000000110;
   7526: result <= 12'b001000000101;
   7527: result <= 12'b001000000101;
   7528: result <= 12'b001000000100;
   7529: result <= 12'b001000000011;
   7530: result <= 12'b001000000010;
   7531: result <= 12'b001000000010;
   7532: result <= 12'b001000000001;
   7533: result <= 12'b001000000000;
   7534: result <= 12'b000111111111;
   7535: result <= 12'b000111111111;
   7536: result <= 12'b000111111110;
   7537: result <= 12'b000111111101;
   7538: result <= 12'b000111111100;
   7539: result <= 12'b000111111100;
   7540: result <= 12'b000111111011;
   7541: result <= 12'b000111111010;
   7542: result <= 12'b000111111001;
   7543: result <= 12'b000111111000;
   7544: result <= 12'b000111111000;
   7545: result <= 12'b000111110111;
   7546: result <= 12'b000111110110;
   7547: result <= 12'b000111110101;
   7548: result <= 12'b000111110101;
   7549: result <= 12'b000111110100;
   7550: result <= 12'b000111110011;
   7551: result <= 12'b000111110010;
   7552: result <= 12'b000111110010;
   7553: result <= 12'b000111110001;
   7554: result <= 12'b000111110000;
   7555: result <= 12'b000111101111;
   7556: result <= 12'b000111101111;
   7557: result <= 12'b000111101110;
   7558: result <= 12'b000111101101;
   7559: result <= 12'b000111101100;
   7560: result <= 12'b000111101100;
   7561: result <= 12'b000111101011;
   7562: result <= 12'b000111101010;
   7563: result <= 12'b000111101001;
   7564: result <= 12'b000111101000;
   7565: result <= 12'b000111101000;
   7566: result <= 12'b000111100111;
   7567: result <= 12'b000111100110;
   7568: result <= 12'b000111100101;
   7569: result <= 12'b000111100101;
   7570: result <= 12'b000111100100;
   7571: result <= 12'b000111100011;
   7572: result <= 12'b000111100010;
   7573: result <= 12'b000111100010;
   7574: result <= 12'b000111100001;
   7575: result <= 12'b000111100000;
   7576: result <= 12'b000111011111;
   7577: result <= 12'b000111011111;
   7578: result <= 12'b000111011110;
   7579: result <= 12'b000111011101;
   7580: result <= 12'b000111011100;
   7581: result <= 12'b000111011011;
   7582: result <= 12'b000111011011;
   7583: result <= 12'b000111011010;
   7584: result <= 12'b000111011001;
   7585: result <= 12'b000111011000;
   7586: result <= 12'b000111011000;
   7587: result <= 12'b000111010111;
   7588: result <= 12'b000111010110;
   7589: result <= 12'b000111010101;
   7590: result <= 12'b000111010101;
   7591: result <= 12'b000111010100;
   7592: result <= 12'b000111010011;
   7593: result <= 12'b000111010010;
   7594: result <= 12'b000111010010;
   7595: result <= 12'b000111010001;
   7596: result <= 12'b000111010000;
   7597: result <= 12'b000111001111;
   7598: result <= 12'b000111001111;
   7599: result <= 12'b000111001110;
   7600: result <= 12'b000111001101;
   7601: result <= 12'b000111001100;
   7602: result <= 12'b000111001011;
   7603: result <= 12'b000111001011;
   7604: result <= 12'b000111001010;
   7605: result <= 12'b000111001001;
   7606: result <= 12'b000111001000;
   7607: result <= 12'b000111001000;
   7608: result <= 12'b000111000111;
   7609: result <= 12'b000111000110;
   7610: result <= 12'b000111000101;
   7611: result <= 12'b000111000101;
   7612: result <= 12'b000111000100;
   7613: result <= 12'b000111000011;
   7614: result <= 12'b000111000010;
   7615: result <= 12'b000111000001;
   7616: result <= 12'b000111000001;
   7617: result <= 12'b000111000000;
   7618: result <= 12'b000110111111;
   7619: result <= 12'b000110111110;
   7620: result <= 12'b000110111110;
   7621: result <= 12'b000110111101;
   7622: result <= 12'b000110111100;
   7623: result <= 12'b000110111011;
   7624: result <= 12'b000110111011;
   7625: result <= 12'b000110111010;
   7626: result <= 12'b000110111001;
   7627: result <= 12'b000110111000;
   7628: result <= 12'b000110111000;
   7629: result <= 12'b000110110111;
   7630: result <= 12'b000110110110;
   7631: result <= 12'b000110110101;
   7632: result <= 12'b000110110100;
   7633: result <= 12'b000110110100;
   7634: result <= 12'b000110110011;
   7635: result <= 12'b000110110010;
   7636: result <= 12'b000110110001;
   7637: result <= 12'b000110110001;
   7638: result <= 12'b000110110000;
   7639: result <= 12'b000110101111;
   7640: result <= 12'b000110101110;
   7641: result <= 12'b000110101110;
   7642: result <= 12'b000110101101;
   7643: result <= 12'b000110101100;
   7644: result <= 12'b000110101011;
   7645: result <= 12'b000110101010;
   7646: result <= 12'b000110101010;
   7647: result <= 12'b000110101001;
   7648: result <= 12'b000110101000;
   7649: result <= 12'b000110100111;
   7650: result <= 12'b000110100111;
   7651: result <= 12'b000110100110;
   7652: result <= 12'b000110100101;
   7653: result <= 12'b000110100100;
   7654: result <= 12'b000110100100;
   7655: result <= 12'b000110100011;
   7656: result <= 12'b000110100010;
   7657: result <= 12'b000110100001;
   7658: result <= 12'b000110100000;
   7659: result <= 12'b000110100000;
   7660: result <= 12'b000110011111;
   7661: result <= 12'b000110011110;
   7662: result <= 12'b000110011101;
   7663: result <= 12'b000110011101;
   7664: result <= 12'b000110011100;
   7665: result <= 12'b000110011011;
   7666: result <= 12'b000110011010;
   7667: result <= 12'b000110011010;
   7668: result <= 12'b000110011001;
   7669: result <= 12'b000110011000;
   7670: result <= 12'b000110010111;
   7671: result <= 12'b000110010110;
   7672: result <= 12'b000110010110;
   7673: result <= 12'b000110010101;
   7674: result <= 12'b000110010100;
   7675: result <= 12'b000110010011;
   7676: result <= 12'b000110010011;
   7677: result <= 12'b000110010010;
   7678: result <= 12'b000110010001;
   7679: result <= 12'b000110010000;
   7680: result <= 12'b000110010000;
   7681: result <= 12'b000110001111;
   7682: result <= 12'b000110001110;
   7683: result <= 12'b000110001101;
   7684: result <= 12'b000110001100;
   7685: result <= 12'b000110001100;
   7686: result <= 12'b000110001011;
   7687: result <= 12'b000110001010;
   7688: result <= 12'b000110001001;
   7689: result <= 12'b000110001001;
   7690: result <= 12'b000110001000;
   7691: result <= 12'b000110000111;
   7692: result <= 12'b000110000110;
   7693: result <= 12'b000110000110;
   7694: result <= 12'b000110000101;
   7695: result <= 12'b000110000100;
   7696: result <= 12'b000110000011;
   7697: result <= 12'b000110000010;
   7698: result <= 12'b000110000010;
   7699: result <= 12'b000110000001;
   7700: result <= 12'b000110000000;
   7701: result <= 12'b000101111111;
   7702: result <= 12'b000101111111;
   7703: result <= 12'b000101111110;
   7704: result <= 12'b000101111101;
   7705: result <= 12'b000101111100;
   7706: result <= 12'b000101111011;
   7707: result <= 12'b000101111011;
   7708: result <= 12'b000101111010;
   7709: result <= 12'b000101111001;
   7710: result <= 12'b000101111000;
   7711: result <= 12'b000101111000;
   7712: result <= 12'b000101110111;
   7713: result <= 12'b000101110110;
   7714: result <= 12'b000101110101;
   7715: result <= 12'b000101110101;
   7716: result <= 12'b000101110100;
   7717: result <= 12'b000101110011;
   7718: result <= 12'b000101110010;
   7719: result <= 12'b000101110001;
   7720: result <= 12'b000101110001;
   7721: result <= 12'b000101110000;
   7722: result <= 12'b000101101111;
   7723: result <= 12'b000101101110;
   7724: result <= 12'b000101101110;
   7725: result <= 12'b000101101101;
   7726: result <= 12'b000101101100;
   7727: result <= 12'b000101101011;
   7728: result <= 12'b000101101011;
   7729: result <= 12'b000101101010;
   7730: result <= 12'b000101101001;
   7731: result <= 12'b000101101000;
   7732: result <= 12'b000101100111;
   7733: result <= 12'b000101100111;
   7734: result <= 12'b000101100110;
   7735: result <= 12'b000101100101;
   7736: result <= 12'b000101100100;
   7737: result <= 12'b000101100100;
   7738: result <= 12'b000101100011;
   7739: result <= 12'b000101100010;
   7740: result <= 12'b000101100001;
   7741: result <= 12'b000101100000;
   7742: result <= 12'b000101100000;
   7743: result <= 12'b000101011111;
   7744: result <= 12'b000101011110;
   7745: result <= 12'b000101011101;
   7746: result <= 12'b000101011101;
   7747: result <= 12'b000101011100;
   7748: result <= 12'b000101011011;
   7749: result <= 12'b000101011010;
   7750: result <= 12'b000101011001;
   7751: result <= 12'b000101011001;
   7752: result <= 12'b000101011000;
   7753: result <= 12'b000101010111;
   7754: result <= 12'b000101010110;
   7755: result <= 12'b000101010110;
   7756: result <= 12'b000101010101;
   7757: result <= 12'b000101010100;
   7758: result <= 12'b000101010011;
   7759: result <= 12'b000101010011;
   7760: result <= 12'b000101010010;
   7761: result <= 12'b000101010001;
   7762: result <= 12'b000101010000;
   7763: result <= 12'b000101001111;
   7764: result <= 12'b000101001111;
   7765: result <= 12'b000101001110;
   7766: result <= 12'b000101001101;
   7767: result <= 12'b000101001100;
   7768: result <= 12'b000101001100;
   7769: result <= 12'b000101001011;
   7770: result <= 12'b000101001010;
   7771: result <= 12'b000101001001;
   7772: result <= 12'b000101001000;
   7773: result <= 12'b000101001000;
   7774: result <= 12'b000101000111;
   7775: result <= 12'b000101000110;
   7776: result <= 12'b000101000101;
   7777: result <= 12'b000101000101;
   7778: result <= 12'b000101000100;
   7779: result <= 12'b000101000011;
   7780: result <= 12'b000101000010;
   7781: result <= 12'b000101000001;
   7782: result <= 12'b000101000001;
   7783: result <= 12'b000101000000;
   7784: result <= 12'b000100111111;
   7785: result <= 12'b000100111110;
   7786: result <= 12'b000100111110;
   7787: result <= 12'b000100111101;
   7788: result <= 12'b000100111100;
   7789: result <= 12'b000100111011;
   7790: result <= 12'b000100111010;
   7791: result <= 12'b000100111010;
   7792: result <= 12'b000100111001;
   7793: result <= 12'b000100111000;
   7794: result <= 12'b000100110111;
   7795: result <= 12'b000100110111;
   7796: result <= 12'b000100110110;
   7797: result <= 12'b000100110101;
   7798: result <= 12'b000100110100;
   7799: result <= 12'b000100110011;
   7800: result <= 12'b000100110011;
   7801: result <= 12'b000100110010;
   7802: result <= 12'b000100110001;
   7803: result <= 12'b000100110000;
   7804: result <= 12'b000100110000;
   7805: result <= 12'b000100101111;
   7806: result <= 12'b000100101110;
   7807: result <= 12'b000100101101;
   7808: result <= 12'b000100101101;
   7809: result <= 12'b000100101100;
   7810: result <= 12'b000100101011;
   7811: result <= 12'b000100101010;
   7812: result <= 12'b000100101001;
   7813: result <= 12'b000100101001;
   7814: result <= 12'b000100101000;
   7815: result <= 12'b000100100111;
   7816: result <= 12'b000100100110;
   7817: result <= 12'b000100100110;
   7818: result <= 12'b000100100101;
   7819: result <= 12'b000100100100;
   7820: result <= 12'b000100100011;
   7821: result <= 12'b000100100010;
   7822: result <= 12'b000100100010;
   7823: result <= 12'b000100100001;
   7824: result <= 12'b000100100000;
   7825: result <= 12'b000100011111;
   7826: result <= 12'b000100011111;
   7827: result <= 12'b000100011110;
   7828: result <= 12'b000100011101;
   7829: result <= 12'b000100011100;
   7830: result <= 12'b000100011011;
   7831: result <= 12'b000100011011;
   7832: result <= 12'b000100011010;
   7833: result <= 12'b000100011001;
   7834: result <= 12'b000100011000;
   7835: result <= 12'b000100011000;
   7836: result <= 12'b000100010111;
   7837: result <= 12'b000100010110;
   7838: result <= 12'b000100010101;
   7839: result <= 12'b000100010100;
   7840: result <= 12'b000100010100;
   7841: result <= 12'b000100010011;
   7842: result <= 12'b000100010010;
   7843: result <= 12'b000100010001;
   7844: result <= 12'b000100010001;
   7845: result <= 12'b000100010000;
   7846: result <= 12'b000100001111;
   7847: result <= 12'b000100001110;
   7848: result <= 12'b000100001101;
   7849: result <= 12'b000100001101;
   7850: result <= 12'b000100001100;
   7851: result <= 12'b000100001011;
   7852: result <= 12'b000100001010;
   7853: result <= 12'b000100001010;
   7854: result <= 12'b000100001001;
   7855: result <= 12'b000100001000;
   7856: result <= 12'b000100000111;
   7857: result <= 12'b000100000110;
   7858: result <= 12'b000100000110;
   7859: result <= 12'b000100000101;
   7860: result <= 12'b000100000100;
   7861: result <= 12'b000100000011;
   7862: result <= 12'b000100000010;
   7863: result <= 12'b000100000010;
   7864: result <= 12'b000100000001;
   7865: result <= 12'b000100000000;
   7866: result <= 12'b000011111111;
   7867: result <= 12'b000011111111;
   7868: result <= 12'b000011111110;
   7869: result <= 12'b000011111101;
   7870: result <= 12'b000011111100;
   7871: result <= 12'b000011111011;
   7872: result <= 12'b000011111011;
   7873: result <= 12'b000011111010;
   7874: result <= 12'b000011111001;
   7875: result <= 12'b000011111000;
   7876: result <= 12'b000011111000;
   7877: result <= 12'b000011110111;
   7878: result <= 12'b000011110110;
   7879: result <= 12'b000011110101;
   7880: result <= 12'b000011110100;
   7881: result <= 12'b000011110100;
   7882: result <= 12'b000011110011;
   7883: result <= 12'b000011110010;
   7884: result <= 12'b000011110001;
   7885: result <= 12'b000011110001;
   7886: result <= 12'b000011110000;
   7887: result <= 12'b000011101111;
   7888: result <= 12'b000011101110;
   7889: result <= 12'b000011101101;
   7890: result <= 12'b000011101101;
   7891: result <= 12'b000011101100;
   7892: result <= 12'b000011101011;
   7893: result <= 12'b000011101010;
   7894: result <= 12'b000011101010;
   7895: result <= 12'b000011101001;
   7896: result <= 12'b000011101000;
   7897: result <= 12'b000011100111;
   7898: result <= 12'b000011100110;
   7899: result <= 12'b000011100110;
   7900: result <= 12'b000011100101;
   7901: result <= 12'b000011100100;
   7902: result <= 12'b000011100011;
   7903: result <= 12'b000011100011;
   7904: result <= 12'b000011100010;
   7905: result <= 12'b000011100001;
   7906: result <= 12'b000011100000;
   7907: result <= 12'b000011011111;
   7908: result <= 12'b000011011111;
   7909: result <= 12'b000011011110;
   7910: result <= 12'b000011011101;
   7911: result <= 12'b000011011100;
   7912: result <= 12'b000011011011;
   7913: result <= 12'b000011011011;
   7914: result <= 12'b000011011010;
   7915: result <= 12'b000011011001;
   7916: result <= 12'b000011011000;
   7917: result <= 12'b000011011000;
   7918: result <= 12'b000011010111;
   7919: result <= 12'b000011010110;
   7920: result <= 12'b000011010101;
   7921: result <= 12'b000011010100;
   7922: result <= 12'b000011010100;
   7923: result <= 12'b000011010011;
   7924: result <= 12'b000011010010;
   7925: result <= 12'b000011010001;
   7926: result <= 12'b000011010001;
   7927: result <= 12'b000011010000;
   7928: result <= 12'b000011001111;
   7929: result <= 12'b000011001110;
   7930: result <= 12'b000011001101;
   7931: result <= 12'b000011001101;
   7932: result <= 12'b000011001100;
   7933: result <= 12'b000011001011;
   7934: result <= 12'b000011001010;
   7935: result <= 12'b000011001010;
   7936: result <= 12'b000011001001;
   7937: result <= 12'b000011001000;
   7938: result <= 12'b000011000111;
   7939: result <= 12'b000011000110;
   7940: result <= 12'b000011000110;
   7941: result <= 12'b000011000101;
   7942: result <= 12'b000011000100;
   7943: result <= 12'b000011000011;
   7944: result <= 12'b000011000010;
   7945: result <= 12'b000011000010;
   7946: result <= 12'b000011000001;
   7947: result <= 12'b000011000000;
   7948: result <= 12'b000010111111;
   7949: result <= 12'b000010111111;
   7950: result <= 12'b000010111110;
   7951: result <= 12'b000010111101;
   7952: result <= 12'b000010111100;
   7953: result <= 12'b000010111011;
   7954: result <= 12'b000010111011;
   7955: result <= 12'b000010111010;
   7956: result <= 12'b000010111001;
   7957: result <= 12'b000010111000;
   7958: result <= 12'b000010111000;
   7959: result <= 12'b000010110111;
   7960: result <= 12'b000010110110;
   7961: result <= 12'b000010110101;
   7962: result <= 12'b000010110100;
   7963: result <= 12'b000010110100;
   7964: result <= 12'b000010110011;
   7965: result <= 12'b000010110010;
   7966: result <= 12'b000010110001;
   7967: result <= 12'b000010110000;
   7968: result <= 12'b000010110000;
   7969: result <= 12'b000010101111;
   7970: result <= 12'b000010101110;
   7971: result <= 12'b000010101101;
   7972: result <= 12'b000010101101;
   7973: result <= 12'b000010101100;
   7974: result <= 12'b000010101011;
   7975: result <= 12'b000010101010;
   7976: result <= 12'b000010101001;
   7977: result <= 12'b000010101001;
   7978: result <= 12'b000010101000;
   7979: result <= 12'b000010100111;
   7980: result <= 12'b000010100110;
   7981: result <= 12'b000010100110;
   7982: result <= 12'b000010100101;
   7983: result <= 12'b000010100100;
   7984: result <= 12'b000010100011;
   7985: result <= 12'b000010100010;
   7986: result <= 12'b000010100010;
   7987: result <= 12'b000010100001;
   7988: result <= 12'b000010100000;
   7989: result <= 12'b000010011111;
   7990: result <= 12'b000010011110;
   7991: result <= 12'b000010011110;
   7992: result <= 12'b000010011101;
   7993: result <= 12'b000010011100;
   7994: result <= 12'b000010011011;
   7995: result <= 12'b000010011011;
   7996: result <= 12'b000010011010;
   7997: result <= 12'b000010011001;
   7998: result <= 12'b000010011000;
   7999: result <= 12'b000010010111;
   8000: result <= 12'b000010010111;
   8001: result <= 12'b000010010110;
   8002: result <= 12'b000010010101;
   8003: result <= 12'b000010010100;
   8004: result <= 12'b000010010100;
   8005: result <= 12'b000010010011;
   8006: result <= 12'b000010010010;
   8007: result <= 12'b000010010001;
   8008: result <= 12'b000010010000;
   8009: result <= 12'b000010010000;
   8010: result <= 12'b000010001111;
   8011: result <= 12'b000010001110;
   8012: result <= 12'b000010001101;
   8013: result <= 12'b000010001100;
   8014: result <= 12'b000010001100;
   8015: result <= 12'b000010001011;
   8016: result <= 12'b000010001010;
   8017: result <= 12'b000010001001;
   8018: result <= 12'b000010001001;
   8019: result <= 12'b000010001000;
   8020: result <= 12'b000010000111;
   8021: result <= 12'b000010000110;
   8022: result <= 12'b000010000101;
   8023: result <= 12'b000010000101;
   8024: result <= 12'b000010000100;
   8025: result <= 12'b000010000011;
   8026: result <= 12'b000010000010;
   8027: result <= 12'b000010000010;
   8028: result <= 12'b000010000001;
   8029: result <= 12'b000010000000;
   8030: result <= 12'b000001111111;
   8031: result <= 12'b000001111110;
   8032: result <= 12'b000001111110;
   8033: result <= 12'b000001111101;
   8034: result <= 12'b000001111100;
   8035: result <= 12'b000001111011;
   8036: result <= 12'b000001111010;
   8037: result <= 12'b000001111010;
   8038: result <= 12'b000001111001;
   8039: result <= 12'b000001111000;
   8040: result <= 12'b000001110111;
   8041: result <= 12'b000001110111;
   8042: result <= 12'b000001110110;
   8043: result <= 12'b000001110101;
   8044: result <= 12'b000001110100;
   8045: result <= 12'b000001110011;
   8046: result <= 12'b000001110011;
   8047: result <= 12'b000001110010;
   8048: result <= 12'b000001110001;
   8049: result <= 12'b000001110000;
   8050: result <= 12'b000001101111;
   8051: result <= 12'b000001101111;
   8052: result <= 12'b000001101110;
   8053: result <= 12'b000001101101;
   8054: result <= 12'b000001101100;
   8055: result <= 12'b000001101100;
   8056: result <= 12'b000001101011;
   8057: result <= 12'b000001101010;
   8058: result <= 12'b000001101001;
   8059: result <= 12'b000001101000;
   8060: result <= 12'b000001101000;
   8061: result <= 12'b000001100111;
   8062: result <= 12'b000001100110;
   8063: result <= 12'b000001100101;
   8064: result <= 12'b000001100100;
   8065: result <= 12'b000001100100;
   8066: result <= 12'b000001100011;
   8067: result <= 12'b000001100010;
   8068: result <= 12'b000001100001;
   8069: result <= 12'b000001100001;
   8070: result <= 12'b000001100000;
   8071: result <= 12'b000001011111;
   8072: result <= 12'b000001011110;
   8073: result <= 12'b000001011101;
   8074: result <= 12'b000001011101;
   8075: result <= 12'b000001011100;
   8076: result <= 12'b000001011011;
   8077: result <= 12'b000001011010;
   8078: result <= 12'b000001011010;
   8079: result <= 12'b000001011001;
   8080: result <= 12'b000001011000;
   8081: result <= 12'b000001010111;
   8082: result <= 12'b000001010110;
   8083: result <= 12'b000001010110;
   8084: result <= 12'b000001010101;
   8085: result <= 12'b000001010100;
   8086: result <= 12'b000001010011;
   8087: result <= 12'b000001010010;
   8088: result <= 12'b000001010010;
   8089: result <= 12'b000001010001;
   8090: result <= 12'b000001010000;
   8091: result <= 12'b000001001111;
   8092: result <= 12'b000001001111;
   8093: result <= 12'b000001001110;
   8094: result <= 12'b000001001101;
   8095: result <= 12'b000001001100;
   8096: result <= 12'b000001001011;
   8097: result <= 12'b000001001011;
   8098: result <= 12'b000001001010;
   8099: result <= 12'b000001001001;
   8100: result <= 12'b000001001000;
   8101: result <= 12'b000001000111;
   8102: result <= 12'b000001000111;
   8103: result <= 12'b000001000110;
   8104: result <= 12'b000001000101;
   8105: result <= 12'b000001000100;
   8106: result <= 12'b000001000100;
   8107: result <= 12'b000001000011;
   8108: result <= 12'b000001000010;
   8109: result <= 12'b000001000001;
   8110: result <= 12'b000001000000;
   8111: result <= 12'b000001000000;
   8112: result <= 12'b000000111111;
   8113: result <= 12'b000000111110;
   8114: result <= 12'b000000111101;
   8115: result <= 12'b000000111100;
   8116: result <= 12'b000000111100;
   8117: result <= 12'b000000111011;
   8118: result <= 12'b000000111010;
   8119: result <= 12'b000000111001;
   8120: result <= 12'b000000111001;
   8121: result <= 12'b000000111000;
   8122: result <= 12'b000000110111;
   8123: result <= 12'b000000110110;
   8124: result <= 12'b000000110101;
   8125: result <= 12'b000000110101;
   8126: result <= 12'b000000110100;
   8127: result <= 12'b000000110011;
   8128: result <= 12'b000000110010;
   8129: result <= 12'b000000110001;
   8130: result <= 12'b000000110001;
   8131: result <= 12'b000000110000;
   8132: result <= 12'b000000101111;
   8133: result <= 12'b000000101110;
   8134: result <= 12'b000000101110;
   8135: result <= 12'b000000101101;
   8136: result <= 12'b000000101100;
   8137: result <= 12'b000000101011;
   8138: result <= 12'b000000101010;
   8139: result <= 12'b000000101010;
   8140: result <= 12'b000000101001;
   8141: result <= 12'b000000101000;
   8142: result <= 12'b000000100111;
   8143: result <= 12'b000000100110;
   8144: result <= 12'b000000100110;
   8145: result <= 12'b000000100101;
   8146: result <= 12'b000000100100;
   8147: result <= 12'b000000100011;
   8148: result <= 12'b000000100011;
   8149: result <= 12'b000000100010;
   8150: result <= 12'b000000100001;
   8151: result <= 12'b000000100000;
   8152: result <= 12'b000000011111;
   8153: result <= 12'b000000011111;
   8154: result <= 12'b000000011110;
   8155: result <= 12'b000000011101;
   8156: result <= 12'b000000011100;
   8157: result <= 12'b000000011011;
   8158: result <= 12'b000000011011;
   8159: result <= 12'b000000011010;
   8160: result <= 12'b000000011001;
   8161: result <= 12'b000000011000;
   8162: result <= 12'b000000011000;
   8163: result <= 12'b000000010111;
   8164: result <= 12'b000000010110;
   8165: result <= 12'b000000010101;
   8166: result <= 12'b000000010100;
   8167: result <= 12'b000000010100;
   8168: result <= 12'b000000010011;
   8169: result <= 12'b000000010010;
   8170: result <= 12'b000000010001;
   8171: result <= 12'b000000010000;
   8172: result <= 12'b000000010000;
   8173: result <= 12'b000000001111;
   8174: result <= 12'b000000001110;
   8175: result <= 12'b000000001101;
   8176: result <= 12'b000000001101;
   8177: result <= 12'b000000001100;
   8178: result <= 12'b000000001011;
   8179: result <= 12'b000000001010;
   8180: result <= 12'b000000001001;
   8181: result <= 12'b000000001001;
   8182: result <= 12'b000000001000;
   8183: result <= 12'b000000000111;
   8184: result <= 12'b000000000110;
   8185: result <= 12'b000000000101;
   8186: result <= 12'b000000000101;
   8187: result <= 12'b000000000100;
   8188: result <= 12'b000000000011;
   8189: result <= 12'b000000000010;
   8190: result <= 12'b000000000010;
   8191: result <= 12'b000000000001;
   8192: result <= 12'b000000000000;
   8193: result <= 12'b111111111111;
   8194: result <= 12'b111111111110;
   8195: result <= 12'b111111111110;
   8196: result <= 12'b111111111101;
   8197: result <= 12'b111111111100;
   8198: result <= 12'b111111111011;
   8199: result <= 12'b111111111011;
   8200: result <= 12'b111111111010;
   8201: result <= 12'b111111111001;
   8202: result <= 12'b111111111000;
   8203: result <= 12'b111111110111;
   8204: result <= 12'b111111110111;
   8205: result <= 12'b111111110110;
   8206: result <= 12'b111111110101;
   8207: result <= 12'b111111110100;
   8208: result <= 12'b111111110011;
   8209: result <= 12'b111111110011;
   8210: result <= 12'b111111110010;
   8211: result <= 12'b111111110001;
   8212: result <= 12'b111111110000;
   8213: result <= 12'b111111110000;
   8214: result <= 12'b111111101111;
   8215: result <= 12'b111111101110;
   8216: result <= 12'b111111101101;
   8217: result <= 12'b111111101100;
   8218: result <= 12'b111111101100;
   8219: result <= 12'b111111101011;
   8220: result <= 12'b111111101010;
   8221: result <= 12'b111111101001;
   8222: result <= 12'b111111101000;
   8223: result <= 12'b111111101000;
   8224: result <= 12'b111111100111;
   8225: result <= 12'b111111100110;
   8226: result <= 12'b111111100101;
   8227: result <= 12'b111111100101;
   8228: result <= 12'b111111100100;
   8229: result <= 12'b111111100011;
   8230: result <= 12'b111111100010;
   8231: result <= 12'b111111100001;
   8232: result <= 12'b111111100001;
   8233: result <= 12'b111111100000;
   8234: result <= 12'b111111011111;
   8235: result <= 12'b111111011110;
   8236: result <= 12'b111111011101;
   8237: result <= 12'b111111011101;
   8238: result <= 12'b111111011100;
   8239: result <= 12'b111111011011;
   8240: result <= 12'b111111011010;
   8241: result <= 12'b111111011010;
   8242: result <= 12'b111111011001;
   8243: result <= 12'b111111011000;
   8244: result <= 12'b111111010111;
   8245: result <= 12'b111111010110;
   8246: result <= 12'b111111010110;
   8247: result <= 12'b111111010101;
   8248: result <= 12'b111111010100;
   8249: result <= 12'b111111010011;
   8250: result <= 12'b111111010010;
   8251: result <= 12'b111111010010;
   8252: result <= 12'b111111010001;
   8253: result <= 12'b111111010000;
   8254: result <= 12'b111111001111;
   8255: result <= 12'b111111001111;
   8256: result <= 12'b111111001110;
   8257: result <= 12'b111111001101;
   8258: result <= 12'b111111001100;
   8259: result <= 12'b111111001011;
   8260: result <= 12'b111111001011;
   8261: result <= 12'b111111001010;
   8262: result <= 12'b111111001001;
   8263: result <= 12'b111111001000;
   8264: result <= 12'b111111000111;
   8265: result <= 12'b111111000111;
   8266: result <= 12'b111111000110;
   8267: result <= 12'b111111000101;
   8268: result <= 12'b111111000100;
   8269: result <= 12'b111111000100;
   8270: result <= 12'b111111000011;
   8271: result <= 12'b111111000010;
   8272: result <= 12'b111111000001;
   8273: result <= 12'b111111000000;
   8274: result <= 12'b111111000000;
   8275: result <= 12'b111110111111;
   8276: result <= 12'b111110111110;
   8277: result <= 12'b111110111101;
   8278: result <= 12'b111110111100;
   8279: result <= 12'b111110111100;
   8280: result <= 12'b111110111011;
   8281: result <= 12'b111110111010;
   8282: result <= 12'b111110111001;
   8283: result <= 12'b111110111001;
   8284: result <= 12'b111110111000;
   8285: result <= 12'b111110110111;
   8286: result <= 12'b111110110110;
   8287: result <= 12'b111110110101;
   8288: result <= 12'b111110110101;
   8289: result <= 12'b111110110100;
   8290: result <= 12'b111110110011;
   8291: result <= 12'b111110110010;
   8292: result <= 12'b111110110001;
   8293: result <= 12'b111110110001;
   8294: result <= 12'b111110110000;
   8295: result <= 12'b111110101111;
   8296: result <= 12'b111110101110;
   8297: result <= 12'b111110101110;
   8298: result <= 12'b111110101101;
   8299: result <= 12'b111110101100;
   8300: result <= 12'b111110101011;
   8301: result <= 12'b111110101010;
   8302: result <= 12'b111110101010;
   8303: result <= 12'b111110101001;
   8304: result <= 12'b111110101000;
   8305: result <= 12'b111110100111;
   8306: result <= 12'b111110100110;
   8307: result <= 12'b111110100110;
   8308: result <= 12'b111110100101;
   8309: result <= 12'b111110100100;
   8310: result <= 12'b111110100011;
   8311: result <= 12'b111110100011;
   8312: result <= 12'b111110100010;
   8313: result <= 12'b111110100001;
   8314: result <= 12'b111110100000;
   8315: result <= 12'b111110011111;
   8316: result <= 12'b111110011111;
   8317: result <= 12'b111110011110;
   8318: result <= 12'b111110011101;
   8319: result <= 12'b111110011100;
   8320: result <= 12'b111110011100;
   8321: result <= 12'b111110011011;
   8322: result <= 12'b111110011010;
   8323: result <= 12'b111110011001;
   8324: result <= 12'b111110011000;
   8325: result <= 12'b111110011000;
   8326: result <= 12'b111110010111;
   8327: result <= 12'b111110010110;
   8328: result <= 12'b111110010101;
   8329: result <= 12'b111110010100;
   8330: result <= 12'b111110010100;
   8331: result <= 12'b111110010011;
   8332: result <= 12'b111110010010;
   8333: result <= 12'b111110010001;
   8334: result <= 12'b111110010001;
   8335: result <= 12'b111110010000;
   8336: result <= 12'b111110001111;
   8337: result <= 12'b111110001110;
   8338: result <= 12'b111110001101;
   8339: result <= 12'b111110001101;
   8340: result <= 12'b111110001100;
   8341: result <= 12'b111110001011;
   8342: result <= 12'b111110001010;
   8343: result <= 12'b111110001001;
   8344: result <= 12'b111110001001;
   8345: result <= 12'b111110001000;
   8346: result <= 12'b111110000111;
   8347: result <= 12'b111110000110;
   8348: result <= 12'b111110000110;
   8349: result <= 12'b111110000101;
   8350: result <= 12'b111110000100;
   8351: result <= 12'b111110000011;
   8352: result <= 12'b111110000010;
   8353: result <= 12'b111110000010;
   8354: result <= 12'b111110000001;
   8355: result <= 12'b111110000000;
   8356: result <= 12'b111101111111;
   8357: result <= 12'b111101111110;
   8358: result <= 12'b111101111110;
   8359: result <= 12'b111101111101;
   8360: result <= 12'b111101111100;
   8361: result <= 12'b111101111011;
   8362: result <= 12'b111101111011;
   8363: result <= 12'b111101111010;
   8364: result <= 12'b111101111001;
   8365: result <= 12'b111101111000;
   8366: result <= 12'b111101110111;
   8367: result <= 12'b111101110111;
   8368: result <= 12'b111101110110;
   8369: result <= 12'b111101110101;
   8370: result <= 12'b111101110100;
   8371: result <= 12'b111101110100;
   8372: result <= 12'b111101110011;
   8373: result <= 12'b111101110010;
   8374: result <= 12'b111101110001;
   8375: result <= 12'b111101110000;
   8376: result <= 12'b111101110000;
   8377: result <= 12'b111101101111;
   8378: result <= 12'b111101101110;
   8379: result <= 12'b111101101101;
   8380: result <= 12'b111101101100;
   8381: result <= 12'b111101101100;
   8382: result <= 12'b111101101011;
   8383: result <= 12'b111101101010;
   8384: result <= 12'b111101101001;
   8385: result <= 12'b111101101001;
   8386: result <= 12'b111101101000;
   8387: result <= 12'b111101100111;
   8388: result <= 12'b111101100110;
   8389: result <= 12'b111101100101;
   8390: result <= 12'b111101100101;
   8391: result <= 12'b111101100100;
   8392: result <= 12'b111101100011;
   8393: result <= 12'b111101100010;
   8394: result <= 12'b111101100010;
   8395: result <= 12'b111101100001;
   8396: result <= 12'b111101100000;
   8397: result <= 12'b111101011111;
   8398: result <= 12'b111101011110;
   8399: result <= 12'b111101011110;
   8400: result <= 12'b111101011101;
   8401: result <= 12'b111101011100;
   8402: result <= 12'b111101011011;
   8403: result <= 12'b111101011010;
   8404: result <= 12'b111101011010;
   8405: result <= 12'b111101011001;
   8406: result <= 12'b111101011000;
   8407: result <= 12'b111101010111;
   8408: result <= 12'b111101010111;
   8409: result <= 12'b111101010110;
   8410: result <= 12'b111101010101;
   8411: result <= 12'b111101010100;
   8412: result <= 12'b111101010011;
   8413: result <= 12'b111101010011;
   8414: result <= 12'b111101010010;
   8415: result <= 12'b111101010001;
   8416: result <= 12'b111101010000;
   8417: result <= 12'b111101010000;
   8418: result <= 12'b111101001111;
   8419: result <= 12'b111101001110;
   8420: result <= 12'b111101001101;
   8421: result <= 12'b111101001100;
   8422: result <= 12'b111101001100;
   8423: result <= 12'b111101001011;
   8424: result <= 12'b111101001010;
   8425: result <= 12'b111101001001;
   8426: result <= 12'b111101001000;
   8427: result <= 12'b111101001000;
   8428: result <= 12'b111101000111;
   8429: result <= 12'b111101000110;
   8430: result <= 12'b111101000101;
   8431: result <= 12'b111101000101;
   8432: result <= 12'b111101000100;
   8433: result <= 12'b111101000011;
   8434: result <= 12'b111101000010;
   8435: result <= 12'b111101000001;
   8436: result <= 12'b111101000001;
   8437: result <= 12'b111101000000;
   8438: result <= 12'b111100111111;
   8439: result <= 12'b111100111110;
   8440: result <= 12'b111100111110;
   8441: result <= 12'b111100111101;
   8442: result <= 12'b111100111100;
   8443: result <= 12'b111100111011;
   8444: result <= 12'b111100111010;
   8445: result <= 12'b111100111010;
   8446: result <= 12'b111100111001;
   8447: result <= 12'b111100111000;
   8448: result <= 12'b111100110111;
   8449: result <= 12'b111100110110;
   8450: result <= 12'b111100110110;
   8451: result <= 12'b111100110101;
   8452: result <= 12'b111100110100;
   8453: result <= 12'b111100110011;
   8454: result <= 12'b111100110011;
   8455: result <= 12'b111100110010;
   8456: result <= 12'b111100110001;
   8457: result <= 12'b111100110000;
   8458: result <= 12'b111100101111;
   8459: result <= 12'b111100101111;
   8460: result <= 12'b111100101110;
   8461: result <= 12'b111100101101;
   8462: result <= 12'b111100101100;
   8463: result <= 12'b111100101100;
   8464: result <= 12'b111100101011;
   8465: result <= 12'b111100101010;
   8466: result <= 12'b111100101001;
   8467: result <= 12'b111100101000;
   8468: result <= 12'b111100101000;
   8469: result <= 12'b111100100111;
   8470: result <= 12'b111100100110;
   8471: result <= 12'b111100100101;
   8472: result <= 12'b111100100101;
   8473: result <= 12'b111100100100;
   8474: result <= 12'b111100100011;
   8475: result <= 12'b111100100010;
   8476: result <= 12'b111100100001;
   8477: result <= 12'b111100100001;
   8478: result <= 12'b111100100000;
   8479: result <= 12'b111100011111;
   8480: result <= 12'b111100011110;
   8481: result <= 12'b111100011101;
   8482: result <= 12'b111100011101;
   8483: result <= 12'b111100011100;
   8484: result <= 12'b111100011011;
   8485: result <= 12'b111100011010;
   8486: result <= 12'b111100011010;
   8487: result <= 12'b111100011001;
   8488: result <= 12'b111100011000;
   8489: result <= 12'b111100010111;
   8490: result <= 12'b111100010110;
   8491: result <= 12'b111100010110;
   8492: result <= 12'b111100010101;
   8493: result <= 12'b111100010100;
   8494: result <= 12'b111100010011;
   8495: result <= 12'b111100010011;
   8496: result <= 12'b111100010010;
   8497: result <= 12'b111100010001;
   8498: result <= 12'b111100010000;
   8499: result <= 12'b111100001111;
   8500: result <= 12'b111100001111;
   8501: result <= 12'b111100001110;
   8502: result <= 12'b111100001101;
   8503: result <= 12'b111100001100;
   8504: result <= 12'b111100001100;
   8505: result <= 12'b111100001011;
   8506: result <= 12'b111100001010;
   8507: result <= 12'b111100001001;
   8508: result <= 12'b111100001000;
   8509: result <= 12'b111100001000;
   8510: result <= 12'b111100000111;
   8511: result <= 12'b111100000110;
   8512: result <= 12'b111100000101;
   8513: result <= 12'b111100000101;
   8514: result <= 12'b111100000100;
   8515: result <= 12'b111100000011;
   8516: result <= 12'b111100000010;
   8517: result <= 12'b111100000001;
   8518: result <= 12'b111100000001;
   8519: result <= 12'b111100000000;
   8520: result <= 12'b111011111111;
   8521: result <= 12'b111011111110;
   8522: result <= 12'b111011111110;
   8523: result <= 12'b111011111101;
   8524: result <= 12'b111011111100;
   8525: result <= 12'b111011111011;
   8526: result <= 12'b111011111010;
   8527: result <= 12'b111011111010;
   8528: result <= 12'b111011111001;
   8529: result <= 12'b111011111000;
   8530: result <= 12'b111011110111;
   8531: result <= 12'b111011110110;
   8532: result <= 12'b111011110110;
   8533: result <= 12'b111011110101;
   8534: result <= 12'b111011110100;
   8535: result <= 12'b111011110011;
   8536: result <= 12'b111011110011;
   8537: result <= 12'b111011110010;
   8538: result <= 12'b111011110001;
   8539: result <= 12'b111011110000;
   8540: result <= 12'b111011101111;
   8541: result <= 12'b111011101111;
   8542: result <= 12'b111011101110;
   8543: result <= 12'b111011101101;
   8544: result <= 12'b111011101100;
   8545: result <= 12'b111011101100;
   8546: result <= 12'b111011101011;
   8547: result <= 12'b111011101010;
   8548: result <= 12'b111011101001;
   8549: result <= 12'b111011101000;
   8550: result <= 12'b111011101000;
   8551: result <= 12'b111011100111;
   8552: result <= 12'b111011100110;
   8553: result <= 12'b111011100101;
   8554: result <= 12'b111011100101;
   8555: result <= 12'b111011100100;
   8556: result <= 12'b111011100011;
   8557: result <= 12'b111011100010;
   8558: result <= 12'b111011100001;
   8559: result <= 12'b111011100001;
   8560: result <= 12'b111011100000;
   8561: result <= 12'b111011011111;
   8562: result <= 12'b111011011110;
   8563: result <= 12'b111011011110;
   8564: result <= 12'b111011011101;
   8565: result <= 12'b111011011100;
   8566: result <= 12'b111011011011;
   8567: result <= 12'b111011011010;
   8568: result <= 12'b111011011010;
   8569: result <= 12'b111011011001;
   8570: result <= 12'b111011011000;
   8571: result <= 12'b111011010111;
   8572: result <= 12'b111011010111;
   8573: result <= 12'b111011010110;
   8574: result <= 12'b111011010101;
   8575: result <= 12'b111011010100;
   8576: result <= 12'b111011010011;
   8577: result <= 12'b111011010011;
   8578: result <= 12'b111011010010;
   8579: result <= 12'b111011010001;
   8580: result <= 12'b111011010000;
   8581: result <= 12'b111011010000;
   8582: result <= 12'b111011001111;
   8583: result <= 12'b111011001110;
   8584: result <= 12'b111011001101;
   8585: result <= 12'b111011001101;
   8586: result <= 12'b111011001100;
   8587: result <= 12'b111011001011;
   8588: result <= 12'b111011001010;
   8589: result <= 12'b111011001001;
   8590: result <= 12'b111011001001;
   8591: result <= 12'b111011001000;
   8592: result <= 12'b111011000111;
   8593: result <= 12'b111011000110;
   8594: result <= 12'b111011000110;
   8595: result <= 12'b111011000101;
   8596: result <= 12'b111011000100;
   8597: result <= 12'b111011000011;
   8598: result <= 12'b111011000010;
   8599: result <= 12'b111011000010;
   8600: result <= 12'b111011000001;
   8601: result <= 12'b111011000000;
   8602: result <= 12'b111010111111;
   8603: result <= 12'b111010111111;
   8604: result <= 12'b111010111110;
   8605: result <= 12'b111010111101;
   8606: result <= 12'b111010111100;
   8607: result <= 12'b111010111011;
   8608: result <= 12'b111010111011;
   8609: result <= 12'b111010111010;
   8610: result <= 12'b111010111001;
   8611: result <= 12'b111010111000;
   8612: result <= 12'b111010111000;
   8613: result <= 12'b111010110111;
   8614: result <= 12'b111010110110;
   8615: result <= 12'b111010110101;
   8616: result <= 12'b111010110100;
   8617: result <= 12'b111010110100;
   8618: result <= 12'b111010110011;
   8619: result <= 12'b111010110010;
   8620: result <= 12'b111010110001;
   8621: result <= 12'b111010110001;
   8622: result <= 12'b111010110000;
   8623: result <= 12'b111010101111;
   8624: result <= 12'b111010101110;
   8625: result <= 12'b111010101101;
   8626: result <= 12'b111010101101;
   8627: result <= 12'b111010101100;
   8628: result <= 12'b111010101011;
   8629: result <= 12'b111010101010;
   8630: result <= 12'b111010101010;
   8631: result <= 12'b111010101001;
   8632: result <= 12'b111010101000;
   8633: result <= 12'b111010100111;
   8634: result <= 12'b111010100111;
   8635: result <= 12'b111010100110;
   8636: result <= 12'b111010100101;
   8637: result <= 12'b111010100100;
   8638: result <= 12'b111010100011;
   8639: result <= 12'b111010100011;
   8640: result <= 12'b111010100010;
   8641: result <= 12'b111010100001;
   8642: result <= 12'b111010100000;
   8643: result <= 12'b111010100000;
   8644: result <= 12'b111010011111;
   8645: result <= 12'b111010011110;
   8646: result <= 12'b111010011101;
   8647: result <= 12'b111010011100;
   8648: result <= 12'b111010011100;
   8649: result <= 12'b111010011011;
   8650: result <= 12'b111010011010;
   8651: result <= 12'b111010011001;
   8652: result <= 12'b111010011001;
   8653: result <= 12'b111010011000;
   8654: result <= 12'b111010010111;
   8655: result <= 12'b111010010110;
   8656: result <= 12'b111010010101;
   8657: result <= 12'b111010010101;
   8658: result <= 12'b111010010100;
   8659: result <= 12'b111010010011;
   8660: result <= 12'b111010010010;
   8661: result <= 12'b111010010010;
   8662: result <= 12'b111010010001;
   8663: result <= 12'b111010010000;
   8664: result <= 12'b111010001111;
   8665: result <= 12'b111010001111;
   8666: result <= 12'b111010001110;
   8667: result <= 12'b111010001101;
   8668: result <= 12'b111010001100;
   8669: result <= 12'b111010001011;
   8670: result <= 12'b111010001011;
   8671: result <= 12'b111010001010;
   8672: result <= 12'b111010001001;
   8673: result <= 12'b111010001000;
   8674: result <= 12'b111010001000;
   8675: result <= 12'b111010000111;
   8676: result <= 12'b111010000110;
   8677: result <= 12'b111010000101;
   8678: result <= 12'b111010000101;
   8679: result <= 12'b111010000100;
   8680: result <= 12'b111010000011;
   8681: result <= 12'b111010000010;
   8682: result <= 12'b111010000001;
   8683: result <= 12'b111010000001;
   8684: result <= 12'b111010000000;
   8685: result <= 12'b111001111111;
   8686: result <= 12'b111001111110;
   8687: result <= 12'b111001111110;
   8688: result <= 12'b111001111101;
   8689: result <= 12'b111001111100;
   8690: result <= 12'b111001111011;
   8691: result <= 12'b111001111010;
   8692: result <= 12'b111001111010;
   8693: result <= 12'b111001111001;
   8694: result <= 12'b111001111000;
   8695: result <= 12'b111001110111;
   8696: result <= 12'b111001110111;
   8697: result <= 12'b111001110110;
   8698: result <= 12'b111001110101;
   8699: result <= 12'b111001110100;
   8700: result <= 12'b111001110100;
   8701: result <= 12'b111001110011;
   8702: result <= 12'b111001110010;
   8703: result <= 12'b111001110001;
   8704: result <= 12'b111001110000;
   8705: result <= 12'b111001110000;
   8706: result <= 12'b111001101111;
   8707: result <= 12'b111001101110;
   8708: result <= 12'b111001101101;
   8709: result <= 12'b111001101101;
   8710: result <= 12'b111001101100;
   8711: result <= 12'b111001101011;
   8712: result <= 12'b111001101010;
   8713: result <= 12'b111001101010;
   8714: result <= 12'b111001101001;
   8715: result <= 12'b111001101000;
   8716: result <= 12'b111001100111;
   8717: result <= 12'b111001100110;
   8718: result <= 12'b111001100110;
   8719: result <= 12'b111001100101;
   8720: result <= 12'b111001100100;
   8721: result <= 12'b111001100011;
   8722: result <= 12'b111001100011;
   8723: result <= 12'b111001100010;
   8724: result <= 12'b111001100001;
   8725: result <= 12'b111001100000;
   8726: result <= 12'b111001100000;
   8727: result <= 12'b111001011111;
   8728: result <= 12'b111001011110;
   8729: result <= 12'b111001011101;
   8730: result <= 12'b111001011100;
   8731: result <= 12'b111001011100;
   8732: result <= 12'b111001011011;
   8733: result <= 12'b111001011010;
   8734: result <= 12'b111001011001;
   8735: result <= 12'b111001011001;
   8736: result <= 12'b111001011000;
   8737: result <= 12'b111001010111;
   8738: result <= 12'b111001010110;
   8739: result <= 12'b111001010110;
   8740: result <= 12'b111001010101;
   8741: result <= 12'b111001010100;
   8742: result <= 12'b111001010011;
   8743: result <= 12'b111001010010;
   8744: result <= 12'b111001010010;
   8745: result <= 12'b111001010001;
   8746: result <= 12'b111001010000;
   8747: result <= 12'b111001001111;
   8748: result <= 12'b111001001111;
   8749: result <= 12'b111001001110;
   8750: result <= 12'b111001001101;
   8751: result <= 12'b111001001100;
   8752: result <= 12'b111001001100;
   8753: result <= 12'b111001001011;
   8754: result <= 12'b111001001010;
   8755: result <= 12'b111001001001;
   8756: result <= 12'b111001001000;
   8757: result <= 12'b111001001000;
   8758: result <= 12'b111001000111;
   8759: result <= 12'b111001000110;
   8760: result <= 12'b111001000101;
   8761: result <= 12'b111001000101;
   8762: result <= 12'b111001000100;
   8763: result <= 12'b111001000011;
   8764: result <= 12'b111001000010;
   8765: result <= 12'b111001000010;
   8766: result <= 12'b111001000001;
   8767: result <= 12'b111001000000;
   8768: result <= 12'b111000111111;
   8769: result <= 12'b111000111111;
   8770: result <= 12'b111000111110;
   8771: result <= 12'b111000111101;
   8772: result <= 12'b111000111100;
   8773: result <= 12'b111000111011;
   8774: result <= 12'b111000111011;
   8775: result <= 12'b111000111010;
   8776: result <= 12'b111000111001;
   8777: result <= 12'b111000111000;
   8778: result <= 12'b111000111000;
   8779: result <= 12'b111000110111;
   8780: result <= 12'b111000110110;
   8781: result <= 12'b111000110101;
   8782: result <= 12'b111000110101;
   8783: result <= 12'b111000110100;
   8784: result <= 12'b111000110011;
   8785: result <= 12'b111000110010;
   8786: result <= 12'b111000110001;
   8787: result <= 12'b111000110001;
   8788: result <= 12'b111000110000;
   8789: result <= 12'b111000101111;
   8790: result <= 12'b111000101110;
   8791: result <= 12'b111000101110;
   8792: result <= 12'b111000101101;
   8793: result <= 12'b111000101100;
   8794: result <= 12'b111000101011;
   8795: result <= 12'b111000101011;
   8796: result <= 12'b111000101010;
   8797: result <= 12'b111000101001;
   8798: result <= 12'b111000101000;
   8799: result <= 12'b111000101000;
   8800: result <= 12'b111000100111;
   8801: result <= 12'b111000100110;
   8802: result <= 12'b111000100101;
   8803: result <= 12'b111000100101;
   8804: result <= 12'b111000100100;
   8805: result <= 12'b111000100011;
   8806: result <= 12'b111000100010;
   8807: result <= 12'b111000100001;
   8808: result <= 12'b111000100001;
   8809: result <= 12'b111000100000;
   8810: result <= 12'b111000011111;
   8811: result <= 12'b111000011110;
   8812: result <= 12'b111000011110;
   8813: result <= 12'b111000011101;
   8814: result <= 12'b111000011100;
   8815: result <= 12'b111000011011;
   8816: result <= 12'b111000011011;
   8817: result <= 12'b111000011010;
   8818: result <= 12'b111000011001;
   8819: result <= 12'b111000011000;
   8820: result <= 12'b111000011000;
   8821: result <= 12'b111000010111;
   8822: result <= 12'b111000010110;
   8823: result <= 12'b111000010101;
   8824: result <= 12'b111000010100;
   8825: result <= 12'b111000010100;
   8826: result <= 12'b111000010011;
   8827: result <= 12'b111000010010;
   8828: result <= 12'b111000010001;
   8829: result <= 12'b111000010001;
   8830: result <= 12'b111000010000;
   8831: result <= 12'b111000001111;
   8832: result <= 12'b111000001110;
   8833: result <= 12'b111000001110;
   8834: result <= 12'b111000001101;
   8835: result <= 12'b111000001100;
   8836: result <= 12'b111000001011;
   8837: result <= 12'b111000001011;
   8838: result <= 12'b111000001010;
   8839: result <= 12'b111000001001;
   8840: result <= 12'b111000001000;
   8841: result <= 12'b111000001000;
   8842: result <= 12'b111000000111;
   8843: result <= 12'b111000000110;
   8844: result <= 12'b111000000101;
   8845: result <= 12'b111000000100;
   8846: result <= 12'b111000000100;
   8847: result <= 12'b111000000011;
   8848: result <= 12'b111000000010;
   8849: result <= 12'b111000000001;
   8850: result <= 12'b111000000001;
   8851: result <= 12'b111000000000;
   8852: result <= 12'b110111111111;
   8853: result <= 12'b110111111110;
   8854: result <= 12'b110111111110;
   8855: result <= 12'b110111111101;
   8856: result <= 12'b110111111100;
   8857: result <= 12'b110111111011;
   8858: result <= 12'b110111111011;
   8859: result <= 12'b110111111010;
   8860: result <= 12'b110111111001;
   8861: result <= 12'b110111111000;
   8862: result <= 12'b110111111000;
   8863: result <= 12'b110111110111;
   8864: result <= 12'b110111110110;
   8865: result <= 12'b110111110101;
   8866: result <= 12'b110111110101;
   8867: result <= 12'b110111110100;
   8868: result <= 12'b110111110011;
   8869: result <= 12'b110111110010;
   8870: result <= 12'b110111110001;
   8871: result <= 12'b110111110001;
   8872: result <= 12'b110111110000;
   8873: result <= 12'b110111101111;
   8874: result <= 12'b110111101110;
   8875: result <= 12'b110111101110;
   8876: result <= 12'b110111101101;
   8877: result <= 12'b110111101100;
   8878: result <= 12'b110111101011;
   8879: result <= 12'b110111101011;
   8880: result <= 12'b110111101010;
   8881: result <= 12'b110111101001;
   8882: result <= 12'b110111101000;
   8883: result <= 12'b110111101000;
   8884: result <= 12'b110111100111;
   8885: result <= 12'b110111100110;
   8886: result <= 12'b110111100101;
   8887: result <= 12'b110111100101;
   8888: result <= 12'b110111100100;
   8889: result <= 12'b110111100011;
   8890: result <= 12'b110111100010;
   8891: result <= 12'b110111100010;
   8892: result <= 12'b110111100001;
   8893: result <= 12'b110111100000;
   8894: result <= 12'b110111011111;
   8895: result <= 12'b110111011111;
   8896: result <= 12'b110111011110;
   8897: result <= 12'b110111011101;
   8898: result <= 12'b110111011100;
   8899: result <= 12'b110111011100;
   8900: result <= 12'b110111011011;
   8901: result <= 12'b110111011010;
   8902: result <= 12'b110111011001;
   8903: result <= 12'b110111011000;
   8904: result <= 12'b110111011000;
   8905: result <= 12'b110111010111;
   8906: result <= 12'b110111010110;
   8907: result <= 12'b110111010101;
   8908: result <= 12'b110111010101;
   8909: result <= 12'b110111010100;
   8910: result <= 12'b110111010011;
   8911: result <= 12'b110111010010;
   8912: result <= 12'b110111010010;
   8913: result <= 12'b110111010001;
   8914: result <= 12'b110111010000;
   8915: result <= 12'b110111001111;
   8916: result <= 12'b110111001111;
   8917: result <= 12'b110111001110;
   8918: result <= 12'b110111001101;
   8919: result <= 12'b110111001100;
   8920: result <= 12'b110111001100;
   8921: result <= 12'b110111001011;
   8922: result <= 12'b110111001010;
   8923: result <= 12'b110111001001;
   8924: result <= 12'b110111001001;
   8925: result <= 12'b110111001000;
   8926: result <= 12'b110111000111;
   8927: result <= 12'b110111000110;
   8928: result <= 12'b110111000110;
   8929: result <= 12'b110111000101;
   8930: result <= 12'b110111000100;
   8931: result <= 12'b110111000011;
   8932: result <= 12'b110111000011;
   8933: result <= 12'b110111000010;
   8934: result <= 12'b110111000001;
   8935: result <= 12'b110111000000;
   8936: result <= 12'b110111000000;
   8937: result <= 12'b110110111111;
   8938: result <= 12'b110110111110;
   8939: result <= 12'b110110111101;
   8940: result <= 12'b110110111101;
   8941: result <= 12'b110110111100;
   8942: result <= 12'b110110111011;
   8943: result <= 12'b110110111010;
   8944: result <= 12'b110110111010;
   8945: result <= 12'b110110111001;
   8946: result <= 12'b110110111000;
   8947: result <= 12'b110110110111;
   8948: result <= 12'b110110110111;
   8949: result <= 12'b110110110110;
   8950: result <= 12'b110110110101;
   8951: result <= 12'b110110110100;
   8952: result <= 12'b110110110100;
   8953: result <= 12'b110110110011;
   8954: result <= 12'b110110110010;
   8955: result <= 12'b110110110001;
   8956: result <= 12'b110110110001;
   8957: result <= 12'b110110110000;
   8958: result <= 12'b110110101111;
   8959: result <= 12'b110110101110;
   8960: result <= 12'b110110101101;
   8961: result <= 12'b110110101101;
   8962: result <= 12'b110110101100;
   8963: result <= 12'b110110101011;
   8964: result <= 12'b110110101010;
   8965: result <= 12'b110110101010;
   8966: result <= 12'b110110101001;
   8967: result <= 12'b110110101000;
   8968: result <= 12'b110110100111;
   8969: result <= 12'b110110100111;
   8970: result <= 12'b110110100110;
   8971: result <= 12'b110110100101;
   8972: result <= 12'b110110100100;
   8973: result <= 12'b110110100100;
   8974: result <= 12'b110110100011;
   8975: result <= 12'b110110100010;
   8976: result <= 12'b110110100001;
   8977: result <= 12'b110110100001;
   8978: result <= 12'b110110100000;
   8979: result <= 12'b110110011111;
   8980: result <= 12'b110110011110;
   8981: result <= 12'b110110011110;
   8982: result <= 12'b110110011101;
   8983: result <= 12'b110110011100;
   8984: result <= 12'b110110011011;
   8985: result <= 12'b110110011011;
   8986: result <= 12'b110110011010;
   8987: result <= 12'b110110011001;
   8988: result <= 12'b110110011000;
   8989: result <= 12'b110110011000;
   8990: result <= 12'b110110010111;
   8991: result <= 12'b110110010110;
   8992: result <= 12'b110110010101;
   8993: result <= 12'b110110010101;
   8994: result <= 12'b110110010100;
   8995: result <= 12'b110110010011;
   8996: result <= 12'b110110010010;
   8997: result <= 12'b110110010010;
   8998: result <= 12'b110110010001;
   8999: result <= 12'b110110010000;
   9000: result <= 12'b110110010000;
   9001: result <= 12'b110110001111;
   9002: result <= 12'b110110001110;
   9003: result <= 12'b110110001101;
   9004: result <= 12'b110110001101;
   9005: result <= 12'b110110001100;
   9006: result <= 12'b110110001011;
   9007: result <= 12'b110110001010;
   9008: result <= 12'b110110001010;
   9009: result <= 12'b110110001001;
   9010: result <= 12'b110110001000;
   9011: result <= 12'b110110000111;
   9012: result <= 12'b110110000111;
   9013: result <= 12'b110110000110;
   9014: result <= 12'b110110000101;
   9015: result <= 12'b110110000100;
   9016: result <= 12'b110110000100;
   9017: result <= 12'b110110000011;
   9018: result <= 12'b110110000010;
   9019: result <= 12'b110110000001;
   9020: result <= 12'b110110000001;
   9021: result <= 12'b110110000000;
   9022: result <= 12'b110101111111;
   9023: result <= 12'b110101111110;
   9024: result <= 12'b110101111110;
   9025: result <= 12'b110101111101;
   9026: result <= 12'b110101111100;
   9027: result <= 12'b110101111011;
   9028: result <= 12'b110101111011;
   9029: result <= 12'b110101111010;
   9030: result <= 12'b110101111001;
   9031: result <= 12'b110101111000;
   9032: result <= 12'b110101111000;
   9033: result <= 12'b110101110111;
   9034: result <= 12'b110101110110;
   9035: result <= 12'b110101110101;
   9036: result <= 12'b110101110101;
   9037: result <= 12'b110101110100;
   9038: result <= 12'b110101110011;
   9039: result <= 12'b110101110010;
   9040: result <= 12'b110101110010;
   9041: result <= 12'b110101110001;
   9042: result <= 12'b110101110000;
   9043: result <= 12'b110101101111;
   9044: result <= 12'b110101101111;
   9045: result <= 12'b110101101110;
   9046: result <= 12'b110101101101;
   9047: result <= 12'b110101101100;
   9048: result <= 12'b110101101100;
   9049: result <= 12'b110101101011;
   9050: result <= 12'b110101101010;
   9051: result <= 12'b110101101001;
   9052: result <= 12'b110101101001;
   9053: result <= 12'b110101101000;
   9054: result <= 12'b110101100111;
   9055: result <= 12'b110101100111;
   9056: result <= 12'b110101100110;
   9057: result <= 12'b110101100101;
   9058: result <= 12'b110101100100;
   9059: result <= 12'b110101100100;
   9060: result <= 12'b110101100011;
   9061: result <= 12'b110101100010;
   9062: result <= 12'b110101100001;
   9063: result <= 12'b110101100001;
   9064: result <= 12'b110101100000;
   9065: result <= 12'b110101011111;
   9066: result <= 12'b110101011110;
   9067: result <= 12'b110101011110;
   9068: result <= 12'b110101011101;
   9069: result <= 12'b110101011100;
   9070: result <= 12'b110101011011;
   9071: result <= 12'b110101011011;
   9072: result <= 12'b110101011010;
   9073: result <= 12'b110101011001;
   9074: result <= 12'b110101011000;
   9075: result <= 12'b110101011000;
   9076: result <= 12'b110101010111;
   9077: result <= 12'b110101010110;
   9078: result <= 12'b110101010101;
   9079: result <= 12'b110101010101;
   9080: result <= 12'b110101010100;
   9081: result <= 12'b110101010011;
   9082: result <= 12'b110101010010;
   9083: result <= 12'b110101010010;
   9084: result <= 12'b110101010001;
   9085: result <= 12'b110101010000;
   9086: result <= 12'b110101010000;
   9087: result <= 12'b110101001111;
   9088: result <= 12'b110101001110;
   9089: result <= 12'b110101001101;
   9090: result <= 12'b110101001101;
   9091: result <= 12'b110101001100;
   9092: result <= 12'b110101001011;
   9093: result <= 12'b110101001010;
   9094: result <= 12'b110101001010;
   9095: result <= 12'b110101001001;
   9096: result <= 12'b110101001000;
   9097: result <= 12'b110101000111;
   9098: result <= 12'b110101000111;
   9099: result <= 12'b110101000110;
   9100: result <= 12'b110101000101;
   9101: result <= 12'b110101000100;
   9102: result <= 12'b110101000100;
   9103: result <= 12'b110101000011;
   9104: result <= 12'b110101000010;
   9105: result <= 12'b110101000001;
   9106: result <= 12'b110101000001;
   9107: result <= 12'b110101000000;
   9108: result <= 12'b110100111111;
   9109: result <= 12'b110100111111;
   9110: result <= 12'b110100111110;
   9111: result <= 12'b110100111101;
   9112: result <= 12'b110100111100;
   9113: result <= 12'b110100111100;
   9114: result <= 12'b110100111011;
   9115: result <= 12'b110100111010;
   9116: result <= 12'b110100111001;
   9117: result <= 12'b110100111001;
   9118: result <= 12'b110100111000;
   9119: result <= 12'b110100110111;
   9120: result <= 12'b110100110110;
   9121: result <= 12'b110100110110;
   9122: result <= 12'b110100110101;
   9123: result <= 12'b110100110100;
   9124: result <= 12'b110100110011;
   9125: result <= 12'b110100110011;
   9126: result <= 12'b110100110010;
   9127: result <= 12'b110100110001;
   9128: result <= 12'b110100110001;
   9129: result <= 12'b110100110000;
   9130: result <= 12'b110100101111;
   9131: result <= 12'b110100101110;
   9132: result <= 12'b110100101110;
   9133: result <= 12'b110100101101;
   9134: result <= 12'b110100101100;
   9135: result <= 12'b110100101011;
   9136: result <= 12'b110100101011;
   9137: result <= 12'b110100101010;
   9138: result <= 12'b110100101001;
   9139: result <= 12'b110100101000;
   9140: result <= 12'b110100101000;
   9141: result <= 12'b110100100111;
   9142: result <= 12'b110100100110;
   9143: result <= 12'b110100100110;
   9144: result <= 12'b110100100101;
   9145: result <= 12'b110100100100;
   9146: result <= 12'b110100100011;
   9147: result <= 12'b110100100011;
   9148: result <= 12'b110100100010;
   9149: result <= 12'b110100100001;
   9150: result <= 12'b110100100000;
   9151: result <= 12'b110100100000;
   9152: result <= 12'b110100011111;
   9153: result <= 12'b110100011110;
   9154: result <= 12'b110100011101;
   9155: result <= 12'b110100011101;
   9156: result <= 12'b110100011100;
   9157: result <= 12'b110100011011;
   9158: result <= 12'b110100011011;
   9159: result <= 12'b110100011010;
   9160: result <= 12'b110100011001;
   9161: result <= 12'b110100011000;
   9162: result <= 12'b110100011000;
   9163: result <= 12'b110100010111;
   9164: result <= 12'b110100010110;
   9165: result <= 12'b110100010101;
   9166: result <= 12'b110100010101;
   9167: result <= 12'b110100010100;
   9168: result <= 12'b110100010011;
   9169: result <= 12'b110100010010;
   9170: result <= 12'b110100010010;
   9171: result <= 12'b110100010001;
   9172: result <= 12'b110100010000;
   9173: result <= 12'b110100010000;
   9174: result <= 12'b110100001111;
   9175: result <= 12'b110100001110;
   9176: result <= 12'b110100001101;
   9177: result <= 12'b110100001101;
   9178: result <= 12'b110100001100;
   9179: result <= 12'b110100001011;
   9180: result <= 12'b110100001010;
   9181: result <= 12'b110100001010;
   9182: result <= 12'b110100001001;
   9183: result <= 12'b110100001000;
   9184: result <= 12'b110100001000;
   9185: result <= 12'b110100000111;
   9186: result <= 12'b110100000110;
   9187: result <= 12'b110100000101;
   9188: result <= 12'b110100000101;
   9189: result <= 12'b110100000100;
   9190: result <= 12'b110100000011;
   9191: result <= 12'b110100000010;
   9192: result <= 12'b110100000010;
   9193: result <= 12'b110100000001;
   9194: result <= 12'b110100000000;
   9195: result <= 12'b110100000000;
   9196: result <= 12'b110011111111;
   9197: result <= 12'b110011111110;
   9198: result <= 12'b110011111101;
   9199: result <= 12'b110011111101;
   9200: result <= 12'b110011111100;
   9201: result <= 12'b110011111011;
   9202: result <= 12'b110011111010;
   9203: result <= 12'b110011111010;
   9204: result <= 12'b110011111001;
   9205: result <= 12'b110011111000;
   9206: result <= 12'b110011111000;
   9207: result <= 12'b110011110111;
   9208: result <= 12'b110011110110;
   9209: result <= 12'b110011110101;
   9210: result <= 12'b110011110101;
   9211: result <= 12'b110011110100;
   9212: result <= 12'b110011110011;
   9213: result <= 12'b110011110010;
   9214: result <= 12'b110011110010;
   9215: result <= 12'b110011110001;
   9216: result <= 12'b110011110000;
   9217: result <= 12'b110011110000;
   9218: result <= 12'b110011101111;
   9219: result <= 12'b110011101110;
   9220: result <= 12'b110011101101;
   9221: result <= 12'b110011101101;
   9222: result <= 12'b110011101100;
   9223: result <= 12'b110011101011;
   9224: result <= 12'b110011101010;
   9225: result <= 12'b110011101010;
   9226: result <= 12'b110011101001;
   9227: result <= 12'b110011101000;
   9228: result <= 12'b110011101000;
   9229: result <= 12'b110011100111;
   9230: result <= 12'b110011100110;
   9231: result <= 12'b110011100101;
   9232: result <= 12'b110011100101;
   9233: result <= 12'b110011100100;
   9234: result <= 12'b110011100011;
   9235: result <= 12'b110011100010;
   9236: result <= 12'b110011100010;
   9237: result <= 12'b110011100001;
   9238: result <= 12'b110011100000;
   9239: result <= 12'b110011100000;
   9240: result <= 12'b110011011111;
   9241: result <= 12'b110011011110;
   9242: result <= 12'b110011011101;
   9243: result <= 12'b110011011101;
   9244: result <= 12'b110011011100;
   9245: result <= 12'b110011011011;
   9246: result <= 12'b110011011011;
   9247: result <= 12'b110011011010;
   9248: result <= 12'b110011011001;
   9249: result <= 12'b110011011000;
   9250: result <= 12'b110011011000;
   9251: result <= 12'b110011010111;
   9252: result <= 12'b110011010110;
   9253: result <= 12'b110011010101;
   9254: result <= 12'b110011010101;
   9255: result <= 12'b110011010100;
   9256: result <= 12'b110011010011;
   9257: result <= 12'b110011010011;
   9258: result <= 12'b110011010010;
   9259: result <= 12'b110011010001;
   9260: result <= 12'b110011010000;
   9261: result <= 12'b110011010000;
   9262: result <= 12'b110011001111;
   9263: result <= 12'b110011001110;
   9264: result <= 12'b110011001110;
   9265: result <= 12'b110011001101;
   9266: result <= 12'b110011001100;
   9267: result <= 12'b110011001011;
   9268: result <= 12'b110011001011;
   9269: result <= 12'b110011001010;
   9270: result <= 12'b110011001001;
   9271: result <= 12'b110011001001;
   9272: result <= 12'b110011001000;
   9273: result <= 12'b110011000111;
   9274: result <= 12'b110011000110;
   9275: result <= 12'b110011000110;
   9276: result <= 12'b110011000101;
   9277: result <= 12'b110011000100;
   9278: result <= 12'b110011000100;
   9279: result <= 12'b110011000011;
   9280: result <= 12'b110011000010;
   9281: result <= 12'b110011000001;
   9282: result <= 12'b110011000001;
   9283: result <= 12'b110011000000;
   9284: result <= 12'b110010111111;
   9285: result <= 12'b110010111110;
   9286: result <= 12'b110010111110;
   9287: result <= 12'b110010111101;
   9288: result <= 12'b110010111100;
   9289: result <= 12'b110010111100;
   9290: result <= 12'b110010111011;
   9291: result <= 12'b110010111010;
   9292: result <= 12'b110010111001;
   9293: result <= 12'b110010111001;
   9294: result <= 12'b110010111000;
   9295: result <= 12'b110010110111;
   9296: result <= 12'b110010110111;
   9297: result <= 12'b110010110110;
   9298: result <= 12'b110010110101;
   9299: result <= 12'b110010110100;
   9300: result <= 12'b110010110100;
   9301: result <= 12'b110010110011;
   9302: result <= 12'b110010110010;
   9303: result <= 12'b110010110010;
   9304: result <= 12'b110010110001;
   9305: result <= 12'b110010110000;
   9306: result <= 12'b110010101111;
   9307: result <= 12'b110010101111;
   9308: result <= 12'b110010101110;
   9309: result <= 12'b110010101101;
   9310: result <= 12'b110010101101;
   9311: result <= 12'b110010101100;
   9312: result <= 12'b110010101011;
   9313: result <= 12'b110010101010;
   9314: result <= 12'b110010101010;
   9315: result <= 12'b110010101001;
   9316: result <= 12'b110010101000;
   9317: result <= 12'b110010101000;
   9318: result <= 12'b110010100111;
   9319: result <= 12'b110010100110;
   9320: result <= 12'b110010100101;
   9321: result <= 12'b110010100101;
   9322: result <= 12'b110010100100;
   9323: result <= 12'b110010100011;
   9324: result <= 12'b110010100011;
   9325: result <= 12'b110010100010;
   9326: result <= 12'b110010100001;
   9327: result <= 12'b110010100000;
   9328: result <= 12'b110010100000;
   9329: result <= 12'b110010011111;
   9330: result <= 12'b110010011110;
   9331: result <= 12'b110010011110;
   9332: result <= 12'b110010011101;
   9333: result <= 12'b110010011100;
   9334: result <= 12'b110010011011;
   9335: result <= 12'b110010011011;
   9336: result <= 12'b110010011010;
   9337: result <= 12'b110010011001;
   9338: result <= 12'b110010011001;
   9339: result <= 12'b110010011000;
   9340: result <= 12'b110010010111;
   9341: result <= 12'b110010010110;
   9342: result <= 12'b110010010110;
   9343: result <= 12'b110010010101;
   9344: result <= 12'b110010010100;
   9345: result <= 12'b110010010100;
   9346: result <= 12'b110010010011;
   9347: result <= 12'b110010010010;
   9348: result <= 12'b110010010010;
   9349: result <= 12'b110010010001;
   9350: result <= 12'b110010010000;
   9351: result <= 12'b110010001111;
   9352: result <= 12'b110010001111;
   9353: result <= 12'b110010001110;
   9354: result <= 12'b110010001101;
   9355: result <= 12'b110010001101;
   9356: result <= 12'b110010001100;
   9357: result <= 12'b110010001011;
   9358: result <= 12'b110010001010;
   9359: result <= 12'b110010001010;
   9360: result <= 12'b110010001001;
   9361: result <= 12'b110010001000;
   9362: result <= 12'b110010001000;
   9363: result <= 12'b110010000111;
   9364: result <= 12'b110010000110;
   9365: result <= 12'b110010000101;
   9366: result <= 12'b110010000101;
   9367: result <= 12'b110010000100;
   9368: result <= 12'b110010000011;
   9369: result <= 12'b110010000011;
   9370: result <= 12'b110010000010;
   9371: result <= 12'b110010000001;
   9372: result <= 12'b110010000001;
   9373: result <= 12'b110010000000;
   9374: result <= 12'b110001111111;
   9375: result <= 12'b110001111110;
   9376: result <= 12'b110001111110;
   9377: result <= 12'b110001111101;
   9378: result <= 12'b110001111100;
   9379: result <= 12'b110001111100;
   9380: result <= 12'b110001111011;
   9381: result <= 12'b110001111010;
   9382: result <= 12'b110001111001;
   9383: result <= 12'b110001111001;
   9384: result <= 12'b110001111000;
   9385: result <= 12'b110001110111;
   9386: result <= 12'b110001110111;
   9387: result <= 12'b110001110110;
   9388: result <= 12'b110001110101;
   9389: result <= 12'b110001110101;
   9390: result <= 12'b110001110100;
   9391: result <= 12'b110001110011;
   9392: result <= 12'b110001110010;
   9393: result <= 12'b110001110010;
   9394: result <= 12'b110001110001;
   9395: result <= 12'b110001110000;
   9396: result <= 12'b110001110000;
   9397: result <= 12'b110001101111;
   9398: result <= 12'b110001101110;
   9399: result <= 12'b110001101110;
   9400: result <= 12'b110001101101;
   9401: result <= 12'b110001101100;
   9402: result <= 12'b110001101011;
   9403: result <= 12'b110001101011;
   9404: result <= 12'b110001101010;
   9405: result <= 12'b110001101001;
   9406: result <= 12'b110001101001;
   9407: result <= 12'b110001101000;
   9408: result <= 12'b110001100111;
   9409: result <= 12'b110001100110;
   9410: result <= 12'b110001100110;
   9411: result <= 12'b110001100101;
   9412: result <= 12'b110001100100;
   9413: result <= 12'b110001100100;
   9414: result <= 12'b110001100011;
   9415: result <= 12'b110001100010;
   9416: result <= 12'b110001100010;
   9417: result <= 12'b110001100001;
   9418: result <= 12'b110001100000;
   9419: result <= 12'b110001011111;
   9420: result <= 12'b110001011111;
   9421: result <= 12'b110001011110;
   9422: result <= 12'b110001011101;
   9423: result <= 12'b110001011101;
   9424: result <= 12'b110001011100;
   9425: result <= 12'b110001011011;
   9426: result <= 12'b110001011011;
   9427: result <= 12'b110001011010;
   9428: result <= 12'b110001011001;
   9429: result <= 12'b110001011000;
   9430: result <= 12'b110001011000;
   9431: result <= 12'b110001010111;
   9432: result <= 12'b110001010110;
   9433: result <= 12'b110001010110;
   9434: result <= 12'b110001010101;
   9435: result <= 12'b110001010100;
   9436: result <= 12'b110001010100;
   9437: result <= 12'b110001010011;
   9438: result <= 12'b110001010010;
   9439: result <= 12'b110001010010;
   9440: result <= 12'b110001010001;
   9441: result <= 12'b110001010000;
   9442: result <= 12'b110001001111;
   9443: result <= 12'b110001001111;
   9444: result <= 12'b110001001110;
   9445: result <= 12'b110001001101;
   9446: result <= 12'b110001001101;
   9447: result <= 12'b110001001100;
   9448: result <= 12'b110001001011;
   9449: result <= 12'b110001001011;
   9450: result <= 12'b110001001010;
   9451: result <= 12'b110001001001;
   9452: result <= 12'b110001001000;
   9453: result <= 12'b110001001000;
   9454: result <= 12'b110001000111;
   9455: result <= 12'b110001000110;
   9456: result <= 12'b110001000110;
   9457: result <= 12'b110001000101;
   9458: result <= 12'b110001000100;
   9459: result <= 12'b110001000100;
   9460: result <= 12'b110001000011;
   9461: result <= 12'b110001000010;
   9462: result <= 12'b110001000010;
   9463: result <= 12'b110001000001;
   9464: result <= 12'b110001000000;
   9465: result <= 12'b110000111111;
   9466: result <= 12'b110000111111;
   9467: result <= 12'b110000111110;
   9468: result <= 12'b110000111101;
   9469: result <= 12'b110000111101;
   9470: result <= 12'b110000111100;
   9471: result <= 12'b110000111011;
   9472: result <= 12'b110000111011;
   9473: result <= 12'b110000111010;
   9474: result <= 12'b110000111001;
   9475: result <= 12'b110000111001;
   9476: result <= 12'b110000111000;
   9477: result <= 12'b110000110111;
   9478: result <= 12'b110000110110;
   9479: result <= 12'b110000110110;
   9480: result <= 12'b110000110101;
   9481: result <= 12'b110000110100;
   9482: result <= 12'b110000110100;
   9483: result <= 12'b110000110011;
   9484: result <= 12'b110000110010;
   9485: result <= 12'b110000110010;
   9486: result <= 12'b110000110001;
   9487: result <= 12'b110000110000;
   9488: result <= 12'b110000110000;
   9489: result <= 12'b110000101111;
   9490: result <= 12'b110000101110;
   9491: result <= 12'b110000101101;
   9492: result <= 12'b110000101101;
   9493: result <= 12'b110000101100;
   9494: result <= 12'b110000101011;
   9495: result <= 12'b110000101011;
   9496: result <= 12'b110000101010;
   9497: result <= 12'b110000101001;
   9498: result <= 12'b110000101001;
   9499: result <= 12'b110000101000;
   9500: result <= 12'b110000100111;
   9501: result <= 12'b110000100111;
   9502: result <= 12'b110000100110;
   9503: result <= 12'b110000100101;
   9504: result <= 12'b110000100100;
   9505: result <= 12'b110000100100;
   9506: result <= 12'b110000100011;
   9507: result <= 12'b110000100010;
   9508: result <= 12'b110000100010;
   9509: result <= 12'b110000100001;
   9510: result <= 12'b110000100000;
   9511: result <= 12'b110000100000;
   9512: result <= 12'b110000011111;
   9513: result <= 12'b110000011110;
   9514: result <= 12'b110000011110;
   9515: result <= 12'b110000011101;
   9516: result <= 12'b110000011100;
   9517: result <= 12'b110000011100;
   9518: result <= 12'b110000011011;
   9519: result <= 12'b110000011010;
   9520: result <= 12'b110000011001;
   9521: result <= 12'b110000011001;
   9522: result <= 12'b110000011000;
   9523: result <= 12'b110000010111;
   9524: result <= 12'b110000010111;
   9525: result <= 12'b110000010110;
   9526: result <= 12'b110000010101;
   9527: result <= 12'b110000010101;
   9528: result <= 12'b110000010100;
   9529: result <= 12'b110000010011;
   9530: result <= 12'b110000010011;
   9531: result <= 12'b110000010010;
   9532: result <= 12'b110000010001;
   9533: result <= 12'b110000010001;
   9534: result <= 12'b110000010000;
   9535: result <= 12'b110000001111;
   9536: result <= 12'b110000001111;
   9537: result <= 12'b110000001110;
   9538: result <= 12'b110000001101;
   9539: result <= 12'b110000001100;
   9540: result <= 12'b110000001100;
   9541: result <= 12'b110000001011;
   9542: result <= 12'b110000001010;
   9543: result <= 12'b110000001010;
   9544: result <= 12'b110000001001;
   9545: result <= 12'b110000001000;
   9546: result <= 12'b110000001000;
   9547: result <= 12'b110000000111;
   9548: result <= 12'b110000000110;
   9549: result <= 12'b110000000110;
   9550: result <= 12'b110000000101;
   9551: result <= 12'b110000000100;
   9552: result <= 12'b110000000100;
   9553: result <= 12'b110000000011;
   9554: result <= 12'b110000000010;
   9555: result <= 12'b110000000010;
   9556: result <= 12'b110000000001;
   9557: result <= 12'b110000000000;
   9558: result <= 12'b110000000000;
   9559: result <= 12'b101111111111;
   9560: result <= 12'b101111111110;
   9561: result <= 12'b101111111110;
   9562: result <= 12'b101111111101;
   9563: result <= 12'b101111111100;
   9564: result <= 12'b101111111011;
   9565: result <= 12'b101111111011;
   9566: result <= 12'b101111111010;
   9567: result <= 12'b101111111001;
   9568: result <= 12'b101111111001;
   9569: result <= 12'b101111111000;
   9570: result <= 12'b101111110111;
   9571: result <= 12'b101111110111;
   9572: result <= 12'b101111110110;
   9573: result <= 12'b101111110101;
   9574: result <= 12'b101111110101;
   9575: result <= 12'b101111110100;
   9576: result <= 12'b101111110011;
   9577: result <= 12'b101111110011;
   9578: result <= 12'b101111110010;
   9579: result <= 12'b101111110001;
   9580: result <= 12'b101111110001;
   9581: result <= 12'b101111110000;
   9582: result <= 12'b101111101111;
   9583: result <= 12'b101111101111;
   9584: result <= 12'b101111101110;
   9585: result <= 12'b101111101101;
   9586: result <= 12'b101111101101;
   9587: result <= 12'b101111101100;
   9588: result <= 12'b101111101011;
   9589: result <= 12'b101111101011;
   9590: result <= 12'b101111101010;
   9591: result <= 12'b101111101001;
   9592: result <= 12'b101111101001;
   9593: result <= 12'b101111101000;
   9594: result <= 12'b101111100111;
   9595: result <= 12'b101111100110;
   9596: result <= 12'b101111100110;
   9597: result <= 12'b101111100101;
   9598: result <= 12'b101111100100;
   9599: result <= 12'b101111100100;
   9600: result <= 12'b101111100011;
   9601: result <= 12'b101111100010;
   9602: result <= 12'b101111100010;
   9603: result <= 12'b101111100001;
   9604: result <= 12'b101111100000;
   9605: result <= 12'b101111100000;
   9606: result <= 12'b101111011111;
   9607: result <= 12'b101111011110;
   9608: result <= 12'b101111011110;
   9609: result <= 12'b101111011101;
   9610: result <= 12'b101111011100;
   9611: result <= 12'b101111011100;
   9612: result <= 12'b101111011011;
   9613: result <= 12'b101111011010;
   9614: result <= 12'b101111011010;
   9615: result <= 12'b101111011001;
   9616: result <= 12'b101111011000;
   9617: result <= 12'b101111011000;
   9618: result <= 12'b101111010111;
   9619: result <= 12'b101111010110;
   9620: result <= 12'b101111010110;
   9621: result <= 12'b101111010101;
   9622: result <= 12'b101111010100;
   9623: result <= 12'b101111010100;
   9624: result <= 12'b101111010011;
   9625: result <= 12'b101111010010;
   9626: result <= 12'b101111010010;
   9627: result <= 12'b101111010001;
   9628: result <= 12'b101111010000;
   9629: result <= 12'b101111010000;
   9630: result <= 12'b101111001111;
   9631: result <= 12'b101111001110;
   9632: result <= 12'b101111001110;
   9633: result <= 12'b101111001101;
   9634: result <= 12'b101111001100;
   9635: result <= 12'b101111001100;
   9636: result <= 12'b101111001011;
   9637: result <= 12'b101111001010;
   9638: result <= 12'b101111001010;
   9639: result <= 12'b101111001001;
   9640: result <= 12'b101111001000;
   9641: result <= 12'b101111001000;
   9642: result <= 12'b101111000111;
   9643: result <= 12'b101111000110;
   9644: result <= 12'b101111000110;
   9645: result <= 12'b101111000101;
   9646: result <= 12'b101111000100;
   9647: result <= 12'b101111000100;
   9648: result <= 12'b101111000011;
   9649: result <= 12'b101111000010;
   9650: result <= 12'b101111000010;
   9651: result <= 12'b101111000001;
   9652: result <= 12'b101111000000;
   9653: result <= 12'b101111000000;
   9654: result <= 12'b101110111111;
   9655: result <= 12'b101110111110;
   9656: result <= 12'b101110111110;
   9657: result <= 12'b101110111101;
   9658: result <= 12'b101110111100;
   9659: result <= 12'b101110111100;
   9660: result <= 12'b101110111011;
   9661: result <= 12'b101110111010;
   9662: result <= 12'b101110111010;
   9663: result <= 12'b101110111001;
   9664: result <= 12'b101110111000;
   9665: result <= 12'b101110111000;
   9666: result <= 12'b101110110111;
   9667: result <= 12'b101110110110;
   9668: result <= 12'b101110110110;
   9669: result <= 12'b101110110101;
   9670: result <= 12'b101110110100;
   9671: result <= 12'b101110110100;
   9672: result <= 12'b101110110011;
   9673: result <= 12'b101110110010;
   9674: result <= 12'b101110110010;
   9675: result <= 12'b101110110001;
   9676: result <= 12'b101110110000;
   9677: result <= 12'b101110110000;
   9678: result <= 12'b101110101111;
   9679: result <= 12'b101110101110;
   9680: result <= 12'b101110101110;
   9681: result <= 12'b101110101101;
   9682: result <= 12'b101110101100;
   9683: result <= 12'b101110101100;
   9684: result <= 12'b101110101011;
   9685: result <= 12'b101110101010;
   9686: result <= 12'b101110101010;
   9687: result <= 12'b101110101001;
   9688: result <= 12'b101110101000;
   9689: result <= 12'b101110101000;
   9690: result <= 12'b101110100111;
   9691: result <= 12'b101110100110;
   9692: result <= 12'b101110100110;
   9693: result <= 12'b101110100101;
   9694: result <= 12'b101110100100;
   9695: result <= 12'b101110100100;
   9696: result <= 12'b101110100011;
   9697: result <= 12'b101110100011;
   9698: result <= 12'b101110100010;
   9699: result <= 12'b101110100001;
   9700: result <= 12'b101110100001;
   9701: result <= 12'b101110100000;
   9702: result <= 12'b101110011111;
   9703: result <= 12'b101110011111;
   9704: result <= 12'b101110011110;
   9705: result <= 12'b101110011101;
   9706: result <= 12'b101110011101;
   9707: result <= 12'b101110011100;
   9708: result <= 12'b101110011011;
   9709: result <= 12'b101110011011;
   9710: result <= 12'b101110011010;
   9711: result <= 12'b101110011001;
   9712: result <= 12'b101110011001;
   9713: result <= 12'b101110011000;
   9714: result <= 12'b101110010111;
   9715: result <= 12'b101110010111;
   9716: result <= 12'b101110010110;
   9717: result <= 12'b101110010101;
   9718: result <= 12'b101110010101;
   9719: result <= 12'b101110010100;
   9720: result <= 12'b101110010011;
   9721: result <= 12'b101110010011;
   9722: result <= 12'b101110010010;
   9723: result <= 12'b101110010001;
   9724: result <= 12'b101110010001;
   9725: result <= 12'b101110010000;
   9726: result <= 12'b101110001111;
   9727: result <= 12'b101110001111;
   9728: result <= 12'b101110001110;
   9729: result <= 12'b101110001110;
   9730: result <= 12'b101110001101;
   9731: result <= 12'b101110001100;
   9732: result <= 12'b101110001100;
   9733: result <= 12'b101110001011;
   9734: result <= 12'b101110001010;
   9735: result <= 12'b101110001010;
   9736: result <= 12'b101110001001;
   9737: result <= 12'b101110001000;
   9738: result <= 12'b101110001000;
   9739: result <= 12'b101110000111;
   9740: result <= 12'b101110000110;
   9741: result <= 12'b101110000110;
   9742: result <= 12'b101110000101;
   9743: result <= 12'b101110000100;
   9744: result <= 12'b101110000100;
   9745: result <= 12'b101110000011;
   9746: result <= 12'b101110000010;
   9747: result <= 12'b101110000010;
   9748: result <= 12'b101110000001;
   9749: result <= 12'b101110000001;
   9750: result <= 12'b101110000000;
   9751: result <= 12'b101101111111;
   9752: result <= 12'b101101111111;
   9753: result <= 12'b101101111110;
   9754: result <= 12'b101101111101;
   9755: result <= 12'b101101111101;
   9756: result <= 12'b101101111100;
   9757: result <= 12'b101101111011;
   9758: result <= 12'b101101111011;
   9759: result <= 12'b101101111010;
   9760: result <= 12'b101101111001;
   9761: result <= 12'b101101111001;
   9762: result <= 12'b101101111000;
   9763: result <= 12'b101101110111;
   9764: result <= 12'b101101110111;
   9765: result <= 12'b101101110110;
   9766: result <= 12'b101101110101;
   9767: result <= 12'b101101110101;
   9768: result <= 12'b101101110100;
   9769: result <= 12'b101101110100;
   9770: result <= 12'b101101110011;
   9771: result <= 12'b101101110010;
   9772: result <= 12'b101101110010;
   9773: result <= 12'b101101110001;
   9774: result <= 12'b101101110000;
   9775: result <= 12'b101101110000;
   9776: result <= 12'b101101101111;
   9777: result <= 12'b101101101110;
   9778: result <= 12'b101101101110;
   9779: result <= 12'b101101101101;
   9780: result <= 12'b101101101100;
   9781: result <= 12'b101101101100;
   9782: result <= 12'b101101101011;
   9783: result <= 12'b101101101011;
   9784: result <= 12'b101101101010;
   9785: result <= 12'b101101101001;
   9786: result <= 12'b101101101001;
   9787: result <= 12'b101101101000;
   9788: result <= 12'b101101100111;
   9789: result <= 12'b101101100111;
   9790: result <= 12'b101101100110;
   9791: result <= 12'b101101100101;
   9792: result <= 12'b101101100101;
   9793: result <= 12'b101101100100;
   9794: result <= 12'b101101100011;
   9795: result <= 12'b101101100011;
   9796: result <= 12'b101101100010;
   9797: result <= 12'b101101100010;
   9798: result <= 12'b101101100001;
   9799: result <= 12'b101101100000;
   9800: result <= 12'b101101100000;
   9801: result <= 12'b101101011111;
   9802: result <= 12'b101101011110;
   9803: result <= 12'b101101011110;
   9804: result <= 12'b101101011101;
   9805: result <= 12'b101101011100;
   9806: result <= 12'b101101011100;
   9807: result <= 12'b101101011011;
   9808: result <= 12'b101101011010;
   9809: result <= 12'b101101011010;
   9810: result <= 12'b101101011001;
   9811: result <= 12'b101101011001;
   9812: result <= 12'b101101011000;
   9813: result <= 12'b101101010111;
   9814: result <= 12'b101101010111;
   9815: result <= 12'b101101010110;
   9816: result <= 12'b101101010101;
   9817: result <= 12'b101101010101;
   9818: result <= 12'b101101010100;
   9819: result <= 12'b101101010011;
   9820: result <= 12'b101101010011;
   9821: result <= 12'b101101010010;
   9822: result <= 12'b101101010010;
   9823: result <= 12'b101101010001;
   9824: result <= 12'b101101010000;
   9825: result <= 12'b101101010000;
   9826: result <= 12'b101101001111;
   9827: result <= 12'b101101001110;
   9828: result <= 12'b101101001110;
   9829: result <= 12'b101101001101;
   9830: result <= 12'b101101001100;
   9831: result <= 12'b101101001100;
   9832: result <= 12'b101101001011;
   9833: result <= 12'b101101001011;
   9834: result <= 12'b101101001010;
   9835: result <= 12'b101101001001;
   9836: result <= 12'b101101001001;
   9837: result <= 12'b101101001000;
   9838: result <= 12'b101101000111;
   9839: result <= 12'b101101000111;
   9840: result <= 12'b101101000110;
   9841: result <= 12'b101101000101;
   9842: result <= 12'b101101000101;
   9843: result <= 12'b101101000100;
   9844: result <= 12'b101101000100;
   9845: result <= 12'b101101000011;
   9846: result <= 12'b101101000010;
   9847: result <= 12'b101101000010;
   9848: result <= 12'b101101000001;
   9849: result <= 12'b101101000000;
   9850: result <= 12'b101101000000;
   9851: result <= 12'b101100111111;
   9852: result <= 12'b101100111111;
   9853: result <= 12'b101100111110;
   9854: result <= 12'b101100111101;
   9855: result <= 12'b101100111101;
   9856: result <= 12'b101100111100;
   9857: result <= 12'b101100111011;
   9858: result <= 12'b101100111011;
   9859: result <= 12'b101100111010;
   9860: result <= 12'b101100111001;
   9861: result <= 12'b101100111001;
   9862: result <= 12'b101100111000;
   9863: result <= 12'b101100111000;
   9864: result <= 12'b101100110111;
   9865: result <= 12'b101100110110;
   9866: result <= 12'b101100110110;
   9867: result <= 12'b101100110101;
   9868: result <= 12'b101100110100;
   9869: result <= 12'b101100110100;
   9870: result <= 12'b101100110011;
   9871: result <= 12'b101100110011;
   9872: result <= 12'b101100110010;
   9873: result <= 12'b101100110001;
   9874: result <= 12'b101100110001;
   9875: result <= 12'b101100110000;
   9876: result <= 12'b101100101111;
   9877: result <= 12'b101100101111;
   9878: result <= 12'b101100101110;
   9879: result <= 12'b101100101110;
   9880: result <= 12'b101100101101;
   9881: result <= 12'b101100101100;
   9882: result <= 12'b101100101100;
   9883: result <= 12'b101100101011;
   9884: result <= 12'b101100101010;
   9885: result <= 12'b101100101010;
   9886: result <= 12'b101100101001;
   9887: result <= 12'b101100101001;
   9888: result <= 12'b101100101000;
   9889: result <= 12'b101100100111;
   9890: result <= 12'b101100100111;
   9891: result <= 12'b101100100110;
   9892: result <= 12'b101100100101;
   9893: result <= 12'b101100100101;
   9894: result <= 12'b101100100100;
   9895: result <= 12'b101100100100;
   9896: result <= 12'b101100100011;
   9897: result <= 12'b101100100010;
   9898: result <= 12'b101100100010;
   9899: result <= 12'b101100100001;
   9900: result <= 12'b101100100000;
   9901: result <= 12'b101100100000;
   9902: result <= 12'b101100011111;
   9903: result <= 12'b101100011111;
   9904: result <= 12'b101100011110;
   9905: result <= 12'b101100011101;
   9906: result <= 12'b101100011101;
   9907: result <= 12'b101100011100;
   9908: result <= 12'b101100011011;
   9909: result <= 12'b101100011011;
   9910: result <= 12'b101100011010;
   9911: result <= 12'b101100011010;
   9912: result <= 12'b101100011001;
   9913: result <= 12'b101100011000;
   9914: result <= 12'b101100011000;
   9915: result <= 12'b101100010111;
   9916: result <= 12'b101100010110;
   9917: result <= 12'b101100010110;
   9918: result <= 12'b101100010101;
   9919: result <= 12'b101100010101;
   9920: result <= 12'b101100010100;
   9921: result <= 12'b101100010011;
   9922: result <= 12'b101100010011;
   9923: result <= 12'b101100010010;
   9924: result <= 12'b101100010010;
   9925: result <= 12'b101100010001;
   9926: result <= 12'b101100010000;
   9927: result <= 12'b101100010000;
   9928: result <= 12'b101100001111;
   9929: result <= 12'b101100001110;
   9930: result <= 12'b101100001110;
   9931: result <= 12'b101100001101;
   9932: result <= 12'b101100001101;
   9933: result <= 12'b101100001100;
   9934: result <= 12'b101100001011;
   9935: result <= 12'b101100001011;
   9936: result <= 12'b101100001010;
   9937: result <= 12'b101100001010;
   9938: result <= 12'b101100001001;
   9939: result <= 12'b101100001000;
   9940: result <= 12'b101100001000;
   9941: result <= 12'b101100000111;
   9942: result <= 12'b101100000110;
   9943: result <= 12'b101100000110;
   9944: result <= 12'b101100000101;
   9945: result <= 12'b101100000101;
   9946: result <= 12'b101100000100;
   9947: result <= 12'b101100000011;
   9948: result <= 12'b101100000011;
   9949: result <= 12'b101100000010;
   9950: result <= 12'b101100000010;
   9951: result <= 12'b101100000001;
   9952: result <= 12'b101100000000;
   9953: result <= 12'b101100000000;
   9954: result <= 12'b101011111111;
   9955: result <= 12'b101011111110;
   9956: result <= 12'b101011111110;
   9957: result <= 12'b101011111101;
   9958: result <= 12'b101011111101;
   9959: result <= 12'b101011111100;
   9960: result <= 12'b101011111011;
   9961: result <= 12'b101011111011;
   9962: result <= 12'b101011111010;
   9963: result <= 12'b101011111010;
   9964: result <= 12'b101011111001;
   9965: result <= 12'b101011111000;
   9966: result <= 12'b101011111000;
   9967: result <= 12'b101011110111;
   9968: result <= 12'b101011110111;
   9969: result <= 12'b101011110110;
   9970: result <= 12'b101011110101;
   9971: result <= 12'b101011110101;
   9972: result <= 12'b101011110100;
   9973: result <= 12'b101011110011;
   9974: result <= 12'b101011110011;
   9975: result <= 12'b101011110010;
   9976: result <= 12'b101011110010;
   9977: result <= 12'b101011110001;
   9978: result <= 12'b101011110000;
   9979: result <= 12'b101011110000;
   9980: result <= 12'b101011101111;
   9981: result <= 12'b101011101111;
   9982: result <= 12'b101011101110;
   9983: result <= 12'b101011101101;
   9984: result <= 12'b101011101101;
   9985: result <= 12'b101011101100;
   9986: result <= 12'b101011101100;
   9987: result <= 12'b101011101011;
   9988: result <= 12'b101011101010;
   9989: result <= 12'b101011101010;
   9990: result <= 12'b101011101001;
   9991: result <= 12'b101011101001;
   9992: result <= 12'b101011101000;
   9993: result <= 12'b101011100111;
   9994: result <= 12'b101011100111;
   9995: result <= 12'b101011100110;
   9996: result <= 12'b101011100101;
   9997: result <= 12'b101011100101;
   9998: result <= 12'b101011100100;
   9999: result <= 12'b101011100100;
   10000: result <= 12'b101011100011;
   10001: result <= 12'b101011100010;
   10002: result <= 12'b101011100010;
   10003: result <= 12'b101011100001;
   10004: result <= 12'b101011100001;
   10005: result <= 12'b101011100000;
   10006: result <= 12'b101011011111;
   10007: result <= 12'b101011011111;
   10008: result <= 12'b101011011110;
   10009: result <= 12'b101011011110;
   10010: result <= 12'b101011011101;
   10011: result <= 12'b101011011100;
   10012: result <= 12'b101011011100;
   10013: result <= 12'b101011011011;
   10014: result <= 12'b101011011011;
   10015: result <= 12'b101011011010;
   10016: result <= 12'b101011011001;
   10017: result <= 12'b101011011001;
   10018: result <= 12'b101011011000;
   10019: result <= 12'b101011011000;
   10020: result <= 12'b101011010111;
   10021: result <= 12'b101011010110;
   10022: result <= 12'b101011010110;
   10023: result <= 12'b101011010101;
   10024: result <= 12'b101011010101;
   10025: result <= 12'b101011010100;
   10026: result <= 12'b101011010011;
   10027: result <= 12'b101011010011;
   10028: result <= 12'b101011010010;
   10029: result <= 12'b101011010010;
   10030: result <= 12'b101011010001;
   10031: result <= 12'b101011010000;
   10032: result <= 12'b101011010000;
   10033: result <= 12'b101011001111;
   10034: result <= 12'b101011001111;
   10035: result <= 12'b101011001110;
   10036: result <= 12'b101011001101;
   10037: result <= 12'b101011001101;
   10038: result <= 12'b101011001100;
   10039: result <= 12'b101011001100;
   10040: result <= 12'b101011001011;
   10041: result <= 12'b101011001010;
   10042: result <= 12'b101011001010;
   10043: result <= 12'b101011001001;
   10044: result <= 12'b101011001001;
   10045: result <= 12'b101011001000;
   10046: result <= 12'b101011000111;
   10047: result <= 12'b101011000111;
   10048: result <= 12'b101011000110;
   10049: result <= 12'b101011000110;
   10050: result <= 12'b101011000101;
   10051: result <= 12'b101011000101;
   10052: result <= 12'b101011000100;
   10053: result <= 12'b101011000011;
   10054: result <= 12'b101011000011;
   10055: result <= 12'b101011000010;
   10056: result <= 12'b101011000010;
   10057: result <= 12'b101011000001;
   10058: result <= 12'b101011000000;
   10059: result <= 12'b101011000000;
   10060: result <= 12'b101010111111;
   10061: result <= 12'b101010111111;
   10062: result <= 12'b101010111110;
   10063: result <= 12'b101010111101;
   10064: result <= 12'b101010111101;
   10065: result <= 12'b101010111100;
   10066: result <= 12'b101010111100;
   10067: result <= 12'b101010111011;
   10068: result <= 12'b101010111010;
   10069: result <= 12'b101010111010;
   10070: result <= 12'b101010111001;
   10071: result <= 12'b101010111001;
   10072: result <= 12'b101010111000;
   10073: result <= 12'b101010110111;
   10074: result <= 12'b101010110111;
   10075: result <= 12'b101010110110;
   10076: result <= 12'b101010110110;
   10077: result <= 12'b101010110101;
   10078: result <= 12'b101010110101;
   10079: result <= 12'b101010110100;
   10080: result <= 12'b101010110011;
   10081: result <= 12'b101010110011;
   10082: result <= 12'b101010110010;
   10083: result <= 12'b101010110010;
   10084: result <= 12'b101010110001;
   10085: result <= 12'b101010110000;
   10086: result <= 12'b101010110000;
   10087: result <= 12'b101010101111;
   10088: result <= 12'b101010101111;
   10089: result <= 12'b101010101110;
   10090: result <= 12'b101010101101;
   10091: result <= 12'b101010101101;
   10092: result <= 12'b101010101100;
   10093: result <= 12'b101010101100;
   10094: result <= 12'b101010101011;
   10095: result <= 12'b101010101011;
   10096: result <= 12'b101010101010;
   10097: result <= 12'b101010101001;
   10098: result <= 12'b101010101001;
   10099: result <= 12'b101010101000;
   10100: result <= 12'b101010101000;
   10101: result <= 12'b101010100111;
   10102: result <= 12'b101010100110;
   10103: result <= 12'b101010100110;
   10104: result <= 12'b101010100101;
   10105: result <= 12'b101010100101;
   10106: result <= 12'b101010100100;
   10107: result <= 12'b101010100100;
   10108: result <= 12'b101010100011;
   10109: result <= 12'b101010100010;
   10110: result <= 12'b101010100010;
   10111: result <= 12'b101010100001;
   10112: result <= 12'b101010100001;
   10113: result <= 12'b101010100000;
   10114: result <= 12'b101010011111;
   10115: result <= 12'b101010011111;
   10116: result <= 12'b101010011110;
   10117: result <= 12'b101010011110;
   10118: result <= 12'b101010011101;
   10119: result <= 12'b101010011101;
   10120: result <= 12'b101010011100;
   10121: result <= 12'b101010011011;
   10122: result <= 12'b101010011011;
   10123: result <= 12'b101010011010;
   10124: result <= 12'b101010011010;
   10125: result <= 12'b101010011001;
   10126: result <= 12'b101010011001;
   10127: result <= 12'b101010011000;
   10128: result <= 12'b101010010111;
   10129: result <= 12'b101010010111;
   10130: result <= 12'b101010010110;
   10131: result <= 12'b101010010110;
   10132: result <= 12'b101010010101;
   10133: result <= 12'b101010010100;
   10134: result <= 12'b101010010100;
   10135: result <= 12'b101010010011;
   10136: result <= 12'b101010010011;
   10137: result <= 12'b101010010010;
   10138: result <= 12'b101010010010;
   10139: result <= 12'b101010010001;
   10140: result <= 12'b101010010000;
   10141: result <= 12'b101010010000;
   10142: result <= 12'b101010001111;
   10143: result <= 12'b101010001111;
   10144: result <= 12'b101010001110;
   10145: result <= 12'b101010001110;
   10146: result <= 12'b101010001101;
   10147: result <= 12'b101010001100;
   10148: result <= 12'b101010001100;
   10149: result <= 12'b101010001011;
   10150: result <= 12'b101010001011;
   10151: result <= 12'b101010001010;
   10152: result <= 12'b101010001010;
   10153: result <= 12'b101010001001;
   10154: result <= 12'b101010001000;
   10155: result <= 12'b101010001000;
   10156: result <= 12'b101010000111;
   10157: result <= 12'b101010000111;
   10158: result <= 12'b101010000110;
   10159: result <= 12'b101010000110;
   10160: result <= 12'b101010000101;
   10161: result <= 12'b101010000100;
   10162: result <= 12'b101010000100;
   10163: result <= 12'b101010000011;
   10164: result <= 12'b101010000011;
   10165: result <= 12'b101010000010;
   10166: result <= 12'b101010000010;
   10167: result <= 12'b101010000001;
   10168: result <= 12'b101010000000;
   10169: result <= 12'b101010000000;
   10170: result <= 12'b101001111111;
   10171: result <= 12'b101001111111;
   10172: result <= 12'b101001111110;
   10173: result <= 12'b101001111110;
   10174: result <= 12'b101001111101;
   10175: result <= 12'b101001111100;
   10176: result <= 12'b101001111100;
   10177: result <= 12'b101001111011;
   10178: result <= 12'b101001111011;
   10179: result <= 12'b101001111010;
   10180: result <= 12'b101001111010;
   10181: result <= 12'b101001111001;
   10182: result <= 12'b101001111000;
   10183: result <= 12'b101001111000;
   10184: result <= 12'b101001110111;
   10185: result <= 12'b101001110111;
   10186: result <= 12'b101001110110;
   10187: result <= 12'b101001110110;
   10188: result <= 12'b101001110101;
   10189: result <= 12'b101001110100;
   10190: result <= 12'b101001110100;
   10191: result <= 12'b101001110011;
   10192: result <= 12'b101001110011;
   10193: result <= 12'b101001110010;
   10194: result <= 12'b101001110010;
   10195: result <= 12'b101001110001;
   10196: result <= 12'b101001110000;
   10197: result <= 12'b101001110000;
   10198: result <= 12'b101001101111;
   10199: result <= 12'b101001101111;
   10200: result <= 12'b101001101110;
   10201: result <= 12'b101001101110;
   10202: result <= 12'b101001101101;
   10203: result <= 12'b101001101101;
   10204: result <= 12'b101001101100;
   10205: result <= 12'b101001101011;
   10206: result <= 12'b101001101011;
   10207: result <= 12'b101001101010;
   10208: result <= 12'b101001101010;
   10209: result <= 12'b101001101001;
   10210: result <= 12'b101001101001;
   10211: result <= 12'b101001101000;
   10212: result <= 12'b101001100111;
   10213: result <= 12'b101001100111;
   10214: result <= 12'b101001100110;
   10215: result <= 12'b101001100110;
   10216: result <= 12'b101001100101;
   10217: result <= 12'b101001100101;
   10218: result <= 12'b101001100100;
   10219: result <= 12'b101001100100;
   10220: result <= 12'b101001100011;
   10221: result <= 12'b101001100010;
   10222: result <= 12'b101001100010;
   10223: result <= 12'b101001100001;
   10224: result <= 12'b101001100001;
   10225: result <= 12'b101001100000;
   10226: result <= 12'b101001100000;
   10227: result <= 12'b101001011111;
   10228: result <= 12'b101001011111;
   10229: result <= 12'b101001011110;
   10230: result <= 12'b101001011101;
   10231: result <= 12'b101001011101;
   10232: result <= 12'b101001011100;
   10233: result <= 12'b101001011100;
   10234: result <= 12'b101001011011;
   10235: result <= 12'b101001011011;
   10236: result <= 12'b101001011010;
   10237: result <= 12'b101001011010;
   10238: result <= 12'b101001011001;
   10239: result <= 12'b101001011000;
   10240: result <= 12'b101001011000;
   10241: result <= 12'b101001010111;
   10242: result <= 12'b101001010111;
   10243: result <= 12'b101001010110;
   10244: result <= 12'b101001010110;
   10245: result <= 12'b101001010101;
   10246: result <= 12'b101001010101;
   10247: result <= 12'b101001010100;
   10248: result <= 12'b101001010011;
   10249: result <= 12'b101001010011;
   10250: result <= 12'b101001010010;
   10251: result <= 12'b101001010010;
   10252: result <= 12'b101001010001;
   10253: result <= 12'b101001010001;
   10254: result <= 12'b101001010000;
   10255: result <= 12'b101001010000;
   10256: result <= 12'b101001001111;
   10257: result <= 12'b101001001110;
   10258: result <= 12'b101001001110;
   10259: result <= 12'b101001001101;
   10260: result <= 12'b101001001101;
   10261: result <= 12'b101001001100;
   10262: result <= 12'b101001001100;
   10263: result <= 12'b101001001011;
   10264: result <= 12'b101001001011;
   10265: result <= 12'b101001001010;
   10266: result <= 12'b101001001001;
   10267: result <= 12'b101001001001;
   10268: result <= 12'b101001001000;
   10269: result <= 12'b101001001000;
   10270: result <= 12'b101001000111;
   10271: result <= 12'b101001000111;
   10272: result <= 12'b101001000110;
   10273: result <= 12'b101001000110;
   10274: result <= 12'b101001000101;
   10275: result <= 12'b101001000101;
   10276: result <= 12'b101001000100;
   10277: result <= 12'b101001000011;
   10278: result <= 12'b101001000011;
   10279: result <= 12'b101001000010;
   10280: result <= 12'b101001000010;
   10281: result <= 12'b101001000001;
   10282: result <= 12'b101001000001;
   10283: result <= 12'b101001000000;
   10284: result <= 12'b101001000000;
   10285: result <= 12'b101000111111;
   10286: result <= 12'b101000111111;
   10287: result <= 12'b101000111110;
   10288: result <= 12'b101000111101;
   10289: result <= 12'b101000111101;
   10290: result <= 12'b101000111100;
   10291: result <= 12'b101000111100;
   10292: result <= 12'b101000111011;
   10293: result <= 12'b101000111011;
   10294: result <= 12'b101000111010;
   10295: result <= 12'b101000111010;
   10296: result <= 12'b101000111001;
   10297: result <= 12'b101000111001;
   10298: result <= 12'b101000111000;
   10299: result <= 12'b101000110111;
   10300: result <= 12'b101000110111;
   10301: result <= 12'b101000110110;
   10302: result <= 12'b101000110110;
   10303: result <= 12'b101000110101;
   10304: result <= 12'b101000110101;
   10305: result <= 12'b101000110100;
   10306: result <= 12'b101000110100;
   10307: result <= 12'b101000110011;
   10308: result <= 12'b101000110011;
   10309: result <= 12'b101000110010;
   10310: result <= 12'b101000110001;
   10311: result <= 12'b101000110001;
   10312: result <= 12'b101000110000;
   10313: result <= 12'b101000110000;
   10314: result <= 12'b101000101111;
   10315: result <= 12'b101000101111;
   10316: result <= 12'b101000101110;
   10317: result <= 12'b101000101110;
   10318: result <= 12'b101000101101;
   10319: result <= 12'b101000101101;
   10320: result <= 12'b101000101100;
   10321: result <= 12'b101000101100;
   10322: result <= 12'b101000101011;
   10323: result <= 12'b101000101010;
   10324: result <= 12'b101000101010;
   10325: result <= 12'b101000101001;
   10326: result <= 12'b101000101001;
   10327: result <= 12'b101000101000;
   10328: result <= 12'b101000101000;
   10329: result <= 12'b101000100111;
   10330: result <= 12'b101000100111;
   10331: result <= 12'b101000100110;
   10332: result <= 12'b101000100110;
   10333: result <= 12'b101000100101;
   10334: result <= 12'b101000100101;
   10335: result <= 12'b101000100100;
   10336: result <= 12'b101000100100;
   10337: result <= 12'b101000100011;
   10338: result <= 12'b101000100010;
   10339: result <= 12'b101000100010;
   10340: result <= 12'b101000100001;
   10341: result <= 12'b101000100001;
   10342: result <= 12'b101000100000;
   10343: result <= 12'b101000100000;
   10344: result <= 12'b101000011111;
   10345: result <= 12'b101000011111;
   10346: result <= 12'b101000011110;
   10347: result <= 12'b101000011110;
   10348: result <= 12'b101000011101;
   10349: result <= 12'b101000011101;
   10350: result <= 12'b101000011100;
   10351: result <= 12'b101000011100;
   10352: result <= 12'b101000011011;
   10353: result <= 12'b101000011010;
   10354: result <= 12'b101000011010;
   10355: result <= 12'b101000011001;
   10356: result <= 12'b101000011001;
   10357: result <= 12'b101000011000;
   10358: result <= 12'b101000011000;
   10359: result <= 12'b101000010111;
   10360: result <= 12'b101000010111;
   10361: result <= 12'b101000010110;
   10362: result <= 12'b101000010110;
   10363: result <= 12'b101000010101;
   10364: result <= 12'b101000010101;
   10365: result <= 12'b101000010100;
   10366: result <= 12'b101000010100;
   10367: result <= 12'b101000010011;
   10368: result <= 12'b101000010011;
   10369: result <= 12'b101000010010;
   10370: result <= 12'b101000010001;
   10371: result <= 12'b101000010001;
   10372: result <= 12'b101000010000;
   10373: result <= 12'b101000010000;
   10374: result <= 12'b101000001111;
   10375: result <= 12'b101000001111;
   10376: result <= 12'b101000001110;
   10377: result <= 12'b101000001110;
   10378: result <= 12'b101000001101;
   10379: result <= 12'b101000001101;
   10380: result <= 12'b101000001100;
   10381: result <= 12'b101000001100;
   10382: result <= 12'b101000001011;
   10383: result <= 12'b101000001011;
   10384: result <= 12'b101000001010;
   10385: result <= 12'b101000001010;
   10386: result <= 12'b101000001001;
   10387: result <= 12'b101000001001;
   10388: result <= 12'b101000001000;
   10389: result <= 12'b101000001000;
   10390: result <= 12'b101000000111;
   10391: result <= 12'b101000000110;
   10392: result <= 12'b101000000110;
   10393: result <= 12'b101000000101;
   10394: result <= 12'b101000000101;
   10395: result <= 12'b101000000100;
   10396: result <= 12'b101000000100;
   10397: result <= 12'b101000000011;
   10398: result <= 12'b101000000011;
   10399: result <= 12'b101000000010;
   10400: result <= 12'b101000000010;
   10401: result <= 12'b101000000001;
   10402: result <= 12'b101000000001;
   10403: result <= 12'b101000000000;
   10404: result <= 12'b101000000000;
   10405: result <= 12'b100111111111;
   10406: result <= 12'b100111111111;
   10407: result <= 12'b100111111110;
   10408: result <= 12'b100111111110;
   10409: result <= 12'b100111111101;
   10410: result <= 12'b100111111101;
   10411: result <= 12'b100111111100;
   10412: result <= 12'b100111111100;
   10413: result <= 12'b100111111011;
   10414: result <= 12'b100111111011;
   10415: result <= 12'b100111111010;
   10416: result <= 12'b100111111001;
   10417: result <= 12'b100111111001;
   10418: result <= 12'b100111111000;
   10419: result <= 12'b100111111000;
   10420: result <= 12'b100111110111;
   10421: result <= 12'b100111110111;
   10422: result <= 12'b100111110110;
   10423: result <= 12'b100111110110;
   10424: result <= 12'b100111110101;
   10425: result <= 12'b100111110101;
   10426: result <= 12'b100111110100;
   10427: result <= 12'b100111110100;
   10428: result <= 12'b100111110011;
   10429: result <= 12'b100111110011;
   10430: result <= 12'b100111110010;
   10431: result <= 12'b100111110010;
   10432: result <= 12'b100111110001;
   10433: result <= 12'b100111110001;
   10434: result <= 12'b100111110000;
   10435: result <= 12'b100111110000;
   10436: result <= 12'b100111101111;
   10437: result <= 12'b100111101111;
   10438: result <= 12'b100111101110;
   10439: result <= 12'b100111101110;
   10440: result <= 12'b100111101101;
   10441: result <= 12'b100111101101;
   10442: result <= 12'b100111101100;
   10443: result <= 12'b100111101100;
   10444: result <= 12'b100111101011;
   10445: result <= 12'b100111101011;
   10446: result <= 12'b100111101010;
   10447: result <= 12'b100111101010;
   10448: result <= 12'b100111101001;
   10449: result <= 12'b100111101001;
   10450: result <= 12'b100111101000;
   10451: result <= 12'b100111101000;
   10452: result <= 12'b100111100111;
   10453: result <= 12'b100111100111;
   10454: result <= 12'b100111100110;
   10455: result <= 12'b100111100101;
   10456: result <= 12'b100111100101;
   10457: result <= 12'b100111100100;
   10458: result <= 12'b100111100100;
   10459: result <= 12'b100111100011;
   10460: result <= 12'b100111100011;
   10461: result <= 12'b100111100010;
   10462: result <= 12'b100111100010;
   10463: result <= 12'b100111100001;
   10464: result <= 12'b100111100001;
   10465: result <= 12'b100111100000;
   10466: result <= 12'b100111100000;
   10467: result <= 12'b100111011111;
   10468: result <= 12'b100111011111;
   10469: result <= 12'b100111011110;
   10470: result <= 12'b100111011110;
   10471: result <= 12'b100111011101;
   10472: result <= 12'b100111011101;
   10473: result <= 12'b100111011100;
   10474: result <= 12'b100111011100;
   10475: result <= 12'b100111011011;
   10476: result <= 12'b100111011011;
   10477: result <= 12'b100111011010;
   10478: result <= 12'b100111011010;
   10479: result <= 12'b100111011001;
   10480: result <= 12'b100111011001;
   10481: result <= 12'b100111011000;
   10482: result <= 12'b100111011000;
   10483: result <= 12'b100111010111;
   10484: result <= 12'b100111010111;
   10485: result <= 12'b100111010110;
   10486: result <= 12'b100111010110;
   10487: result <= 12'b100111010101;
   10488: result <= 12'b100111010101;
   10489: result <= 12'b100111010100;
   10490: result <= 12'b100111010100;
   10491: result <= 12'b100111010011;
   10492: result <= 12'b100111010011;
   10493: result <= 12'b100111010010;
   10494: result <= 12'b100111010010;
   10495: result <= 12'b100111010001;
   10496: result <= 12'b100111010001;
   10497: result <= 12'b100111010000;
   10498: result <= 12'b100111010000;
   10499: result <= 12'b100111001111;
   10500: result <= 12'b100111001111;
   10501: result <= 12'b100111001110;
   10502: result <= 12'b100111001110;
   10503: result <= 12'b100111001101;
   10504: result <= 12'b100111001101;
   10505: result <= 12'b100111001100;
   10506: result <= 12'b100111001100;
   10507: result <= 12'b100111001011;
   10508: result <= 12'b100111001011;
   10509: result <= 12'b100111001010;
   10510: result <= 12'b100111001010;
   10511: result <= 12'b100111001001;
   10512: result <= 12'b100111001001;
   10513: result <= 12'b100111001000;
   10514: result <= 12'b100111001000;
   10515: result <= 12'b100111000111;
   10516: result <= 12'b100111000111;
   10517: result <= 12'b100111000110;
   10518: result <= 12'b100111000110;
   10519: result <= 12'b100111000101;
   10520: result <= 12'b100111000101;
   10521: result <= 12'b100111000100;
   10522: result <= 12'b100111000100;
   10523: result <= 12'b100111000100;
   10524: result <= 12'b100111000011;
   10525: result <= 12'b100111000011;
   10526: result <= 12'b100111000010;
   10527: result <= 12'b100111000010;
   10528: result <= 12'b100111000001;
   10529: result <= 12'b100111000001;
   10530: result <= 12'b100111000000;
   10531: result <= 12'b100111000000;
   10532: result <= 12'b100110111111;
   10533: result <= 12'b100110111111;
   10534: result <= 12'b100110111110;
   10535: result <= 12'b100110111110;
   10536: result <= 12'b100110111101;
   10537: result <= 12'b100110111101;
   10538: result <= 12'b100110111100;
   10539: result <= 12'b100110111100;
   10540: result <= 12'b100110111011;
   10541: result <= 12'b100110111011;
   10542: result <= 12'b100110111010;
   10543: result <= 12'b100110111010;
   10544: result <= 12'b100110111001;
   10545: result <= 12'b100110111001;
   10546: result <= 12'b100110111000;
   10547: result <= 12'b100110111000;
   10548: result <= 12'b100110110111;
   10549: result <= 12'b100110110111;
   10550: result <= 12'b100110110110;
   10551: result <= 12'b100110110110;
   10552: result <= 12'b100110110101;
   10553: result <= 12'b100110110101;
   10554: result <= 12'b100110110100;
   10555: result <= 12'b100110110100;
   10556: result <= 12'b100110110011;
   10557: result <= 12'b100110110011;
   10558: result <= 12'b100110110010;
   10559: result <= 12'b100110110010;
   10560: result <= 12'b100110110001;
   10561: result <= 12'b100110110001;
   10562: result <= 12'b100110110001;
   10563: result <= 12'b100110110000;
   10564: result <= 12'b100110110000;
   10565: result <= 12'b100110101111;
   10566: result <= 12'b100110101111;
   10567: result <= 12'b100110101110;
   10568: result <= 12'b100110101110;
   10569: result <= 12'b100110101101;
   10570: result <= 12'b100110101101;
   10571: result <= 12'b100110101100;
   10572: result <= 12'b100110101100;
   10573: result <= 12'b100110101011;
   10574: result <= 12'b100110101011;
   10575: result <= 12'b100110101010;
   10576: result <= 12'b100110101010;
   10577: result <= 12'b100110101001;
   10578: result <= 12'b100110101001;
   10579: result <= 12'b100110101000;
   10580: result <= 12'b100110101000;
   10581: result <= 12'b100110100111;
   10582: result <= 12'b100110100111;
   10583: result <= 12'b100110100110;
   10584: result <= 12'b100110100110;
   10585: result <= 12'b100110100101;
   10586: result <= 12'b100110100101;
   10587: result <= 12'b100110100101;
   10588: result <= 12'b100110100100;
   10589: result <= 12'b100110100100;
   10590: result <= 12'b100110100011;
   10591: result <= 12'b100110100011;
   10592: result <= 12'b100110100010;
   10593: result <= 12'b100110100010;
   10594: result <= 12'b100110100001;
   10595: result <= 12'b100110100001;
   10596: result <= 12'b100110100000;
   10597: result <= 12'b100110100000;
   10598: result <= 12'b100110011111;
   10599: result <= 12'b100110011111;
   10600: result <= 12'b100110011110;
   10601: result <= 12'b100110011110;
   10602: result <= 12'b100110011101;
   10603: result <= 12'b100110011101;
   10604: result <= 12'b100110011100;
   10605: result <= 12'b100110011100;
   10606: result <= 12'b100110011011;
   10607: result <= 12'b100110011011;
   10608: result <= 12'b100110011011;
   10609: result <= 12'b100110011010;
   10610: result <= 12'b100110011010;
   10611: result <= 12'b100110011001;
   10612: result <= 12'b100110011001;
   10613: result <= 12'b100110011000;
   10614: result <= 12'b100110011000;
   10615: result <= 12'b100110010111;
   10616: result <= 12'b100110010111;
   10617: result <= 12'b100110010110;
   10618: result <= 12'b100110010110;
   10619: result <= 12'b100110010101;
   10620: result <= 12'b100110010101;
   10621: result <= 12'b100110010100;
   10622: result <= 12'b100110010100;
   10623: result <= 12'b100110010011;
   10624: result <= 12'b100110010011;
   10625: result <= 12'b100110010011;
   10626: result <= 12'b100110010010;
   10627: result <= 12'b100110010010;
   10628: result <= 12'b100110010001;
   10629: result <= 12'b100110010001;
   10630: result <= 12'b100110010000;
   10631: result <= 12'b100110010000;
   10632: result <= 12'b100110001111;
   10633: result <= 12'b100110001111;
   10634: result <= 12'b100110001110;
   10635: result <= 12'b100110001110;
   10636: result <= 12'b100110001101;
   10637: result <= 12'b100110001101;
   10638: result <= 12'b100110001101;
   10639: result <= 12'b100110001100;
   10640: result <= 12'b100110001100;
   10641: result <= 12'b100110001011;
   10642: result <= 12'b100110001011;
   10643: result <= 12'b100110001010;
   10644: result <= 12'b100110001010;
   10645: result <= 12'b100110001001;
   10646: result <= 12'b100110001001;
   10647: result <= 12'b100110001000;
   10648: result <= 12'b100110001000;
   10649: result <= 12'b100110000111;
   10650: result <= 12'b100110000111;
   10651: result <= 12'b100110000110;
   10652: result <= 12'b100110000110;
   10653: result <= 12'b100110000110;
   10654: result <= 12'b100110000101;
   10655: result <= 12'b100110000101;
   10656: result <= 12'b100110000100;
   10657: result <= 12'b100110000100;
   10658: result <= 12'b100110000011;
   10659: result <= 12'b100110000011;
   10660: result <= 12'b100110000010;
   10661: result <= 12'b100110000010;
   10662: result <= 12'b100110000001;
   10663: result <= 12'b100110000001;
   10664: result <= 12'b100110000001;
   10665: result <= 12'b100110000000;
   10666: result <= 12'b100110000000;
   10667: result <= 12'b100101111111;
   10668: result <= 12'b100101111111;
   10669: result <= 12'b100101111110;
   10670: result <= 12'b100101111110;
   10671: result <= 12'b100101111101;
   10672: result <= 12'b100101111101;
   10673: result <= 12'b100101111100;
   10674: result <= 12'b100101111100;
   10675: result <= 12'b100101111011;
   10676: result <= 12'b100101111011;
   10677: result <= 12'b100101111011;
   10678: result <= 12'b100101111010;
   10679: result <= 12'b100101111010;
   10680: result <= 12'b100101111001;
   10681: result <= 12'b100101111001;
   10682: result <= 12'b100101111000;
   10683: result <= 12'b100101111000;
   10684: result <= 12'b100101110111;
   10685: result <= 12'b100101110111;
   10686: result <= 12'b100101110110;
   10687: result <= 12'b100101110110;
   10688: result <= 12'b100101110110;
   10689: result <= 12'b100101110101;
   10690: result <= 12'b100101110101;
   10691: result <= 12'b100101110100;
   10692: result <= 12'b100101110100;
   10693: result <= 12'b100101110011;
   10694: result <= 12'b100101110011;
   10695: result <= 12'b100101110010;
   10696: result <= 12'b100101110010;
   10697: result <= 12'b100101110010;
   10698: result <= 12'b100101110001;
   10699: result <= 12'b100101110001;
   10700: result <= 12'b100101110000;
   10701: result <= 12'b100101110000;
   10702: result <= 12'b100101101111;
   10703: result <= 12'b100101101111;
   10704: result <= 12'b100101101110;
   10705: result <= 12'b100101101110;
   10706: result <= 12'b100101101101;
   10707: result <= 12'b100101101101;
   10708: result <= 12'b100101101101;
   10709: result <= 12'b100101101100;
   10710: result <= 12'b100101101100;
   10711: result <= 12'b100101101011;
   10712: result <= 12'b100101101011;
   10713: result <= 12'b100101101010;
   10714: result <= 12'b100101101010;
   10715: result <= 12'b100101101001;
   10716: result <= 12'b100101101001;
   10717: result <= 12'b100101101001;
   10718: result <= 12'b100101101000;
   10719: result <= 12'b100101101000;
   10720: result <= 12'b100101100111;
   10721: result <= 12'b100101100111;
   10722: result <= 12'b100101100110;
   10723: result <= 12'b100101100110;
   10724: result <= 12'b100101100101;
   10725: result <= 12'b100101100101;
   10726: result <= 12'b100101100101;
   10727: result <= 12'b100101100100;
   10728: result <= 12'b100101100100;
   10729: result <= 12'b100101100011;
   10730: result <= 12'b100101100011;
   10731: result <= 12'b100101100010;
   10732: result <= 12'b100101100010;
   10733: result <= 12'b100101100001;
   10734: result <= 12'b100101100001;
   10735: result <= 12'b100101100001;
   10736: result <= 12'b100101100000;
   10737: result <= 12'b100101100000;
   10738: result <= 12'b100101011111;
   10739: result <= 12'b100101011111;
   10740: result <= 12'b100101011110;
   10741: result <= 12'b100101011110;
   10742: result <= 12'b100101011110;
   10743: result <= 12'b100101011101;
   10744: result <= 12'b100101011101;
   10745: result <= 12'b100101011100;
   10746: result <= 12'b100101011100;
   10747: result <= 12'b100101011011;
   10748: result <= 12'b100101011011;
   10749: result <= 12'b100101011010;
   10750: result <= 12'b100101011010;
   10751: result <= 12'b100101011010;
   10752: result <= 12'b100101011001;
   10753: result <= 12'b100101011001;
   10754: result <= 12'b100101011000;
   10755: result <= 12'b100101011000;
   10756: result <= 12'b100101010111;
   10757: result <= 12'b100101010111;
   10758: result <= 12'b100101010111;
   10759: result <= 12'b100101010110;
   10760: result <= 12'b100101010110;
   10761: result <= 12'b100101010101;
   10762: result <= 12'b100101010101;
   10763: result <= 12'b100101010100;
   10764: result <= 12'b100101010100;
   10765: result <= 12'b100101010011;
   10766: result <= 12'b100101010011;
   10767: result <= 12'b100101010011;
   10768: result <= 12'b100101010010;
   10769: result <= 12'b100101010010;
   10770: result <= 12'b100101010001;
   10771: result <= 12'b100101010001;
   10772: result <= 12'b100101010000;
   10773: result <= 12'b100101010000;
   10774: result <= 12'b100101010000;
   10775: result <= 12'b100101001111;
   10776: result <= 12'b100101001111;
   10777: result <= 12'b100101001110;
   10778: result <= 12'b100101001110;
   10779: result <= 12'b100101001101;
   10780: result <= 12'b100101001101;
   10781: result <= 12'b100101001101;
   10782: result <= 12'b100101001100;
   10783: result <= 12'b100101001100;
   10784: result <= 12'b100101001011;
   10785: result <= 12'b100101001011;
   10786: result <= 12'b100101001010;
   10787: result <= 12'b100101001010;
   10788: result <= 12'b100101001010;
   10789: result <= 12'b100101001001;
   10790: result <= 12'b100101001001;
   10791: result <= 12'b100101001000;
   10792: result <= 12'b100101001000;
   10793: result <= 12'b100101000111;
   10794: result <= 12'b100101000111;
   10795: result <= 12'b100101000111;
   10796: result <= 12'b100101000110;
   10797: result <= 12'b100101000110;
   10798: result <= 12'b100101000101;
   10799: result <= 12'b100101000101;
   10800: result <= 12'b100101000100;
   10801: result <= 12'b100101000100;
   10802: result <= 12'b100101000100;
   10803: result <= 12'b100101000011;
   10804: result <= 12'b100101000011;
   10805: result <= 12'b100101000010;
   10806: result <= 12'b100101000010;
   10807: result <= 12'b100101000010;
   10808: result <= 12'b100101000001;
   10809: result <= 12'b100101000001;
   10810: result <= 12'b100101000000;
   10811: result <= 12'b100101000000;
   10812: result <= 12'b100100111111;
   10813: result <= 12'b100100111111;
   10814: result <= 12'b100100111111;
   10815: result <= 12'b100100111110;
   10816: result <= 12'b100100111110;
   10817: result <= 12'b100100111101;
   10818: result <= 12'b100100111101;
   10819: result <= 12'b100100111100;
   10820: result <= 12'b100100111100;
   10821: result <= 12'b100100111100;
   10822: result <= 12'b100100111011;
   10823: result <= 12'b100100111011;
   10824: result <= 12'b100100111010;
   10825: result <= 12'b100100111010;
   10826: result <= 12'b100100111010;
   10827: result <= 12'b100100111001;
   10828: result <= 12'b100100111001;
   10829: result <= 12'b100100111000;
   10830: result <= 12'b100100111000;
   10831: result <= 12'b100100110111;
   10832: result <= 12'b100100110111;
   10833: result <= 12'b100100110111;
   10834: result <= 12'b100100110110;
   10835: result <= 12'b100100110110;
   10836: result <= 12'b100100110101;
   10837: result <= 12'b100100110101;
   10838: result <= 12'b100100110101;
   10839: result <= 12'b100100110100;
   10840: result <= 12'b100100110100;
   10841: result <= 12'b100100110011;
   10842: result <= 12'b100100110011;
   10843: result <= 12'b100100110010;
   10844: result <= 12'b100100110010;
   10845: result <= 12'b100100110010;
   10846: result <= 12'b100100110001;
   10847: result <= 12'b100100110001;
   10848: result <= 12'b100100110000;
   10849: result <= 12'b100100110000;
   10850: result <= 12'b100100110000;
   10851: result <= 12'b100100101111;
   10852: result <= 12'b100100101111;
   10853: result <= 12'b100100101110;
   10854: result <= 12'b100100101110;
   10855: result <= 12'b100100101110;
   10856: result <= 12'b100100101101;
   10857: result <= 12'b100100101101;
   10858: result <= 12'b100100101100;
   10859: result <= 12'b100100101100;
   10860: result <= 12'b100100101011;
   10861: result <= 12'b100100101011;
   10862: result <= 12'b100100101011;
   10863: result <= 12'b100100101010;
   10864: result <= 12'b100100101010;
   10865: result <= 12'b100100101001;
   10866: result <= 12'b100100101001;
   10867: result <= 12'b100100101001;
   10868: result <= 12'b100100101000;
   10869: result <= 12'b100100101000;
   10870: result <= 12'b100100100111;
   10871: result <= 12'b100100100111;
   10872: result <= 12'b100100100111;
   10873: result <= 12'b100100100110;
   10874: result <= 12'b100100100110;
   10875: result <= 12'b100100100101;
   10876: result <= 12'b100100100101;
   10877: result <= 12'b100100100101;
   10878: result <= 12'b100100100100;
   10879: result <= 12'b100100100100;
   10880: result <= 12'b100100100011;
   10881: result <= 12'b100100100011;
   10882: result <= 12'b100100100011;
   10883: result <= 12'b100100100010;
   10884: result <= 12'b100100100010;
   10885: result <= 12'b100100100001;
   10886: result <= 12'b100100100001;
   10887: result <= 12'b100100100001;
   10888: result <= 12'b100100100000;
   10889: result <= 12'b100100100000;
   10890: result <= 12'b100100011111;
   10891: result <= 12'b100100011111;
   10892: result <= 12'b100100011111;
   10893: result <= 12'b100100011110;
   10894: result <= 12'b100100011110;
   10895: result <= 12'b100100011101;
   10896: result <= 12'b100100011101;
   10897: result <= 12'b100100011101;
   10898: result <= 12'b100100011100;
   10899: result <= 12'b100100011100;
   10900: result <= 12'b100100011011;
   10901: result <= 12'b100100011011;
   10902: result <= 12'b100100011011;
   10903: result <= 12'b100100011010;
   10904: result <= 12'b100100011010;
   10905: result <= 12'b100100011001;
   10906: result <= 12'b100100011001;
   10907: result <= 12'b100100011001;
   10908: result <= 12'b100100011000;
   10909: result <= 12'b100100011000;
   10910: result <= 12'b100100010111;
   10911: result <= 12'b100100010111;
   10912: result <= 12'b100100010111;
   10913: result <= 12'b100100010110;
   10914: result <= 12'b100100010110;
   10915: result <= 12'b100100010101;
   10916: result <= 12'b100100010101;
   10917: result <= 12'b100100010101;
   10918: result <= 12'b100100010100;
   10919: result <= 12'b100100010100;
   10920: result <= 12'b100100010011;
   10921: result <= 12'b100100010011;
   10922: result <= 12'b100100010011;
   10923: result <= 12'b100100010010;
   10924: result <= 12'b100100010010;
   10925: result <= 12'b100100010001;
   10926: result <= 12'b100100010001;
   10927: result <= 12'b100100010001;
   10928: result <= 12'b100100010000;
   10929: result <= 12'b100100010000;
   10930: result <= 12'b100100010000;
   10931: result <= 12'b100100001111;
   10932: result <= 12'b100100001111;
   10933: result <= 12'b100100001110;
   10934: result <= 12'b100100001110;
   10935: result <= 12'b100100001110;
   10936: result <= 12'b100100001101;
   10937: result <= 12'b100100001101;
   10938: result <= 12'b100100001100;
   10939: result <= 12'b100100001100;
   10940: result <= 12'b100100001100;
   10941: result <= 12'b100100001011;
   10942: result <= 12'b100100001011;
   10943: result <= 12'b100100001010;
   10944: result <= 12'b100100001010;
   10945: result <= 12'b100100001010;
   10946: result <= 12'b100100001001;
   10947: result <= 12'b100100001001;
   10948: result <= 12'b100100001001;
   10949: result <= 12'b100100001000;
   10950: result <= 12'b100100001000;
   10951: result <= 12'b100100000111;
   10952: result <= 12'b100100000111;
   10953: result <= 12'b100100000111;
   10954: result <= 12'b100100000110;
   10955: result <= 12'b100100000110;
   10956: result <= 12'b100100000101;
   10957: result <= 12'b100100000101;
   10958: result <= 12'b100100000101;
   10959: result <= 12'b100100000100;
   10960: result <= 12'b100100000100;
   10961: result <= 12'b100100000100;
   10962: result <= 12'b100100000011;
   10963: result <= 12'b100100000011;
   10964: result <= 12'b100100000010;
   10965: result <= 12'b100100000010;
   10966: result <= 12'b100100000010;
   10967: result <= 12'b100100000001;
   10968: result <= 12'b100100000001;
   10969: result <= 12'b100100000000;
   10970: result <= 12'b100100000000;
   10971: result <= 12'b100100000000;
   10972: result <= 12'b100011111111;
   10973: result <= 12'b100011111111;
   10974: result <= 12'b100011111111;
   10975: result <= 12'b100011111110;
   10976: result <= 12'b100011111110;
   10977: result <= 12'b100011111101;
   10978: result <= 12'b100011111101;
   10979: result <= 12'b100011111101;
   10980: result <= 12'b100011111100;
   10981: result <= 12'b100011111100;
   10982: result <= 12'b100011111100;
   10983: result <= 12'b100011111011;
   10984: result <= 12'b100011111011;
   10985: result <= 12'b100011111010;
   10986: result <= 12'b100011111010;
   10987: result <= 12'b100011111010;
   10988: result <= 12'b100011111001;
   10989: result <= 12'b100011111001;
   10990: result <= 12'b100011111001;
   10991: result <= 12'b100011111000;
   10992: result <= 12'b100011111000;
   10993: result <= 12'b100011110111;
   10994: result <= 12'b100011110111;
   10995: result <= 12'b100011110111;
   10996: result <= 12'b100011110110;
   10997: result <= 12'b100011110110;
   10998: result <= 12'b100011110110;
   10999: result <= 12'b100011110101;
   11000: result <= 12'b100011110101;
   11001: result <= 12'b100011110100;
   11002: result <= 12'b100011110100;
   11003: result <= 12'b100011110100;
   11004: result <= 12'b100011110011;
   11005: result <= 12'b100011110011;
   11006: result <= 12'b100011110011;
   11007: result <= 12'b100011110010;
   11008: result <= 12'b100011110010;
   11009: result <= 12'b100011110001;
   11010: result <= 12'b100011110001;
   11011: result <= 12'b100011110001;
   11012: result <= 12'b100011110000;
   11013: result <= 12'b100011110000;
   11014: result <= 12'b100011110000;
   11015: result <= 12'b100011101111;
   11016: result <= 12'b100011101111;
   11017: result <= 12'b100011101111;
   11018: result <= 12'b100011101110;
   11019: result <= 12'b100011101110;
   11020: result <= 12'b100011101101;
   11021: result <= 12'b100011101101;
   11022: result <= 12'b100011101101;
   11023: result <= 12'b100011101100;
   11024: result <= 12'b100011101100;
   11025: result <= 12'b100011101100;
   11026: result <= 12'b100011101011;
   11027: result <= 12'b100011101011;
   11028: result <= 12'b100011101010;
   11029: result <= 12'b100011101010;
   11030: result <= 12'b100011101010;
   11031: result <= 12'b100011101001;
   11032: result <= 12'b100011101001;
   11033: result <= 12'b100011101001;
   11034: result <= 12'b100011101000;
   11035: result <= 12'b100011101000;
   11036: result <= 12'b100011101000;
   11037: result <= 12'b100011100111;
   11038: result <= 12'b100011100111;
   11039: result <= 12'b100011100110;
   11040: result <= 12'b100011100110;
   11041: result <= 12'b100011100110;
   11042: result <= 12'b100011100101;
   11043: result <= 12'b100011100101;
   11044: result <= 12'b100011100101;
   11045: result <= 12'b100011100100;
   11046: result <= 12'b100011100100;
   11047: result <= 12'b100011100100;
   11048: result <= 12'b100011100011;
   11049: result <= 12'b100011100011;
   11050: result <= 12'b100011100011;
   11051: result <= 12'b100011100010;
   11052: result <= 12'b100011100010;
   11053: result <= 12'b100011100001;
   11054: result <= 12'b100011100001;
   11055: result <= 12'b100011100001;
   11056: result <= 12'b100011100000;
   11057: result <= 12'b100011100000;
   11058: result <= 12'b100011100000;
   11059: result <= 12'b100011011111;
   11060: result <= 12'b100011011111;
   11061: result <= 12'b100011011111;
   11062: result <= 12'b100011011110;
   11063: result <= 12'b100011011110;
   11064: result <= 12'b100011011110;
   11065: result <= 12'b100011011101;
   11066: result <= 12'b100011011101;
   11067: result <= 12'b100011011100;
   11068: result <= 12'b100011011100;
   11069: result <= 12'b100011011100;
   11070: result <= 12'b100011011011;
   11071: result <= 12'b100011011011;
   11072: result <= 12'b100011011011;
   11073: result <= 12'b100011011010;
   11074: result <= 12'b100011011010;
   11075: result <= 12'b100011011010;
   11076: result <= 12'b100011011001;
   11077: result <= 12'b100011011001;
   11078: result <= 12'b100011011001;
   11079: result <= 12'b100011011000;
   11080: result <= 12'b100011011000;
   11081: result <= 12'b100011011000;
   11082: result <= 12'b100011010111;
   11083: result <= 12'b100011010111;
   11084: result <= 12'b100011010110;
   11085: result <= 12'b100011010110;
   11086: result <= 12'b100011010110;
   11087: result <= 12'b100011010101;
   11088: result <= 12'b100011010101;
   11089: result <= 12'b100011010101;
   11090: result <= 12'b100011010100;
   11091: result <= 12'b100011010100;
   11092: result <= 12'b100011010100;
   11093: result <= 12'b100011010011;
   11094: result <= 12'b100011010011;
   11095: result <= 12'b100011010011;
   11096: result <= 12'b100011010010;
   11097: result <= 12'b100011010010;
   11098: result <= 12'b100011010010;
   11099: result <= 12'b100011010001;
   11100: result <= 12'b100011010001;
   11101: result <= 12'b100011010001;
   11102: result <= 12'b100011010000;
   11103: result <= 12'b100011010000;
   11104: result <= 12'b100011010000;
   11105: result <= 12'b100011001111;
   11106: result <= 12'b100011001111;
   11107: result <= 12'b100011001110;
   11108: result <= 12'b100011001110;
   11109: result <= 12'b100011001110;
   11110: result <= 12'b100011001101;
   11111: result <= 12'b100011001101;
   11112: result <= 12'b100011001101;
   11113: result <= 12'b100011001100;
   11114: result <= 12'b100011001100;
   11115: result <= 12'b100011001100;
   11116: result <= 12'b100011001011;
   11117: result <= 12'b100011001011;
   11118: result <= 12'b100011001011;
   11119: result <= 12'b100011001010;
   11120: result <= 12'b100011001010;
   11121: result <= 12'b100011001010;
   11122: result <= 12'b100011001001;
   11123: result <= 12'b100011001001;
   11124: result <= 12'b100011001001;
   11125: result <= 12'b100011001000;
   11126: result <= 12'b100011001000;
   11127: result <= 12'b100011001000;
   11128: result <= 12'b100011000111;
   11129: result <= 12'b100011000111;
   11130: result <= 12'b100011000111;
   11131: result <= 12'b100011000110;
   11132: result <= 12'b100011000110;
   11133: result <= 12'b100011000110;
   11134: result <= 12'b100011000101;
   11135: result <= 12'b100011000101;
   11136: result <= 12'b100011000101;
   11137: result <= 12'b100011000100;
   11138: result <= 12'b100011000100;
   11139: result <= 12'b100011000100;
   11140: result <= 12'b100011000011;
   11141: result <= 12'b100011000011;
   11142: result <= 12'b100011000011;
   11143: result <= 12'b100011000010;
   11144: result <= 12'b100011000010;
   11145: result <= 12'b100011000010;
   11146: result <= 12'b100011000001;
   11147: result <= 12'b100011000001;
   11148: result <= 12'b100011000001;
   11149: result <= 12'b100011000000;
   11150: result <= 12'b100011000000;
   11151: result <= 12'b100011000000;
   11152: result <= 12'b100010111111;
   11153: result <= 12'b100010111111;
   11154: result <= 12'b100010111111;
   11155: result <= 12'b100010111110;
   11156: result <= 12'b100010111110;
   11157: result <= 12'b100010111110;
   11158: result <= 12'b100010111101;
   11159: result <= 12'b100010111101;
   11160: result <= 12'b100010111101;
   11161: result <= 12'b100010111100;
   11162: result <= 12'b100010111100;
   11163: result <= 12'b100010111100;
   11164: result <= 12'b100010111011;
   11165: result <= 12'b100010111011;
   11166: result <= 12'b100010111011;
   11167: result <= 12'b100010111010;
   11168: result <= 12'b100010111010;
   11169: result <= 12'b100010111010;
   11170: result <= 12'b100010111001;
   11171: result <= 12'b100010111001;
   11172: result <= 12'b100010111001;
   11173: result <= 12'b100010111000;
   11174: result <= 12'b100010111000;
   11175: result <= 12'b100010111000;
   11176: result <= 12'b100010110111;
   11177: result <= 12'b100010110111;
   11178: result <= 12'b100010110111;
   11179: result <= 12'b100010110110;
   11180: result <= 12'b100010110110;
   11181: result <= 12'b100010110110;
   11182: result <= 12'b100010110101;
   11183: result <= 12'b100010110101;
   11184: result <= 12'b100010110101;
   11185: result <= 12'b100010110101;
   11186: result <= 12'b100010110100;
   11187: result <= 12'b100010110100;
   11188: result <= 12'b100010110100;
   11189: result <= 12'b100010110011;
   11190: result <= 12'b100010110011;
   11191: result <= 12'b100010110011;
   11192: result <= 12'b100010110010;
   11193: result <= 12'b100010110010;
   11194: result <= 12'b100010110010;
   11195: result <= 12'b100010110001;
   11196: result <= 12'b100010110001;
   11197: result <= 12'b100010110001;
   11198: result <= 12'b100010110000;
   11199: result <= 12'b100010110000;
   11200: result <= 12'b100010110000;
   11201: result <= 12'b100010101111;
   11202: result <= 12'b100010101111;
   11203: result <= 12'b100010101111;
   11204: result <= 12'b100010101110;
   11205: result <= 12'b100010101110;
   11206: result <= 12'b100010101110;
   11207: result <= 12'b100010101101;
   11208: result <= 12'b100010101101;
   11209: result <= 12'b100010101101;
   11210: result <= 12'b100010101101;
   11211: result <= 12'b100010101100;
   11212: result <= 12'b100010101100;
   11213: result <= 12'b100010101100;
   11214: result <= 12'b100010101011;
   11215: result <= 12'b100010101011;
   11216: result <= 12'b100010101011;
   11217: result <= 12'b100010101010;
   11218: result <= 12'b100010101010;
   11219: result <= 12'b100010101010;
   11220: result <= 12'b100010101001;
   11221: result <= 12'b100010101001;
   11222: result <= 12'b100010101001;
   11223: result <= 12'b100010101000;
   11224: result <= 12'b100010101000;
   11225: result <= 12'b100010101000;
   11226: result <= 12'b100010101000;
   11227: result <= 12'b100010100111;
   11228: result <= 12'b100010100111;
   11229: result <= 12'b100010100111;
   11230: result <= 12'b100010100110;
   11231: result <= 12'b100010100110;
   11232: result <= 12'b100010100110;
   11233: result <= 12'b100010100101;
   11234: result <= 12'b100010100101;
   11235: result <= 12'b100010100101;
   11236: result <= 12'b100010100100;
   11237: result <= 12'b100010100100;
   11238: result <= 12'b100010100100;
   11239: result <= 12'b100010100011;
   11240: result <= 12'b100010100011;
   11241: result <= 12'b100010100011;
   11242: result <= 12'b100010100011;
   11243: result <= 12'b100010100010;
   11244: result <= 12'b100010100010;
   11245: result <= 12'b100010100010;
   11246: result <= 12'b100010100001;
   11247: result <= 12'b100010100001;
   11248: result <= 12'b100010100001;
   11249: result <= 12'b100010100000;
   11250: result <= 12'b100010100000;
   11251: result <= 12'b100010100000;
   11252: result <= 12'b100010100000;
   11253: result <= 12'b100010011111;
   11254: result <= 12'b100010011111;
   11255: result <= 12'b100010011111;
   11256: result <= 12'b100010011110;
   11257: result <= 12'b100010011110;
   11258: result <= 12'b100010011110;
   11259: result <= 12'b100010011101;
   11260: result <= 12'b100010011101;
   11261: result <= 12'b100010011101;
   11262: result <= 12'b100010011100;
   11263: result <= 12'b100010011100;
   11264: result <= 12'b100010011100;
   11265: result <= 12'b100010011100;
   11266: result <= 12'b100010011011;
   11267: result <= 12'b100010011011;
   11268: result <= 12'b100010011011;
   11269: result <= 12'b100010011010;
   11270: result <= 12'b100010011010;
   11271: result <= 12'b100010011010;
   11272: result <= 12'b100010011001;
   11273: result <= 12'b100010011001;
   11274: result <= 12'b100010011001;
   11275: result <= 12'b100010011001;
   11276: result <= 12'b100010011000;
   11277: result <= 12'b100010011000;
   11278: result <= 12'b100010011000;
   11279: result <= 12'b100010010111;
   11280: result <= 12'b100010010111;
   11281: result <= 12'b100010010111;
   11282: result <= 12'b100010010111;
   11283: result <= 12'b100010010110;
   11284: result <= 12'b100010010110;
   11285: result <= 12'b100010010110;
   11286: result <= 12'b100010010101;
   11287: result <= 12'b100010010101;
   11288: result <= 12'b100010010101;
   11289: result <= 12'b100010010100;
   11290: result <= 12'b100010010100;
   11291: result <= 12'b100010010100;
   11292: result <= 12'b100010010100;
   11293: result <= 12'b100010010011;
   11294: result <= 12'b100010010011;
   11295: result <= 12'b100010010011;
   11296: result <= 12'b100010010010;
   11297: result <= 12'b100010010010;
   11298: result <= 12'b100010010010;
   11299: result <= 12'b100010010010;
   11300: result <= 12'b100010010001;
   11301: result <= 12'b100010010001;
   11302: result <= 12'b100010010001;
   11303: result <= 12'b100010010000;
   11304: result <= 12'b100010010000;
   11305: result <= 12'b100010010000;
   11306: result <= 12'b100010010000;
   11307: result <= 12'b100010001111;
   11308: result <= 12'b100010001111;
   11309: result <= 12'b100010001111;
   11310: result <= 12'b100010001110;
   11311: result <= 12'b100010001110;
   11312: result <= 12'b100010001110;
   11313: result <= 12'b100010001110;
   11314: result <= 12'b100010001101;
   11315: result <= 12'b100010001101;
   11316: result <= 12'b100010001101;
   11317: result <= 12'b100010001100;
   11318: result <= 12'b100010001100;
   11319: result <= 12'b100010001100;
   11320: result <= 12'b100010001100;
   11321: result <= 12'b100010001011;
   11322: result <= 12'b100010001011;
   11323: result <= 12'b100010001011;
   11324: result <= 12'b100010001010;
   11325: result <= 12'b100010001010;
   11326: result <= 12'b100010001010;
   11327: result <= 12'b100010001010;
   11328: result <= 12'b100010001001;
   11329: result <= 12'b100010001001;
   11330: result <= 12'b100010001001;
   11331: result <= 12'b100010001000;
   11332: result <= 12'b100010001000;
   11333: result <= 12'b100010001000;
   11334: result <= 12'b100010001000;
   11335: result <= 12'b100010000111;
   11336: result <= 12'b100010000111;
   11337: result <= 12'b100010000111;
   11338: result <= 12'b100010000110;
   11339: result <= 12'b100010000110;
   11340: result <= 12'b100010000110;
   11341: result <= 12'b100010000110;
   11342: result <= 12'b100010000101;
   11343: result <= 12'b100010000101;
   11344: result <= 12'b100010000101;
   11345: result <= 12'b100010000100;
   11346: result <= 12'b100010000100;
   11347: result <= 12'b100010000100;
   11348: result <= 12'b100010000100;
   11349: result <= 12'b100010000011;
   11350: result <= 12'b100010000011;
   11351: result <= 12'b100010000011;
   11352: result <= 12'b100010000011;
   11353: result <= 12'b100010000010;
   11354: result <= 12'b100010000010;
   11355: result <= 12'b100010000010;
   11356: result <= 12'b100010000001;
   11357: result <= 12'b100010000001;
   11358: result <= 12'b100010000001;
   11359: result <= 12'b100010000001;
   11360: result <= 12'b100010000000;
   11361: result <= 12'b100010000000;
   11362: result <= 12'b100010000000;
   11363: result <= 12'b100010000000;
   11364: result <= 12'b100001111111;
   11365: result <= 12'b100001111111;
   11366: result <= 12'b100001111111;
   11367: result <= 12'b100001111110;
   11368: result <= 12'b100001111110;
   11369: result <= 12'b100001111110;
   11370: result <= 12'b100001111110;
   11371: result <= 12'b100001111101;
   11372: result <= 12'b100001111101;
   11373: result <= 12'b100001111101;
   11374: result <= 12'b100001111101;
   11375: result <= 12'b100001111100;
   11376: result <= 12'b100001111100;
   11377: result <= 12'b100001111100;
   11378: result <= 12'b100001111011;
   11379: result <= 12'b100001111011;
   11380: result <= 12'b100001111011;
   11381: result <= 12'b100001111011;
   11382: result <= 12'b100001111010;
   11383: result <= 12'b100001111010;
   11384: result <= 12'b100001111010;
   11385: result <= 12'b100001111010;
   11386: result <= 12'b100001111001;
   11387: result <= 12'b100001111001;
   11388: result <= 12'b100001111001;
   11389: result <= 12'b100001111001;
   11390: result <= 12'b100001111000;
   11391: result <= 12'b100001111000;
   11392: result <= 12'b100001111000;
   11393: result <= 12'b100001110111;
   11394: result <= 12'b100001110111;
   11395: result <= 12'b100001110111;
   11396: result <= 12'b100001110111;
   11397: result <= 12'b100001110110;
   11398: result <= 12'b100001110110;
   11399: result <= 12'b100001110110;
   11400: result <= 12'b100001110110;
   11401: result <= 12'b100001110101;
   11402: result <= 12'b100001110101;
   11403: result <= 12'b100001110101;
   11404: result <= 12'b100001110101;
   11405: result <= 12'b100001110100;
   11406: result <= 12'b100001110100;
   11407: result <= 12'b100001110100;
   11408: result <= 12'b100001110100;
   11409: result <= 12'b100001110011;
   11410: result <= 12'b100001110011;
   11411: result <= 12'b100001110011;
   11412: result <= 12'b100001110010;
   11413: result <= 12'b100001110010;
   11414: result <= 12'b100001110010;
   11415: result <= 12'b100001110010;
   11416: result <= 12'b100001110001;
   11417: result <= 12'b100001110001;
   11418: result <= 12'b100001110001;
   11419: result <= 12'b100001110001;
   11420: result <= 12'b100001110000;
   11421: result <= 12'b100001110000;
   11422: result <= 12'b100001110000;
   11423: result <= 12'b100001110000;
   11424: result <= 12'b100001101111;
   11425: result <= 12'b100001101111;
   11426: result <= 12'b100001101111;
   11427: result <= 12'b100001101111;
   11428: result <= 12'b100001101110;
   11429: result <= 12'b100001101110;
   11430: result <= 12'b100001101110;
   11431: result <= 12'b100001101110;
   11432: result <= 12'b100001101101;
   11433: result <= 12'b100001101101;
   11434: result <= 12'b100001101101;
   11435: result <= 12'b100001101101;
   11436: result <= 12'b100001101100;
   11437: result <= 12'b100001101100;
   11438: result <= 12'b100001101100;
   11439: result <= 12'b100001101100;
   11440: result <= 12'b100001101011;
   11441: result <= 12'b100001101011;
   11442: result <= 12'b100001101011;
   11443: result <= 12'b100001101011;
   11444: result <= 12'b100001101010;
   11445: result <= 12'b100001101010;
   11446: result <= 12'b100001101010;
   11447: result <= 12'b100001101010;
   11448: result <= 12'b100001101001;
   11449: result <= 12'b100001101001;
   11450: result <= 12'b100001101001;
   11451: result <= 12'b100001101001;
   11452: result <= 12'b100001101000;
   11453: result <= 12'b100001101000;
   11454: result <= 12'b100001101000;
   11455: result <= 12'b100001101000;
   11456: result <= 12'b100001100111;
   11457: result <= 12'b100001100111;
   11458: result <= 12'b100001100111;
   11459: result <= 12'b100001100111;
   11460: result <= 12'b100001100110;
   11461: result <= 12'b100001100110;
   11462: result <= 12'b100001100110;
   11463: result <= 12'b100001100110;
   11464: result <= 12'b100001100101;
   11465: result <= 12'b100001100101;
   11466: result <= 12'b100001100101;
   11467: result <= 12'b100001100101;
   11468: result <= 12'b100001100100;
   11469: result <= 12'b100001100100;
   11470: result <= 12'b100001100100;
   11471: result <= 12'b100001100100;
   11472: result <= 12'b100001100011;
   11473: result <= 12'b100001100011;
   11474: result <= 12'b100001100011;
   11475: result <= 12'b100001100011;
   11476: result <= 12'b100001100010;
   11477: result <= 12'b100001100010;
   11478: result <= 12'b100001100010;
   11479: result <= 12'b100001100010;
   11480: result <= 12'b100001100010;
   11481: result <= 12'b100001100001;
   11482: result <= 12'b100001100001;
   11483: result <= 12'b100001100001;
   11484: result <= 12'b100001100001;
   11485: result <= 12'b100001100000;
   11486: result <= 12'b100001100000;
   11487: result <= 12'b100001100000;
   11488: result <= 12'b100001100000;
   11489: result <= 12'b100001011111;
   11490: result <= 12'b100001011111;
   11491: result <= 12'b100001011111;
   11492: result <= 12'b100001011111;
   11493: result <= 12'b100001011110;
   11494: result <= 12'b100001011110;
   11495: result <= 12'b100001011110;
   11496: result <= 12'b100001011110;
   11497: result <= 12'b100001011110;
   11498: result <= 12'b100001011101;
   11499: result <= 12'b100001011101;
   11500: result <= 12'b100001011101;
   11501: result <= 12'b100001011101;
   11502: result <= 12'b100001011100;
   11503: result <= 12'b100001011100;
   11504: result <= 12'b100001011100;
   11505: result <= 12'b100001011100;
   11506: result <= 12'b100001011011;
   11507: result <= 12'b100001011011;
   11508: result <= 12'b100001011011;
   11509: result <= 12'b100001011011;
   11510: result <= 12'b100001011010;
   11511: result <= 12'b100001011010;
   11512: result <= 12'b100001011010;
   11513: result <= 12'b100001011010;
   11514: result <= 12'b100001011010;
   11515: result <= 12'b100001011001;
   11516: result <= 12'b100001011001;
   11517: result <= 12'b100001011001;
   11518: result <= 12'b100001011001;
   11519: result <= 12'b100001011000;
   11520: result <= 12'b100001011000;
   11521: result <= 12'b100001011000;
   11522: result <= 12'b100001011000;
   11523: result <= 12'b100001011000;
   11524: result <= 12'b100001010111;
   11525: result <= 12'b100001010111;
   11526: result <= 12'b100001010111;
   11527: result <= 12'b100001010111;
   11528: result <= 12'b100001010110;
   11529: result <= 12'b100001010110;
   11530: result <= 12'b100001010110;
   11531: result <= 12'b100001010110;
   11532: result <= 12'b100001010101;
   11533: result <= 12'b100001010101;
   11534: result <= 12'b100001010101;
   11535: result <= 12'b100001010101;
   11536: result <= 12'b100001010101;
   11537: result <= 12'b100001010100;
   11538: result <= 12'b100001010100;
   11539: result <= 12'b100001010100;
   11540: result <= 12'b100001010100;
   11541: result <= 12'b100001010011;
   11542: result <= 12'b100001010011;
   11543: result <= 12'b100001010011;
   11544: result <= 12'b100001010011;
   11545: result <= 12'b100001010011;
   11546: result <= 12'b100001010010;
   11547: result <= 12'b100001010010;
   11548: result <= 12'b100001010010;
   11549: result <= 12'b100001010010;
   11550: result <= 12'b100001010001;
   11551: result <= 12'b100001010001;
   11552: result <= 12'b100001010001;
   11553: result <= 12'b100001010001;
   11554: result <= 12'b100001010001;
   11555: result <= 12'b100001010000;
   11556: result <= 12'b100001010000;
   11557: result <= 12'b100001010000;
   11558: result <= 12'b100001010000;
   11559: result <= 12'b100001010000;
   11560: result <= 12'b100001001111;
   11561: result <= 12'b100001001111;
   11562: result <= 12'b100001001111;
   11563: result <= 12'b100001001111;
   11564: result <= 12'b100001001110;
   11565: result <= 12'b100001001110;
   11566: result <= 12'b100001001110;
   11567: result <= 12'b100001001110;
   11568: result <= 12'b100001001110;
   11569: result <= 12'b100001001101;
   11570: result <= 12'b100001001101;
   11571: result <= 12'b100001001101;
   11572: result <= 12'b100001001101;
   11573: result <= 12'b100001001101;
   11574: result <= 12'b100001001100;
   11575: result <= 12'b100001001100;
   11576: result <= 12'b100001001100;
   11577: result <= 12'b100001001100;
   11578: result <= 12'b100001001011;
   11579: result <= 12'b100001001011;
   11580: result <= 12'b100001001011;
   11581: result <= 12'b100001001011;
   11582: result <= 12'b100001001011;
   11583: result <= 12'b100001001010;
   11584: result <= 12'b100001001010;
   11585: result <= 12'b100001001010;
   11586: result <= 12'b100001001010;
   11587: result <= 12'b100001001010;
   11588: result <= 12'b100001001001;
   11589: result <= 12'b100001001001;
   11590: result <= 12'b100001001001;
   11591: result <= 12'b100001001001;
   11592: result <= 12'b100001001001;
   11593: result <= 12'b100001001000;
   11594: result <= 12'b100001001000;
   11595: result <= 12'b100001001000;
   11596: result <= 12'b100001001000;
   11597: result <= 12'b100001000111;
   11598: result <= 12'b100001000111;
   11599: result <= 12'b100001000111;
   11600: result <= 12'b100001000111;
   11601: result <= 12'b100001000111;
   11602: result <= 12'b100001000110;
   11603: result <= 12'b100001000110;
   11604: result <= 12'b100001000110;
   11605: result <= 12'b100001000110;
   11606: result <= 12'b100001000110;
   11607: result <= 12'b100001000101;
   11608: result <= 12'b100001000101;
   11609: result <= 12'b100001000101;
   11610: result <= 12'b100001000101;
   11611: result <= 12'b100001000101;
   11612: result <= 12'b100001000100;
   11613: result <= 12'b100001000100;
   11614: result <= 12'b100001000100;
   11615: result <= 12'b100001000100;
   11616: result <= 12'b100001000100;
   11617: result <= 12'b100001000011;
   11618: result <= 12'b100001000011;
   11619: result <= 12'b100001000011;
   11620: result <= 12'b100001000011;
   11621: result <= 12'b100001000011;
   11622: result <= 12'b100001000010;
   11623: result <= 12'b100001000010;
   11624: result <= 12'b100001000010;
   11625: result <= 12'b100001000010;
   11626: result <= 12'b100001000010;
   11627: result <= 12'b100001000001;
   11628: result <= 12'b100001000001;
   11629: result <= 12'b100001000001;
   11630: result <= 12'b100001000001;
   11631: result <= 12'b100001000001;
   11632: result <= 12'b100001000000;
   11633: result <= 12'b100001000000;
   11634: result <= 12'b100001000000;
   11635: result <= 12'b100001000000;
   11636: result <= 12'b100001000000;
   11637: result <= 12'b100000111111;
   11638: result <= 12'b100000111111;
   11639: result <= 12'b100000111111;
   11640: result <= 12'b100000111111;
   11641: result <= 12'b100000111111;
   11642: result <= 12'b100000111111;
   11643: result <= 12'b100000111110;
   11644: result <= 12'b100000111110;
   11645: result <= 12'b100000111110;
   11646: result <= 12'b100000111110;
   11647: result <= 12'b100000111110;
   11648: result <= 12'b100000111101;
   11649: result <= 12'b100000111101;
   11650: result <= 12'b100000111101;
   11651: result <= 12'b100000111101;
   11652: result <= 12'b100000111101;
   11653: result <= 12'b100000111100;
   11654: result <= 12'b100000111100;
   11655: result <= 12'b100000111100;
   11656: result <= 12'b100000111100;
   11657: result <= 12'b100000111100;
   11658: result <= 12'b100000111011;
   11659: result <= 12'b100000111011;
   11660: result <= 12'b100000111011;
   11661: result <= 12'b100000111011;
   11662: result <= 12'b100000111011;
   11663: result <= 12'b100000111011;
   11664: result <= 12'b100000111010;
   11665: result <= 12'b100000111010;
   11666: result <= 12'b100000111010;
   11667: result <= 12'b100000111010;
   11668: result <= 12'b100000111010;
   11669: result <= 12'b100000111001;
   11670: result <= 12'b100000111001;
   11671: result <= 12'b100000111001;
   11672: result <= 12'b100000111001;
   11673: result <= 12'b100000111001;
   11674: result <= 12'b100000111001;
   11675: result <= 12'b100000111000;
   11676: result <= 12'b100000111000;
   11677: result <= 12'b100000111000;
   11678: result <= 12'b100000111000;
   11679: result <= 12'b100000111000;
   11680: result <= 12'b100000110111;
   11681: result <= 12'b100000110111;
   11682: result <= 12'b100000110111;
   11683: result <= 12'b100000110111;
   11684: result <= 12'b100000110111;
   11685: result <= 12'b100000110111;
   11686: result <= 12'b100000110110;
   11687: result <= 12'b100000110110;
   11688: result <= 12'b100000110110;
   11689: result <= 12'b100000110110;
   11690: result <= 12'b100000110110;
   11691: result <= 12'b100000110101;
   11692: result <= 12'b100000110101;
   11693: result <= 12'b100000110101;
   11694: result <= 12'b100000110101;
   11695: result <= 12'b100000110101;
   11696: result <= 12'b100000110101;
   11697: result <= 12'b100000110100;
   11698: result <= 12'b100000110100;
   11699: result <= 12'b100000110100;
   11700: result <= 12'b100000110100;
   11701: result <= 12'b100000110100;
   11702: result <= 12'b100000110011;
   11703: result <= 12'b100000110011;
   11704: result <= 12'b100000110011;
   11705: result <= 12'b100000110011;
   11706: result <= 12'b100000110011;
   11707: result <= 12'b100000110011;
   11708: result <= 12'b100000110010;
   11709: result <= 12'b100000110010;
   11710: result <= 12'b100000110010;
   11711: result <= 12'b100000110010;
   11712: result <= 12'b100000110010;
   11713: result <= 12'b100000110010;
   11714: result <= 12'b100000110001;
   11715: result <= 12'b100000110001;
   11716: result <= 12'b100000110001;
   11717: result <= 12'b100000110001;
   11718: result <= 12'b100000110001;
   11719: result <= 12'b100000110001;
   11720: result <= 12'b100000110000;
   11721: result <= 12'b100000110000;
   11722: result <= 12'b100000110000;
   11723: result <= 12'b100000110000;
   11724: result <= 12'b100000110000;
   11725: result <= 12'b100000110000;
   11726: result <= 12'b100000101111;
   11727: result <= 12'b100000101111;
   11728: result <= 12'b100000101111;
   11729: result <= 12'b100000101111;
   11730: result <= 12'b100000101111;
   11731: result <= 12'b100000101111;
   11732: result <= 12'b100000101110;
   11733: result <= 12'b100000101110;
   11734: result <= 12'b100000101110;
   11735: result <= 12'b100000101110;
   11736: result <= 12'b100000101110;
   11737: result <= 12'b100000101110;
   11738: result <= 12'b100000101101;
   11739: result <= 12'b100000101101;
   11740: result <= 12'b100000101101;
   11741: result <= 12'b100000101101;
   11742: result <= 12'b100000101101;
   11743: result <= 12'b100000101101;
   11744: result <= 12'b100000101100;
   11745: result <= 12'b100000101100;
   11746: result <= 12'b100000101100;
   11747: result <= 12'b100000101100;
   11748: result <= 12'b100000101100;
   11749: result <= 12'b100000101100;
   11750: result <= 12'b100000101011;
   11751: result <= 12'b100000101011;
   11752: result <= 12'b100000101011;
   11753: result <= 12'b100000101011;
   11754: result <= 12'b100000101011;
   11755: result <= 12'b100000101011;
   11756: result <= 12'b100000101010;
   11757: result <= 12'b100000101010;
   11758: result <= 12'b100000101010;
   11759: result <= 12'b100000101010;
   11760: result <= 12'b100000101010;
   11761: result <= 12'b100000101010;
   11762: result <= 12'b100000101010;
   11763: result <= 12'b100000101001;
   11764: result <= 12'b100000101001;
   11765: result <= 12'b100000101001;
   11766: result <= 12'b100000101001;
   11767: result <= 12'b100000101001;
   11768: result <= 12'b100000101001;
   11769: result <= 12'b100000101000;
   11770: result <= 12'b100000101000;
   11771: result <= 12'b100000101000;
   11772: result <= 12'b100000101000;
   11773: result <= 12'b100000101000;
   11774: result <= 12'b100000101000;
   11775: result <= 12'b100000101000;
   11776: result <= 12'b100000100111;
   11777: result <= 12'b100000100111;
   11778: result <= 12'b100000100111;
   11779: result <= 12'b100000100111;
   11780: result <= 12'b100000100111;
   11781: result <= 12'b100000100111;
   11782: result <= 12'b100000100110;
   11783: result <= 12'b100000100110;
   11784: result <= 12'b100000100110;
   11785: result <= 12'b100000100110;
   11786: result <= 12'b100000100110;
   11787: result <= 12'b100000100110;
   11788: result <= 12'b100000100110;
   11789: result <= 12'b100000100101;
   11790: result <= 12'b100000100101;
   11791: result <= 12'b100000100101;
   11792: result <= 12'b100000100101;
   11793: result <= 12'b100000100101;
   11794: result <= 12'b100000100101;
   11795: result <= 12'b100000100100;
   11796: result <= 12'b100000100100;
   11797: result <= 12'b100000100100;
   11798: result <= 12'b100000100100;
   11799: result <= 12'b100000100100;
   11800: result <= 12'b100000100100;
   11801: result <= 12'b100000100100;
   11802: result <= 12'b100000100011;
   11803: result <= 12'b100000100011;
   11804: result <= 12'b100000100011;
   11805: result <= 12'b100000100011;
   11806: result <= 12'b100000100011;
   11807: result <= 12'b100000100011;
   11808: result <= 12'b100000100011;
   11809: result <= 12'b100000100010;
   11810: result <= 12'b100000100010;
   11811: result <= 12'b100000100010;
   11812: result <= 12'b100000100010;
   11813: result <= 12'b100000100010;
   11814: result <= 12'b100000100010;
   11815: result <= 12'b100000100010;
   11816: result <= 12'b100000100001;
   11817: result <= 12'b100000100001;
   11818: result <= 12'b100000100001;
   11819: result <= 12'b100000100001;
   11820: result <= 12'b100000100001;
   11821: result <= 12'b100000100001;
   11822: result <= 12'b100000100001;
   11823: result <= 12'b100000100000;
   11824: result <= 12'b100000100000;
   11825: result <= 12'b100000100000;
   11826: result <= 12'b100000100000;
   11827: result <= 12'b100000100000;
   11828: result <= 12'b100000100000;
   11829: result <= 12'b100000100000;
   11830: result <= 12'b100000100000;
   11831: result <= 12'b100000011111;
   11832: result <= 12'b100000011111;
   11833: result <= 12'b100000011111;
   11834: result <= 12'b100000011111;
   11835: result <= 12'b100000011111;
   11836: result <= 12'b100000011111;
   11837: result <= 12'b100000011111;
   11838: result <= 12'b100000011110;
   11839: result <= 12'b100000011110;
   11840: result <= 12'b100000011110;
   11841: result <= 12'b100000011110;
   11842: result <= 12'b100000011110;
   11843: result <= 12'b100000011110;
   11844: result <= 12'b100000011110;
   11845: result <= 12'b100000011101;
   11846: result <= 12'b100000011101;
   11847: result <= 12'b100000011101;
   11848: result <= 12'b100000011101;
   11849: result <= 12'b100000011101;
   11850: result <= 12'b100000011101;
   11851: result <= 12'b100000011101;
   11852: result <= 12'b100000011101;
   11853: result <= 12'b100000011100;
   11854: result <= 12'b100000011100;
   11855: result <= 12'b100000011100;
   11856: result <= 12'b100000011100;
   11857: result <= 12'b100000011100;
   11858: result <= 12'b100000011100;
   11859: result <= 12'b100000011100;
   11860: result <= 12'b100000011100;
   11861: result <= 12'b100000011011;
   11862: result <= 12'b100000011011;
   11863: result <= 12'b100000011011;
   11864: result <= 12'b100000011011;
   11865: result <= 12'b100000011011;
   11866: result <= 12'b100000011011;
   11867: result <= 12'b100000011011;
   11868: result <= 12'b100000011011;
   11869: result <= 12'b100000011010;
   11870: result <= 12'b100000011010;
   11871: result <= 12'b100000011010;
   11872: result <= 12'b100000011010;
   11873: result <= 12'b100000011010;
   11874: result <= 12'b100000011010;
   11875: result <= 12'b100000011010;
   11876: result <= 12'b100000011010;
   11877: result <= 12'b100000011001;
   11878: result <= 12'b100000011001;
   11879: result <= 12'b100000011001;
   11880: result <= 12'b100000011001;
   11881: result <= 12'b100000011001;
   11882: result <= 12'b100000011001;
   11883: result <= 12'b100000011001;
   11884: result <= 12'b100000011001;
   11885: result <= 12'b100000011000;
   11886: result <= 12'b100000011000;
   11887: result <= 12'b100000011000;
   11888: result <= 12'b100000011000;
   11889: result <= 12'b100000011000;
   11890: result <= 12'b100000011000;
   11891: result <= 12'b100000011000;
   11892: result <= 12'b100000011000;
   11893: result <= 12'b100000010111;
   11894: result <= 12'b100000010111;
   11895: result <= 12'b100000010111;
   11896: result <= 12'b100000010111;
   11897: result <= 12'b100000010111;
   11898: result <= 12'b100000010111;
   11899: result <= 12'b100000010111;
   11900: result <= 12'b100000010111;
   11901: result <= 12'b100000010111;
   11902: result <= 12'b100000010110;
   11903: result <= 12'b100000010110;
   11904: result <= 12'b100000010110;
   11905: result <= 12'b100000010110;
   11906: result <= 12'b100000010110;
   11907: result <= 12'b100000010110;
   11908: result <= 12'b100000010110;
   11909: result <= 12'b100000010110;
   11910: result <= 12'b100000010101;
   11911: result <= 12'b100000010101;
   11912: result <= 12'b100000010101;
   11913: result <= 12'b100000010101;
   11914: result <= 12'b100000010101;
   11915: result <= 12'b100000010101;
   11916: result <= 12'b100000010101;
   11917: result <= 12'b100000010101;
   11918: result <= 12'b100000010101;
   11919: result <= 12'b100000010100;
   11920: result <= 12'b100000010100;
   11921: result <= 12'b100000010100;
   11922: result <= 12'b100000010100;
   11923: result <= 12'b100000010100;
   11924: result <= 12'b100000010100;
   11925: result <= 12'b100000010100;
   11926: result <= 12'b100000010100;
   11927: result <= 12'b100000010100;
   11928: result <= 12'b100000010011;
   11929: result <= 12'b100000010011;
   11930: result <= 12'b100000010011;
   11931: result <= 12'b100000010011;
   11932: result <= 12'b100000010011;
   11933: result <= 12'b100000010011;
   11934: result <= 12'b100000010011;
   11935: result <= 12'b100000010011;
   11936: result <= 12'b100000010011;
   11937: result <= 12'b100000010011;
   11938: result <= 12'b100000010010;
   11939: result <= 12'b100000010010;
   11940: result <= 12'b100000010010;
   11941: result <= 12'b100000010010;
   11942: result <= 12'b100000010010;
   11943: result <= 12'b100000010010;
   11944: result <= 12'b100000010010;
   11945: result <= 12'b100000010010;
   11946: result <= 12'b100000010010;
   11947: result <= 12'b100000010001;
   11948: result <= 12'b100000010001;
   11949: result <= 12'b100000010001;
   11950: result <= 12'b100000010001;
   11951: result <= 12'b100000010001;
   11952: result <= 12'b100000010001;
   11953: result <= 12'b100000010001;
   11954: result <= 12'b100000010001;
   11955: result <= 12'b100000010001;
   11956: result <= 12'b100000010001;
   11957: result <= 12'b100000010000;
   11958: result <= 12'b100000010000;
   11959: result <= 12'b100000010000;
   11960: result <= 12'b100000010000;
   11961: result <= 12'b100000010000;
   11962: result <= 12'b100000010000;
   11963: result <= 12'b100000010000;
   11964: result <= 12'b100000010000;
   11965: result <= 12'b100000010000;
   11966: result <= 12'b100000010000;
   11967: result <= 12'b100000001111;
   11968: result <= 12'b100000001111;
   11969: result <= 12'b100000001111;
   11970: result <= 12'b100000001111;
   11971: result <= 12'b100000001111;
   11972: result <= 12'b100000001111;
   11973: result <= 12'b100000001111;
   11974: result <= 12'b100000001111;
   11975: result <= 12'b100000001111;
   11976: result <= 12'b100000001111;
   11977: result <= 12'b100000001111;
   11978: result <= 12'b100000001110;
   11979: result <= 12'b100000001110;
   11980: result <= 12'b100000001110;
   11981: result <= 12'b100000001110;
   11982: result <= 12'b100000001110;
   11983: result <= 12'b100000001110;
   11984: result <= 12'b100000001110;
   11985: result <= 12'b100000001110;
   11986: result <= 12'b100000001110;
   11987: result <= 12'b100000001110;
   11988: result <= 12'b100000001110;
   11989: result <= 12'b100000001101;
   11990: result <= 12'b100000001101;
   11991: result <= 12'b100000001101;
   11992: result <= 12'b100000001101;
   11993: result <= 12'b100000001101;
   11994: result <= 12'b100000001101;
   11995: result <= 12'b100000001101;
   11996: result <= 12'b100000001101;
   11997: result <= 12'b100000001101;
   11998: result <= 12'b100000001101;
   11999: result <= 12'b100000001101;
   12000: result <= 12'b100000001100;
   12001: result <= 12'b100000001100;
   12002: result <= 12'b100000001100;
   12003: result <= 12'b100000001100;
   12004: result <= 12'b100000001100;
   12005: result <= 12'b100000001100;
   12006: result <= 12'b100000001100;
   12007: result <= 12'b100000001100;
   12008: result <= 12'b100000001100;
   12009: result <= 12'b100000001100;
   12010: result <= 12'b100000001100;
   12011: result <= 12'b100000001100;
   12012: result <= 12'b100000001011;
   12013: result <= 12'b100000001011;
   12014: result <= 12'b100000001011;
   12015: result <= 12'b100000001011;
   12016: result <= 12'b100000001011;
   12017: result <= 12'b100000001011;
   12018: result <= 12'b100000001011;
   12019: result <= 12'b100000001011;
   12020: result <= 12'b100000001011;
   12021: result <= 12'b100000001011;
   12022: result <= 12'b100000001011;
   12023: result <= 12'b100000001011;
   12024: result <= 12'b100000001010;
   12025: result <= 12'b100000001010;
   12026: result <= 12'b100000001010;
   12027: result <= 12'b100000001010;
   12028: result <= 12'b100000001010;
   12029: result <= 12'b100000001010;
   12030: result <= 12'b100000001010;
   12031: result <= 12'b100000001010;
   12032: result <= 12'b100000001010;
   12033: result <= 12'b100000001010;
   12034: result <= 12'b100000001010;
   12035: result <= 12'b100000001010;
   12036: result <= 12'b100000001010;
   12037: result <= 12'b100000001001;
   12038: result <= 12'b100000001001;
   12039: result <= 12'b100000001001;
   12040: result <= 12'b100000001001;
   12041: result <= 12'b100000001001;
   12042: result <= 12'b100000001001;
   12043: result <= 12'b100000001001;
   12044: result <= 12'b100000001001;
   12045: result <= 12'b100000001001;
   12046: result <= 12'b100000001001;
   12047: result <= 12'b100000001001;
   12048: result <= 12'b100000001001;
   12049: result <= 12'b100000001001;
   12050: result <= 12'b100000001001;
   12051: result <= 12'b100000001000;
   12052: result <= 12'b100000001000;
   12053: result <= 12'b100000001000;
   12054: result <= 12'b100000001000;
   12055: result <= 12'b100000001000;
   12056: result <= 12'b100000001000;
   12057: result <= 12'b100000001000;
   12058: result <= 12'b100000001000;
   12059: result <= 12'b100000001000;
   12060: result <= 12'b100000001000;
   12061: result <= 12'b100000001000;
   12062: result <= 12'b100000001000;
   12063: result <= 12'b100000001000;
   12064: result <= 12'b100000001000;
   12065: result <= 12'b100000000111;
   12066: result <= 12'b100000000111;
   12067: result <= 12'b100000000111;
   12068: result <= 12'b100000000111;
   12069: result <= 12'b100000000111;
   12070: result <= 12'b100000000111;
   12071: result <= 12'b100000000111;
   12072: result <= 12'b100000000111;
   12073: result <= 12'b100000000111;
   12074: result <= 12'b100000000111;
   12075: result <= 12'b100000000111;
   12076: result <= 12'b100000000111;
   12077: result <= 12'b100000000111;
   12078: result <= 12'b100000000111;
   12079: result <= 12'b100000000111;
   12080: result <= 12'b100000000111;
   12081: result <= 12'b100000000110;
   12082: result <= 12'b100000000110;
   12083: result <= 12'b100000000110;
   12084: result <= 12'b100000000110;
   12085: result <= 12'b100000000110;
   12086: result <= 12'b100000000110;
   12087: result <= 12'b100000000110;
   12088: result <= 12'b100000000110;
   12089: result <= 12'b100000000110;
   12090: result <= 12'b100000000110;
   12091: result <= 12'b100000000110;
   12092: result <= 12'b100000000110;
   12093: result <= 12'b100000000110;
   12094: result <= 12'b100000000110;
   12095: result <= 12'b100000000110;
   12096: result <= 12'b100000000110;
   12097: result <= 12'b100000000101;
   12098: result <= 12'b100000000101;
   12099: result <= 12'b100000000101;
   12100: result <= 12'b100000000101;
   12101: result <= 12'b100000000101;
   12102: result <= 12'b100000000101;
   12103: result <= 12'b100000000101;
   12104: result <= 12'b100000000101;
   12105: result <= 12'b100000000101;
   12106: result <= 12'b100000000101;
   12107: result <= 12'b100000000101;
   12108: result <= 12'b100000000101;
   12109: result <= 12'b100000000101;
   12110: result <= 12'b100000000101;
   12111: result <= 12'b100000000101;
   12112: result <= 12'b100000000101;
   12113: result <= 12'b100000000101;
   12114: result <= 12'b100000000101;
   12115: result <= 12'b100000000101;
   12116: result <= 12'b100000000100;
   12117: result <= 12'b100000000100;
   12118: result <= 12'b100000000100;
   12119: result <= 12'b100000000100;
   12120: result <= 12'b100000000100;
   12121: result <= 12'b100000000100;
   12122: result <= 12'b100000000100;
   12123: result <= 12'b100000000100;
   12124: result <= 12'b100000000100;
   12125: result <= 12'b100000000100;
   12126: result <= 12'b100000000100;
   12127: result <= 12'b100000000100;
   12128: result <= 12'b100000000100;
   12129: result <= 12'b100000000100;
   12130: result <= 12'b100000000100;
   12131: result <= 12'b100000000100;
   12132: result <= 12'b100000000100;
   12133: result <= 12'b100000000100;
   12134: result <= 12'b100000000100;
   12135: result <= 12'b100000000100;
   12136: result <= 12'b100000000011;
   12137: result <= 12'b100000000011;
   12138: result <= 12'b100000000011;
   12139: result <= 12'b100000000011;
   12140: result <= 12'b100000000011;
   12141: result <= 12'b100000000011;
   12142: result <= 12'b100000000011;
   12143: result <= 12'b100000000011;
   12144: result <= 12'b100000000011;
   12145: result <= 12'b100000000011;
   12146: result <= 12'b100000000011;
   12147: result <= 12'b100000000011;
   12148: result <= 12'b100000000011;
   12149: result <= 12'b100000000011;
   12150: result <= 12'b100000000011;
   12151: result <= 12'b100000000011;
   12152: result <= 12'b100000000011;
   12153: result <= 12'b100000000011;
   12154: result <= 12'b100000000011;
   12155: result <= 12'b100000000011;
   12156: result <= 12'b100000000011;
   12157: result <= 12'b100000000011;
   12158: result <= 12'b100000000011;
   12159: result <= 12'b100000000011;
   12160: result <= 12'b100000000010;
   12161: result <= 12'b100000000010;
   12162: result <= 12'b100000000010;
   12163: result <= 12'b100000000010;
   12164: result <= 12'b100000000010;
   12165: result <= 12'b100000000010;
   12166: result <= 12'b100000000010;
   12167: result <= 12'b100000000010;
   12168: result <= 12'b100000000010;
   12169: result <= 12'b100000000010;
   12170: result <= 12'b100000000010;
   12171: result <= 12'b100000000010;
   12172: result <= 12'b100000000010;
   12173: result <= 12'b100000000010;
   12174: result <= 12'b100000000010;
   12175: result <= 12'b100000000010;
   12176: result <= 12'b100000000010;
   12177: result <= 12'b100000000010;
   12178: result <= 12'b100000000010;
   12179: result <= 12'b100000000010;
   12180: result <= 12'b100000000010;
   12181: result <= 12'b100000000010;
   12182: result <= 12'b100000000010;
   12183: result <= 12'b100000000010;
   12184: result <= 12'b100000000010;
   12185: result <= 12'b100000000010;
   12186: result <= 12'b100000000010;
   12187: result <= 12'b100000000010;
   12188: result <= 12'b100000000010;
   12189: result <= 12'b100000000001;
   12190: result <= 12'b100000000001;
   12191: result <= 12'b100000000001;
   12192: result <= 12'b100000000001;
   12193: result <= 12'b100000000001;
   12194: result <= 12'b100000000001;
   12195: result <= 12'b100000000001;
   12196: result <= 12'b100000000001;
   12197: result <= 12'b100000000001;
   12198: result <= 12'b100000000001;
   12199: result <= 12'b100000000001;
   12200: result <= 12'b100000000001;
   12201: result <= 12'b100000000001;
   12202: result <= 12'b100000000001;
   12203: result <= 12'b100000000001;
   12204: result <= 12'b100000000001;
   12205: result <= 12'b100000000001;
   12206: result <= 12'b100000000001;
   12207: result <= 12'b100000000001;
   12208: result <= 12'b100000000001;
   12209: result <= 12'b100000000001;
   12210: result <= 12'b100000000001;
   12211: result <= 12'b100000000001;
   12212: result <= 12'b100000000001;
   12213: result <= 12'b100000000001;
   12214: result <= 12'b100000000001;
   12215: result <= 12'b100000000001;
   12216: result <= 12'b100000000001;
   12217: result <= 12'b100000000001;
   12218: result <= 12'b100000000001;
   12219: result <= 12'b100000000001;
   12220: result <= 12'b100000000001;
   12221: result <= 12'b100000000001;
   12222: result <= 12'b100000000001;
   12223: result <= 12'b100000000001;
   12224: result <= 12'b100000000001;
   12225: result <= 12'b100000000001;
   12226: result <= 12'b100000000001;
   12227: result <= 12'b100000000001;
   12228: result <= 12'b100000000001;
   12229: result <= 12'b100000000001;
   12230: result <= 12'b100000000001;
   12231: result <= 12'b100000000000;
   12232: result <= 12'b100000000000;
   12233: result <= 12'b100000000000;
   12234: result <= 12'b100000000000;
   12235: result <= 12'b100000000000;
   12236: result <= 12'b100000000000;
   12237: result <= 12'b100000000000;
   12238: result <= 12'b100000000000;
   12239: result <= 12'b100000000000;
   12240: result <= 12'b100000000000;
   12241: result <= 12'b100000000000;
   12242: result <= 12'b100000000000;
   12243: result <= 12'b100000000000;
   12244: result <= 12'b100000000000;
   12245: result <= 12'b100000000000;
   12246: result <= 12'b100000000000;
   12247: result <= 12'b100000000000;
   12248: result <= 12'b100000000000;
   12249: result <= 12'b100000000000;
   12250: result <= 12'b100000000000;
   12251: result <= 12'b100000000000;
   12252: result <= 12'b100000000000;
   12253: result <= 12'b100000000000;
   12254: result <= 12'b100000000000;
   12255: result <= 12'b100000000000;
   12256: result <= 12'b100000000000;
   12257: result <= 12'b100000000000;
   12258: result <= 12'b100000000000;
   12259: result <= 12'b100000000000;
   12260: result <= 12'b100000000000;
   12261: result <= 12'b100000000000;
   12262: result <= 12'b100000000000;
   12263: result <= 12'b100000000000;
   12264: result <= 12'b100000000000;
   12265: result <= 12'b100000000000;
   12266: result <= 12'b100000000000;
   12267: result <= 12'b100000000000;
   12268: result <= 12'b100000000000;
   12269: result <= 12'b100000000000;
   12270: result <= 12'b100000000000;
   12271: result <= 12'b100000000000;
   12272: result <= 12'b100000000000;
   12273: result <= 12'b100000000000;
   12274: result <= 12'b100000000000;
   12275: result <= 12'b100000000000;
   12276: result <= 12'b100000000000;
   12277: result <= 12'b100000000000;
   12278: result <= 12'b100000000000;
   12279: result <= 12'b100000000000;
   12280: result <= 12'b100000000000;
   12281: result <= 12'b100000000000;
   12282: result <= 12'b100000000000;
   12283: result <= 12'b100000000000;
   12284: result <= 12'b100000000000;
   12285: result <= 12'b100000000000;
   12286: result <= 12'b100000000000;
   12287: result <= 12'b100000000000;
   12288: result <= 12'b100000000000;
   12289: result <= 12'b100000000000;
   12290: result <= 12'b100000000000;
   12291: result <= 12'b100000000000;
   12292: result <= 12'b100000000000;
   12293: result <= 12'b100000000000;
   12294: result <= 12'b100000000000;
   12295: result <= 12'b100000000000;
   12296: result <= 12'b100000000000;
   12297: result <= 12'b100000000000;
   12298: result <= 12'b100000000000;
   12299: result <= 12'b100000000000;
   12300: result <= 12'b100000000000;
   12301: result <= 12'b100000000000;
   12302: result <= 12'b100000000000;
   12303: result <= 12'b100000000000;
   12304: result <= 12'b100000000000;
   12305: result <= 12'b100000000000;
   12306: result <= 12'b100000000000;
   12307: result <= 12'b100000000000;
   12308: result <= 12'b100000000000;
   12309: result <= 12'b100000000000;
   12310: result <= 12'b100000000000;
   12311: result <= 12'b100000000000;
   12312: result <= 12'b100000000000;
   12313: result <= 12'b100000000000;
   12314: result <= 12'b100000000000;
   12315: result <= 12'b100000000000;
   12316: result <= 12'b100000000000;
   12317: result <= 12'b100000000000;
   12318: result <= 12'b100000000000;
   12319: result <= 12'b100000000000;
   12320: result <= 12'b100000000000;
   12321: result <= 12'b100000000000;
   12322: result <= 12'b100000000000;
   12323: result <= 12'b100000000000;
   12324: result <= 12'b100000000000;
   12325: result <= 12'b100000000000;
   12326: result <= 12'b100000000000;
   12327: result <= 12'b100000000000;
   12328: result <= 12'b100000000000;
   12329: result <= 12'b100000000000;
   12330: result <= 12'b100000000000;
   12331: result <= 12'b100000000000;
   12332: result <= 12'b100000000000;
   12333: result <= 12'b100000000000;
   12334: result <= 12'b100000000000;
   12335: result <= 12'b100000000000;
   12336: result <= 12'b100000000000;
   12337: result <= 12'b100000000000;
   12338: result <= 12'b100000000000;
   12339: result <= 12'b100000000000;
   12340: result <= 12'b100000000000;
   12341: result <= 12'b100000000000;
   12342: result <= 12'b100000000000;
   12343: result <= 12'b100000000000;
   12344: result <= 12'b100000000000;
   12345: result <= 12'b100000000000;
   12346: result <= 12'b100000000001;
   12347: result <= 12'b100000000001;
   12348: result <= 12'b100000000001;
   12349: result <= 12'b100000000001;
   12350: result <= 12'b100000000001;
   12351: result <= 12'b100000000001;
   12352: result <= 12'b100000000001;
   12353: result <= 12'b100000000001;
   12354: result <= 12'b100000000001;
   12355: result <= 12'b100000000001;
   12356: result <= 12'b100000000001;
   12357: result <= 12'b100000000001;
   12358: result <= 12'b100000000001;
   12359: result <= 12'b100000000001;
   12360: result <= 12'b100000000001;
   12361: result <= 12'b100000000001;
   12362: result <= 12'b100000000001;
   12363: result <= 12'b100000000001;
   12364: result <= 12'b100000000001;
   12365: result <= 12'b100000000001;
   12366: result <= 12'b100000000001;
   12367: result <= 12'b100000000001;
   12368: result <= 12'b100000000001;
   12369: result <= 12'b100000000001;
   12370: result <= 12'b100000000001;
   12371: result <= 12'b100000000001;
   12372: result <= 12'b100000000001;
   12373: result <= 12'b100000000001;
   12374: result <= 12'b100000000001;
   12375: result <= 12'b100000000001;
   12376: result <= 12'b100000000001;
   12377: result <= 12'b100000000001;
   12378: result <= 12'b100000000001;
   12379: result <= 12'b100000000001;
   12380: result <= 12'b100000000001;
   12381: result <= 12'b100000000001;
   12382: result <= 12'b100000000001;
   12383: result <= 12'b100000000001;
   12384: result <= 12'b100000000001;
   12385: result <= 12'b100000000001;
   12386: result <= 12'b100000000001;
   12387: result <= 12'b100000000001;
   12388: result <= 12'b100000000010;
   12389: result <= 12'b100000000010;
   12390: result <= 12'b100000000010;
   12391: result <= 12'b100000000010;
   12392: result <= 12'b100000000010;
   12393: result <= 12'b100000000010;
   12394: result <= 12'b100000000010;
   12395: result <= 12'b100000000010;
   12396: result <= 12'b100000000010;
   12397: result <= 12'b100000000010;
   12398: result <= 12'b100000000010;
   12399: result <= 12'b100000000010;
   12400: result <= 12'b100000000010;
   12401: result <= 12'b100000000010;
   12402: result <= 12'b100000000010;
   12403: result <= 12'b100000000010;
   12404: result <= 12'b100000000010;
   12405: result <= 12'b100000000010;
   12406: result <= 12'b100000000010;
   12407: result <= 12'b100000000010;
   12408: result <= 12'b100000000010;
   12409: result <= 12'b100000000010;
   12410: result <= 12'b100000000010;
   12411: result <= 12'b100000000010;
   12412: result <= 12'b100000000010;
   12413: result <= 12'b100000000010;
   12414: result <= 12'b100000000010;
   12415: result <= 12'b100000000010;
   12416: result <= 12'b100000000010;
   12417: result <= 12'b100000000011;
   12418: result <= 12'b100000000011;
   12419: result <= 12'b100000000011;
   12420: result <= 12'b100000000011;
   12421: result <= 12'b100000000011;
   12422: result <= 12'b100000000011;
   12423: result <= 12'b100000000011;
   12424: result <= 12'b100000000011;
   12425: result <= 12'b100000000011;
   12426: result <= 12'b100000000011;
   12427: result <= 12'b100000000011;
   12428: result <= 12'b100000000011;
   12429: result <= 12'b100000000011;
   12430: result <= 12'b100000000011;
   12431: result <= 12'b100000000011;
   12432: result <= 12'b100000000011;
   12433: result <= 12'b100000000011;
   12434: result <= 12'b100000000011;
   12435: result <= 12'b100000000011;
   12436: result <= 12'b100000000011;
   12437: result <= 12'b100000000011;
   12438: result <= 12'b100000000011;
   12439: result <= 12'b100000000011;
   12440: result <= 12'b100000000011;
   12441: result <= 12'b100000000100;
   12442: result <= 12'b100000000100;
   12443: result <= 12'b100000000100;
   12444: result <= 12'b100000000100;
   12445: result <= 12'b100000000100;
   12446: result <= 12'b100000000100;
   12447: result <= 12'b100000000100;
   12448: result <= 12'b100000000100;
   12449: result <= 12'b100000000100;
   12450: result <= 12'b100000000100;
   12451: result <= 12'b100000000100;
   12452: result <= 12'b100000000100;
   12453: result <= 12'b100000000100;
   12454: result <= 12'b100000000100;
   12455: result <= 12'b100000000100;
   12456: result <= 12'b100000000100;
   12457: result <= 12'b100000000100;
   12458: result <= 12'b100000000100;
   12459: result <= 12'b100000000100;
   12460: result <= 12'b100000000100;
   12461: result <= 12'b100000000101;
   12462: result <= 12'b100000000101;
   12463: result <= 12'b100000000101;
   12464: result <= 12'b100000000101;
   12465: result <= 12'b100000000101;
   12466: result <= 12'b100000000101;
   12467: result <= 12'b100000000101;
   12468: result <= 12'b100000000101;
   12469: result <= 12'b100000000101;
   12470: result <= 12'b100000000101;
   12471: result <= 12'b100000000101;
   12472: result <= 12'b100000000101;
   12473: result <= 12'b100000000101;
   12474: result <= 12'b100000000101;
   12475: result <= 12'b100000000101;
   12476: result <= 12'b100000000101;
   12477: result <= 12'b100000000101;
   12478: result <= 12'b100000000101;
   12479: result <= 12'b100000000101;
   12480: result <= 12'b100000000110;
   12481: result <= 12'b100000000110;
   12482: result <= 12'b100000000110;
   12483: result <= 12'b100000000110;
   12484: result <= 12'b100000000110;
   12485: result <= 12'b100000000110;
   12486: result <= 12'b100000000110;
   12487: result <= 12'b100000000110;
   12488: result <= 12'b100000000110;
   12489: result <= 12'b100000000110;
   12490: result <= 12'b100000000110;
   12491: result <= 12'b100000000110;
   12492: result <= 12'b100000000110;
   12493: result <= 12'b100000000110;
   12494: result <= 12'b100000000110;
   12495: result <= 12'b100000000110;
   12496: result <= 12'b100000000111;
   12497: result <= 12'b100000000111;
   12498: result <= 12'b100000000111;
   12499: result <= 12'b100000000111;
   12500: result <= 12'b100000000111;
   12501: result <= 12'b100000000111;
   12502: result <= 12'b100000000111;
   12503: result <= 12'b100000000111;
   12504: result <= 12'b100000000111;
   12505: result <= 12'b100000000111;
   12506: result <= 12'b100000000111;
   12507: result <= 12'b100000000111;
   12508: result <= 12'b100000000111;
   12509: result <= 12'b100000000111;
   12510: result <= 12'b100000000111;
   12511: result <= 12'b100000000111;
   12512: result <= 12'b100000001000;
   12513: result <= 12'b100000001000;
   12514: result <= 12'b100000001000;
   12515: result <= 12'b100000001000;
   12516: result <= 12'b100000001000;
   12517: result <= 12'b100000001000;
   12518: result <= 12'b100000001000;
   12519: result <= 12'b100000001000;
   12520: result <= 12'b100000001000;
   12521: result <= 12'b100000001000;
   12522: result <= 12'b100000001000;
   12523: result <= 12'b100000001000;
   12524: result <= 12'b100000001000;
   12525: result <= 12'b100000001000;
   12526: result <= 12'b100000001001;
   12527: result <= 12'b100000001001;
   12528: result <= 12'b100000001001;
   12529: result <= 12'b100000001001;
   12530: result <= 12'b100000001001;
   12531: result <= 12'b100000001001;
   12532: result <= 12'b100000001001;
   12533: result <= 12'b100000001001;
   12534: result <= 12'b100000001001;
   12535: result <= 12'b100000001001;
   12536: result <= 12'b100000001001;
   12537: result <= 12'b100000001001;
   12538: result <= 12'b100000001001;
   12539: result <= 12'b100000001001;
   12540: result <= 12'b100000001010;
   12541: result <= 12'b100000001010;
   12542: result <= 12'b100000001010;
   12543: result <= 12'b100000001010;
   12544: result <= 12'b100000001010;
   12545: result <= 12'b100000001010;
   12546: result <= 12'b100000001010;
   12547: result <= 12'b100000001010;
   12548: result <= 12'b100000001010;
   12549: result <= 12'b100000001010;
   12550: result <= 12'b100000001010;
   12551: result <= 12'b100000001010;
   12552: result <= 12'b100000001010;
   12553: result <= 12'b100000001011;
   12554: result <= 12'b100000001011;
   12555: result <= 12'b100000001011;
   12556: result <= 12'b100000001011;
   12557: result <= 12'b100000001011;
   12558: result <= 12'b100000001011;
   12559: result <= 12'b100000001011;
   12560: result <= 12'b100000001011;
   12561: result <= 12'b100000001011;
   12562: result <= 12'b100000001011;
   12563: result <= 12'b100000001011;
   12564: result <= 12'b100000001011;
   12565: result <= 12'b100000001100;
   12566: result <= 12'b100000001100;
   12567: result <= 12'b100000001100;
   12568: result <= 12'b100000001100;
   12569: result <= 12'b100000001100;
   12570: result <= 12'b100000001100;
   12571: result <= 12'b100000001100;
   12572: result <= 12'b100000001100;
   12573: result <= 12'b100000001100;
   12574: result <= 12'b100000001100;
   12575: result <= 12'b100000001100;
   12576: result <= 12'b100000001100;
   12577: result <= 12'b100000001101;
   12578: result <= 12'b100000001101;
   12579: result <= 12'b100000001101;
   12580: result <= 12'b100000001101;
   12581: result <= 12'b100000001101;
   12582: result <= 12'b100000001101;
   12583: result <= 12'b100000001101;
   12584: result <= 12'b100000001101;
   12585: result <= 12'b100000001101;
   12586: result <= 12'b100000001101;
   12587: result <= 12'b100000001101;
   12588: result <= 12'b100000001110;
   12589: result <= 12'b100000001110;
   12590: result <= 12'b100000001110;
   12591: result <= 12'b100000001110;
   12592: result <= 12'b100000001110;
   12593: result <= 12'b100000001110;
   12594: result <= 12'b100000001110;
   12595: result <= 12'b100000001110;
   12596: result <= 12'b100000001110;
   12597: result <= 12'b100000001110;
   12598: result <= 12'b100000001110;
   12599: result <= 12'b100000001111;
   12600: result <= 12'b100000001111;
   12601: result <= 12'b100000001111;
   12602: result <= 12'b100000001111;
   12603: result <= 12'b100000001111;
   12604: result <= 12'b100000001111;
   12605: result <= 12'b100000001111;
   12606: result <= 12'b100000001111;
   12607: result <= 12'b100000001111;
   12608: result <= 12'b100000001111;
   12609: result <= 12'b100000001111;
   12610: result <= 12'b100000010000;
   12611: result <= 12'b100000010000;
   12612: result <= 12'b100000010000;
   12613: result <= 12'b100000010000;
   12614: result <= 12'b100000010000;
   12615: result <= 12'b100000010000;
   12616: result <= 12'b100000010000;
   12617: result <= 12'b100000010000;
   12618: result <= 12'b100000010000;
   12619: result <= 12'b100000010000;
   12620: result <= 12'b100000010001;
   12621: result <= 12'b100000010001;
   12622: result <= 12'b100000010001;
   12623: result <= 12'b100000010001;
   12624: result <= 12'b100000010001;
   12625: result <= 12'b100000010001;
   12626: result <= 12'b100000010001;
   12627: result <= 12'b100000010001;
   12628: result <= 12'b100000010001;
   12629: result <= 12'b100000010001;
   12630: result <= 12'b100000010010;
   12631: result <= 12'b100000010010;
   12632: result <= 12'b100000010010;
   12633: result <= 12'b100000010010;
   12634: result <= 12'b100000010010;
   12635: result <= 12'b100000010010;
   12636: result <= 12'b100000010010;
   12637: result <= 12'b100000010010;
   12638: result <= 12'b100000010010;
   12639: result <= 12'b100000010011;
   12640: result <= 12'b100000010011;
   12641: result <= 12'b100000010011;
   12642: result <= 12'b100000010011;
   12643: result <= 12'b100000010011;
   12644: result <= 12'b100000010011;
   12645: result <= 12'b100000010011;
   12646: result <= 12'b100000010011;
   12647: result <= 12'b100000010011;
   12648: result <= 12'b100000010011;
   12649: result <= 12'b100000010100;
   12650: result <= 12'b100000010100;
   12651: result <= 12'b100000010100;
   12652: result <= 12'b100000010100;
   12653: result <= 12'b100000010100;
   12654: result <= 12'b100000010100;
   12655: result <= 12'b100000010100;
   12656: result <= 12'b100000010100;
   12657: result <= 12'b100000010100;
   12658: result <= 12'b100000010101;
   12659: result <= 12'b100000010101;
   12660: result <= 12'b100000010101;
   12661: result <= 12'b100000010101;
   12662: result <= 12'b100000010101;
   12663: result <= 12'b100000010101;
   12664: result <= 12'b100000010101;
   12665: result <= 12'b100000010101;
   12666: result <= 12'b100000010101;
   12667: result <= 12'b100000010110;
   12668: result <= 12'b100000010110;
   12669: result <= 12'b100000010110;
   12670: result <= 12'b100000010110;
   12671: result <= 12'b100000010110;
   12672: result <= 12'b100000010110;
   12673: result <= 12'b100000010110;
   12674: result <= 12'b100000010110;
   12675: result <= 12'b100000010111;
   12676: result <= 12'b100000010111;
   12677: result <= 12'b100000010111;
   12678: result <= 12'b100000010111;
   12679: result <= 12'b100000010111;
   12680: result <= 12'b100000010111;
   12681: result <= 12'b100000010111;
   12682: result <= 12'b100000010111;
   12683: result <= 12'b100000010111;
   12684: result <= 12'b100000011000;
   12685: result <= 12'b100000011000;
   12686: result <= 12'b100000011000;
   12687: result <= 12'b100000011000;
   12688: result <= 12'b100000011000;
   12689: result <= 12'b100000011000;
   12690: result <= 12'b100000011000;
   12691: result <= 12'b100000011000;
   12692: result <= 12'b100000011001;
   12693: result <= 12'b100000011001;
   12694: result <= 12'b100000011001;
   12695: result <= 12'b100000011001;
   12696: result <= 12'b100000011001;
   12697: result <= 12'b100000011001;
   12698: result <= 12'b100000011001;
   12699: result <= 12'b100000011001;
   12700: result <= 12'b100000011010;
   12701: result <= 12'b100000011010;
   12702: result <= 12'b100000011010;
   12703: result <= 12'b100000011010;
   12704: result <= 12'b100000011010;
   12705: result <= 12'b100000011010;
   12706: result <= 12'b100000011010;
   12707: result <= 12'b100000011010;
   12708: result <= 12'b100000011011;
   12709: result <= 12'b100000011011;
   12710: result <= 12'b100000011011;
   12711: result <= 12'b100000011011;
   12712: result <= 12'b100000011011;
   12713: result <= 12'b100000011011;
   12714: result <= 12'b100000011011;
   12715: result <= 12'b100000011011;
   12716: result <= 12'b100000011100;
   12717: result <= 12'b100000011100;
   12718: result <= 12'b100000011100;
   12719: result <= 12'b100000011100;
   12720: result <= 12'b100000011100;
   12721: result <= 12'b100000011100;
   12722: result <= 12'b100000011100;
   12723: result <= 12'b100000011100;
   12724: result <= 12'b100000011101;
   12725: result <= 12'b100000011101;
   12726: result <= 12'b100000011101;
   12727: result <= 12'b100000011101;
   12728: result <= 12'b100000011101;
   12729: result <= 12'b100000011101;
   12730: result <= 12'b100000011101;
   12731: result <= 12'b100000011101;
   12732: result <= 12'b100000011110;
   12733: result <= 12'b100000011110;
   12734: result <= 12'b100000011110;
   12735: result <= 12'b100000011110;
   12736: result <= 12'b100000011110;
   12737: result <= 12'b100000011110;
   12738: result <= 12'b100000011110;
   12739: result <= 12'b100000011111;
   12740: result <= 12'b100000011111;
   12741: result <= 12'b100000011111;
   12742: result <= 12'b100000011111;
   12743: result <= 12'b100000011111;
   12744: result <= 12'b100000011111;
   12745: result <= 12'b100000011111;
   12746: result <= 12'b100000100000;
   12747: result <= 12'b100000100000;
   12748: result <= 12'b100000100000;
   12749: result <= 12'b100000100000;
   12750: result <= 12'b100000100000;
   12751: result <= 12'b100000100000;
   12752: result <= 12'b100000100000;
   12753: result <= 12'b100000100000;
   12754: result <= 12'b100000100001;
   12755: result <= 12'b100000100001;
   12756: result <= 12'b100000100001;
   12757: result <= 12'b100000100001;
   12758: result <= 12'b100000100001;
   12759: result <= 12'b100000100001;
   12760: result <= 12'b100000100001;
   12761: result <= 12'b100000100010;
   12762: result <= 12'b100000100010;
   12763: result <= 12'b100000100010;
   12764: result <= 12'b100000100010;
   12765: result <= 12'b100000100010;
   12766: result <= 12'b100000100010;
   12767: result <= 12'b100000100010;
   12768: result <= 12'b100000100011;
   12769: result <= 12'b100000100011;
   12770: result <= 12'b100000100011;
   12771: result <= 12'b100000100011;
   12772: result <= 12'b100000100011;
   12773: result <= 12'b100000100011;
   12774: result <= 12'b100000100011;
   12775: result <= 12'b100000100100;
   12776: result <= 12'b100000100100;
   12777: result <= 12'b100000100100;
   12778: result <= 12'b100000100100;
   12779: result <= 12'b100000100100;
   12780: result <= 12'b100000100100;
   12781: result <= 12'b100000100100;
   12782: result <= 12'b100000100101;
   12783: result <= 12'b100000100101;
   12784: result <= 12'b100000100101;
   12785: result <= 12'b100000100101;
   12786: result <= 12'b100000100101;
   12787: result <= 12'b100000100101;
   12788: result <= 12'b100000100110;
   12789: result <= 12'b100000100110;
   12790: result <= 12'b100000100110;
   12791: result <= 12'b100000100110;
   12792: result <= 12'b100000100110;
   12793: result <= 12'b100000100110;
   12794: result <= 12'b100000100110;
   12795: result <= 12'b100000100111;
   12796: result <= 12'b100000100111;
   12797: result <= 12'b100000100111;
   12798: result <= 12'b100000100111;
   12799: result <= 12'b100000100111;
   12800: result <= 12'b100000100111;
   12801: result <= 12'b100000101000;
   12802: result <= 12'b100000101000;
   12803: result <= 12'b100000101000;
   12804: result <= 12'b100000101000;
   12805: result <= 12'b100000101000;
   12806: result <= 12'b100000101000;
   12807: result <= 12'b100000101000;
   12808: result <= 12'b100000101001;
   12809: result <= 12'b100000101001;
   12810: result <= 12'b100000101001;
   12811: result <= 12'b100000101001;
   12812: result <= 12'b100000101001;
   12813: result <= 12'b100000101001;
   12814: result <= 12'b100000101010;
   12815: result <= 12'b100000101010;
   12816: result <= 12'b100000101010;
   12817: result <= 12'b100000101010;
   12818: result <= 12'b100000101010;
   12819: result <= 12'b100000101010;
   12820: result <= 12'b100000101010;
   12821: result <= 12'b100000101011;
   12822: result <= 12'b100000101011;
   12823: result <= 12'b100000101011;
   12824: result <= 12'b100000101011;
   12825: result <= 12'b100000101011;
   12826: result <= 12'b100000101011;
   12827: result <= 12'b100000101100;
   12828: result <= 12'b100000101100;
   12829: result <= 12'b100000101100;
   12830: result <= 12'b100000101100;
   12831: result <= 12'b100000101100;
   12832: result <= 12'b100000101100;
   12833: result <= 12'b100000101101;
   12834: result <= 12'b100000101101;
   12835: result <= 12'b100000101101;
   12836: result <= 12'b100000101101;
   12837: result <= 12'b100000101101;
   12838: result <= 12'b100000101101;
   12839: result <= 12'b100000101110;
   12840: result <= 12'b100000101110;
   12841: result <= 12'b100000101110;
   12842: result <= 12'b100000101110;
   12843: result <= 12'b100000101110;
   12844: result <= 12'b100000101110;
   12845: result <= 12'b100000101111;
   12846: result <= 12'b100000101111;
   12847: result <= 12'b100000101111;
   12848: result <= 12'b100000101111;
   12849: result <= 12'b100000101111;
   12850: result <= 12'b100000101111;
   12851: result <= 12'b100000110000;
   12852: result <= 12'b100000110000;
   12853: result <= 12'b100000110000;
   12854: result <= 12'b100000110000;
   12855: result <= 12'b100000110000;
   12856: result <= 12'b100000110000;
   12857: result <= 12'b100000110001;
   12858: result <= 12'b100000110001;
   12859: result <= 12'b100000110001;
   12860: result <= 12'b100000110001;
   12861: result <= 12'b100000110001;
   12862: result <= 12'b100000110001;
   12863: result <= 12'b100000110010;
   12864: result <= 12'b100000110010;
   12865: result <= 12'b100000110010;
   12866: result <= 12'b100000110010;
   12867: result <= 12'b100000110010;
   12868: result <= 12'b100000110010;
   12869: result <= 12'b100000110011;
   12870: result <= 12'b100000110011;
   12871: result <= 12'b100000110011;
   12872: result <= 12'b100000110011;
   12873: result <= 12'b100000110011;
   12874: result <= 12'b100000110011;
   12875: result <= 12'b100000110100;
   12876: result <= 12'b100000110100;
   12877: result <= 12'b100000110100;
   12878: result <= 12'b100000110100;
   12879: result <= 12'b100000110100;
   12880: result <= 12'b100000110101;
   12881: result <= 12'b100000110101;
   12882: result <= 12'b100000110101;
   12883: result <= 12'b100000110101;
   12884: result <= 12'b100000110101;
   12885: result <= 12'b100000110101;
   12886: result <= 12'b100000110110;
   12887: result <= 12'b100000110110;
   12888: result <= 12'b100000110110;
   12889: result <= 12'b100000110110;
   12890: result <= 12'b100000110110;
   12891: result <= 12'b100000110111;
   12892: result <= 12'b100000110111;
   12893: result <= 12'b100000110111;
   12894: result <= 12'b100000110111;
   12895: result <= 12'b100000110111;
   12896: result <= 12'b100000110111;
   12897: result <= 12'b100000111000;
   12898: result <= 12'b100000111000;
   12899: result <= 12'b100000111000;
   12900: result <= 12'b100000111000;
   12901: result <= 12'b100000111000;
   12902: result <= 12'b100000111001;
   12903: result <= 12'b100000111001;
   12904: result <= 12'b100000111001;
   12905: result <= 12'b100000111001;
   12906: result <= 12'b100000111001;
   12907: result <= 12'b100000111001;
   12908: result <= 12'b100000111010;
   12909: result <= 12'b100000111010;
   12910: result <= 12'b100000111010;
   12911: result <= 12'b100000111010;
   12912: result <= 12'b100000111010;
   12913: result <= 12'b100000111011;
   12914: result <= 12'b100000111011;
   12915: result <= 12'b100000111011;
   12916: result <= 12'b100000111011;
   12917: result <= 12'b100000111011;
   12918: result <= 12'b100000111011;
   12919: result <= 12'b100000111100;
   12920: result <= 12'b100000111100;
   12921: result <= 12'b100000111100;
   12922: result <= 12'b100000111100;
   12923: result <= 12'b100000111100;
   12924: result <= 12'b100000111101;
   12925: result <= 12'b100000111101;
   12926: result <= 12'b100000111101;
   12927: result <= 12'b100000111101;
   12928: result <= 12'b100000111101;
   12929: result <= 12'b100000111110;
   12930: result <= 12'b100000111110;
   12931: result <= 12'b100000111110;
   12932: result <= 12'b100000111110;
   12933: result <= 12'b100000111110;
   12934: result <= 12'b100000111111;
   12935: result <= 12'b100000111111;
   12936: result <= 12'b100000111111;
   12937: result <= 12'b100000111111;
   12938: result <= 12'b100000111111;
   12939: result <= 12'b100000111111;
   12940: result <= 12'b100001000000;
   12941: result <= 12'b100001000000;
   12942: result <= 12'b100001000000;
   12943: result <= 12'b100001000000;
   12944: result <= 12'b100001000000;
   12945: result <= 12'b100001000001;
   12946: result <= 12'b100001000001;
   12947: result <= 12'b100001000001;
   12948: result <= 12'b100001000001;
   12949: result <= 12'b100001000001;
   12950: result <= 12'b100001000010;
   12951: result <= 12'b100001000010;
   12952: result <= 12'b100001000010;
   12953: result <= 12'b100001000010;
   12954: result <= 12'b100001000010;
   12955: result <= 12'b100001000011;
   12956: result <= 12'b100001000011;
   12957: result <= 12'b100001000011;
   12958: result <= 12'b100001000011;
   12959: result <= 12'b100001000011;
   12960: result <= 12'b100001000100;
   12961: result <= 12'b100001000100;
   12962: result <= 12'b100001000100;
   12963: result <= 12'b100001000100;
   12964: result <= 12'b100001000100;
   12965: result <= 12'b100001000101;
   12966: result <= 12'b100001000101;
   12967: result <= 12'b100001000101;
   12968: result <= 12'b100001000101;
   12969: result <= 12'b100001000101;
   12970: result <= 12'b100001000110;
   12971: result <= 12'b100001000110;
   12972: result <= 12'b100001000110;
   12973: result <= 12'b100001000110;
   12974: result <= 12'b100001000110;
   12975: result <= 12'b100001000111;
   12976: result <= 12'b100001000111;
   12977: result <= 12'b100001000111;
   12978: result <= 12'b100001000111;
   12979: result <= 12'b100001000111;
   12980: result <= 12'b100001001000;
   12981: result <= 12'b100001001000;
   12982: result <= 12'b100001001000;
   12983: result <= 12'b100001001000;
   12984: result <= 12'b100001001001;
   12985: result <= 12'b100001001001;
   12986: result <= 12'b100001001001;
   12987: result <= 12'b100001001001;
   12988: result <= 12'b100001001001;
   12989: result <= 12'b100001001010;
   12990: result <= 12'b100001001010;
   12991: result <= 12'b100001001010;
   12992: result <= 12'b100001001010;
   12993: result <= 12'b100001001010;
   12994: result <= 12'b100001001011;
   12995: result <= 12'b100001001011;
   12996: result <= 12'b100001001011;
   12997: result <= 12'b100001001011;
   12998: result <= 12'b100001001011;
   12999: result <= 12'b100001001100;
   13000: result <= 12'b100001001100;
   13001: result <= 12'b100001001100;
   13002: result <= 12'b100001001100;
   13003: result <= 12'b100001001101;
   13004: result <= 12'b100001001101;
   13005: result <= 12'b100001001101;
   13006: result <= 12'b100001001101;
   13007: result <= 12'b100001001101;
   13008: result <= 12'b100001001110;
   13009: result <= 12'b100001001110;
   13010: result <= 12'b100001001110;
   13011: result <= 12'b100001001110;
   13012: result <= 12'b100001001110;
   13013: result <= 12'b100001001111;
   13014: result <= 12'b100001001111;
   13015: result <= 12'b100001001111;
   13016: result <= 12'b100001001111;
   13017: result <= 12'b100001010000;
   13018: result <= 12'b100001010000;
   13019: result <= 12'b100001010000;
   13020: result <= 12'b100001010000;
   13021: result <= 12'b100001010000;
   13022: result <= 12'b100001010001;
   13023: result <= 12'b100001010001;
   13024: result <= 12'b100001010001;
   13025: result <= 12'b100001010001;
   13026: result <= 12'b100001010001;
   13027: result <= 12'b100001010010;
   13028: result <= 12'b100001010010;
   13029: result <= 12'b100001010010;
   13030: result <= 12'b100001010010;
   13031: result <= 12'b100001010011;
   13032: result <= 12'b100001010011;
   13033: result <= 12'b100001010011;
   13034: result <= 12'b100001010011;
   13035: result <= 12'b100001010011;
   13036: result <= 12'b100001010100;
   13037: result <= 12'b100001010100;
   13038: result <= 12'b100001010100;
   13039: result <= 12'b100001010100;
   13040: result <= 12'b100001010101;
   13041: result <= 12'b100001010101;
   13042: result <= 12'b100001010101;
   13043: result <= 12'b100001010101;
   13044: result <= 12'b100001010101;
   13045: result <= 12'b100001010110;
   13046: result <= 12'b100001010110;
   13047: result <= 12'b100001010110;
   13048: result <= 12'b100001010110;
   13049: result <= 12'b100001010111;
   13050: result <= 12'b100001010111;
   13051: result <= 12'b100001010111;
   13052: result <= 12'b100001010111;
   13053: result <= 12'b100001011000;
   13054: result <= 12'b100001011000;
   13055: result <= 12'b100001011000;
   13056: result <= 12'b100001011000;
   13057: result <= 12'b100001011000;
   13058: result <= 12'b100001011001;
   13059: result <= 12'b100001011001;
   13060: result <= 12'b100001011001;
   13061: result <= 12'b100001011001;
   13062: result <= 12'b100001011010;
   13063: result <= 12'b100001011010;
   13064: result <= 12'b100001011010;
   13065: result <= 12'b100001011010;
   13066: result <= 12'b100001011010;
   13067: result <= 12'b100001011011;
   13068: result <= 12'b100001011011;
   13069: result <= 12'b100001011011;
   13070: result <= 12'b100001011011;
   13071: result <= 12'b100001011100;
   13072: result <= 12'b100001011100;
   13073: result <= 12'b100001011100;
   13074: result <= 12'b100001011100;
   13075: result <= 12'b100001011101;
   13076: result <= 12'b100001011101;
   13077: result <= 12'b100001011101;
   13078: result <= 12'b100001011101;
   13079: result <= 12'b100001011110;
   13080: result <= 12'b100001011110;
   13081: result <= 12'b100001011110;
   13082: result <= 12'b100001011110;
   13083: result <= 12'b100001011110;
   13084: result <= 12'b100001011111;
   13085: result <= 12'b100001011111;
   13086: result <= 12'b100001011111;
   13087: result <= 12'b100001011111;
   13088: result <= 12'b100001100000;
   13089: result <= 12'b100001100000;
   13090: result <= 12'b100001100000;
   13091: result <= 12'b100001100000;
   13092: result <= 12'b100001100001;
   13093: result <= 12'b100001100001;
   13094: result <= 12'b100001100001;
   13095: result <= 12'b100001100001;
   13096: result <= 12'b100001100010;
   13097: result <= 12'b100001100010;
   13098: result <= 12'b100001100010;
   13099: result <= 12'b100001100010;
   13100: result <= 12'b100001100010;
   13101: result <= 12'b100001100011;
   13102: result <= 12'b100001100011;
   13103: result <= 12'b100001100011;
   13104: result <= 12'b100001100011;
   13105: result <= 12'b100001100100;
   13106: result <= 12'b100001100100;
   13107: result <= 12'b100001100100;
   13108: result <= 12'b100001100100;
   13109: result <= 12'b100001100101;
   13110: result <= 12'b100001100101;
   13111: result <= 12'b100001100101;
   13112: result <= 12'b100001100101;
   13113: result <= 12'b100001100110;
   13114: result <= 12'b100001100110;
   13115: result <= 12'b100001100110;
   13116: result <= 12'b100001100110;
   13117: result <= 12'b100001100111;
   13118: result <= 12'b100001100111;
   13119: result <= 12'b100001100111;
   13120: result <= 12'b100001100111;
   13121: result <= 12'b100001101000;
   13122: result <= 12'b100001101000;
   13123: result <= 12'b100001101000;
   13124: result <= 12'b100001101000;
   13125: result <= 12'b100001101001;
   13126: result <= 12'b100001101001;
   13127: result <= 12'b100001101001;
   13128: result <= 12'b100001101001;
   13129: result <= 12'b100001101010;
   13130: result <= 12'b100001101010;
   13131: result <= 12'b100001101010;
   13132: result <= 12'b100001101010;
   13133: result <= 12'b100001101011;
   13134: result <= 12'b100001101011;
   13135: result <= 12'b100001101011;
   13136: result <= 12'b100001101011;
   13137: result <= 12'b100001101100;
   13138: result <= 12'b100001101100;
   13139: result <= 12'b100001101100;
   13140: result <= 12'b100001101100;
   13141: result <= 12'b100001101101;
   13142: result <= 12'b100001101101;
   13143: result <= 12'b100001101101;
   13144: result <= 12'b100001101101;
   13145: result <= 12'b100001101110;
   13146: result <= 12'b100001101110;
   13147: result <= 12'b100001101110;
   13148: result <= 12'b100001101110;
   13149: result <= 12'b100001101111;
   13150: result <= 12'b100001101111;
   13151: result <= 12'b100001101111;
   13152: result <= 12'b100001101111;
   13153: result <= 12'b100001110000;
   13154: result <= 12'b100001110000;
   13155: result <= 12'b100001110000;
   13156: result <= 12'b100001110000;
   13157: result <= 12'b100001110001;
   13158: result <= 12'b100001110001;
   13159: result <= 12'b100001110001;
   13160: result <= 12'b100001110001;
   13161: result <= 12'b100001110010;
   13162: result <= 12'b100001110010;
   13163: result <= 12'b100001110010;
   13164: result <= 12'b100001110010;
   13165: result <= 12'b100001110011;
   13166: result <= 12'b100001110011;
   13167: result <= 12'b100001110011;
   13168: result <= 12'b100001110100;
   13169: result <= 12'b100001110100;
   13170: result <= 12'b100001110100;
   13171: result <= 12'b100001110100;
   13172: result <= 12'b100001110101;
   13173: result <= 12'b100001110101;
   13174: result <= 12'b100001110101;
   13175: result <= 12'b100001110101;
   13176: result <= 12'b100001110110;
   13177: result <= 12'b100001110110;
   13178: result <= 12'b100001110110;
   13179: result <= 12'b100001110110;
   13180: result <= 12'b100001110111;
   13181: result <= 12'b100001110111;
   13182: result <= 12'b100001110111;
   13183: result <= 12'b100001110111;
   13184: result <= 12'b100001111000;
   13185: result <= 12'b100001111000;
   13186: result <= 12'b100001111000;
   13187: result <= 12'b100001111001;
   13188: result <= 12'b100001111001;
   13189: result <= 12'b100001111001;
   13190: result <= 12'b100001111001;
   13191: result <= 12'b100001111010;
   13192: result <= 12'b100001111010;
   13193: result <= 12'b100001111010;
   13194: result <= 12'b100001111010;
   13195: result <= 12'b100001111011;
   13196: result <= 12'b100001111011;
   13197: result <= 12'b100001111011;
   13198: result <= 12'b100001111011;
   13199: result <= 12'b100001111100;
   13200: result <= 12'b100001111100;
   13201: result <= 12'b100001111100;
   13202: result <= 12'b100001111101;
   13203: result <= 12'b100001111101;
   13204: result <= 12'b100001111101;
   13205: result <= 12'b100001111101;
   13206: result <= 12'b100001111110;
   13207: result <= 12'b100001111110;
   13208: result <= 12'b100001111110;
   13209: result <= 12'b100001111110;
   13210: result <= 12'b100001111111;
   13211: result <= 12'b100001111111;
   13212: result <= 12'b100001111111;
   13213: result <= 12'b100010000000;
   13214: result <= 12'b100010000000;
   13215: result <= 12'b100010000000;
   13216: result <= 12'b100010000000;
   13217: result <= 12'b100010000001;
   13218: result <= 12'b100010000001;
   13219: result <= 12'b100010000001;
   13220: result <= 12'b100010000001;
   13221: result <= 12'b100010000010;
   13222: result <= 12'b100010000010;
   13223: result <= 12'b100010000010;
   13224: result <= 12'b100010000011;
   13225: result <= 12'b100010000011;
   13226: result <= 12'b100010000011;
   13227: result <= 12'b100010000011;
   13228: result <= 12'b100010000100;
   13229: result <= 12'b100010000100;
   13230: result <= 12'b100010000100;
   13231: result <= 12'b100010000100;
   13232: result <= 12'b100010000101;
   13233: result <= 12'b100010000101;
   13234: result <= 12'b100010000101;
   13235: result <= 12'b100010000110;
   13236: result <= 12'b100010000110;
   13237: result <= 12'b100010000110;
   13238: result <= 12'b100010000110;
   13239: result <= 12'b100010000111;
   13240: result <= 12'b100010000111;
   13241: result <= 12'b100010000111;
   13242: result <= 12'b100010001000;
   13243: result <= 12'b100010001000;
   13244: result <= 12'b100010001000;
   13245: result <= 12'b100010001000;
   13246: result <= 12'b100010001001;
   13247: result <= 12'b100010001001;
   13248: result <= 12'b100010001001;
   13249: result <= 12'b100010001010;
   13250: result <= 12'b100010001010;
   13251: result <= 12'b100010001010;
   13252: result <= 12'b100010001010;
   13253: result <= 12'b100010001011;
   13254: result <= 12'b100010001011;
   13255: result <= 12'b100010001011;
   13256: result <= 12'b100010001100;
   13257: result <= 12'b100010001100;
   13258: result <= 12'b100010001100;
   13259: result <= 12'b100010001100;
   13260: result <= 12'b100010001101;
   13261: result <= 12'b100010001101;
   13262: result <= 12'b100010001101;
   13263: result <= 12'b100010001110;
   13264: result <= 12'b100010001110;
   13265: result <= 12'b100010001110;
   13266: result <= 12'b100010001110;
   13267: result <= 12'b100010001111;
   13268: result <= 12'b100010001111;
   13269: result <= 12'b100010001111;
   13270: result <= 12'b100010010000;
   13271: result <= 12'b100010010000;
   13272: result <= 12'b100010010000;
   13273: result <= 12'b100010010000;
   13274: result <= 12'b100010010001;
   13275: result <= 12'b100010010001;
   13276: result <= 12'b100010010001;
   13277: result <= 12'b100010010010;
   13278: result <= 12'b100010010010;
   13279: result <= 12'b100010010010;
   13280: result <= 12'b100010010010;
   13281: result <= 12'b100010010011;
   13282: result <= 12'b100010010011;
   13283: result <= 12'b100010010011;
   13284: result <= 12'b100010010100;
   13285: result <= 12'b100010010100;
   13286: result <= 12'b100010010100;
   13287: result <= 12'b100010010100;
   13288: result <= 12'b100010010101;
   13289: result <= 12'b100010010101;
   13290: result <= 12'b100010010101;
   13291: result <= 12'b100010010110;
   13292: result <= 12'b100010010110;
   13293: result <= 12'b100010010110;
   13294: result <= 12'b100010010111;
   13295: result <= 12'b100010010111;
   13296: result <= 12'b100010010111;
   13297: result <= 12'b100010010111;
   13298: result <= 12'b100010011000;
   13299: result <= 12'b100010011000;
   13300: result <= 12'b100010011000;
   13301: result <= 12'b100010011001;
   13302: result <= 12'b100010011001;
   13303: result <= 12'b100010011001;
   13304: result <= 12'b100010011001;
   13305: result <= 12'b100010011010;
   13306: result <= 12'b100010011010;
   13307: result <= 12'b100010011010;
   13308: result <= 12'b100010011011;
   13309: result <= 12'b100010011011;
   13310: result <= 12'b100010011011;
   13311: result <= 12'b100010011100;
   13312: result <= 12'b100010011100;
   13313: result <= 12'b100010011100;
   13314: result <= 12'b100010011100;
   13315: result <= 12'b100010011101;
   13316: result <= 12'b100010011101;
   13317: result <= 12'b100010011101;
   13318: result <= 12'b100010011110;
   13319: result <= 12'b100010011110;
   13320: result <= 12'b100010011110;
   13321: result <= 12'b100010011111;
   13322: result <= 12'b100010011111;
   13323: result <= 12'b100010011111;
   13324: result <= 12'b100010100000;
   13325: result <= 12'b100010100000;
   13326: result <= 12'b100010100000;
   13327: result <= 12'b100010100000;
   13328: result <= 12'b100010100001;
   13329: result <= 12'b100010100001;
   13330: result <= 12'b100010100001;
   13331: result <= 12'b100010100010;
   13332: result <= 12'b100010100010;
   13333: result <= 12'b100010100010;
   13334: result <= 12'b100010100011;
   13335: result <= 12'b100010100011;
   13336: result <= 12'b100010100011;
   13337: result <= 12'b100010100011;
   13338: result <= 12'b100010100100;
   13339: result <= 12'b100010100100;
   13340: result <= 12'b100010100100;
   13341: result <= 12'b100010100101;
   13342: result <= 12'b100010100101;
   13343: result <= 12'b100010100101;
   13344: result <= 12'b100010100110;
   13345: result <= 12'b100010100110;
   13346: result <= 12'b100010100110;
   13347: result <= 12'b100010100111;
   13348: result <= 12'b100010100111;
   13349: result <= 12'b100010100111;
   13350: result <= 12'b100010101000;
   13351: result <= 12'b100010101000;
   13352: result <= 12'b100010101000;
   13353: result <= 12'b100010101000;
   13354: result <= 12'b100010101001;
   13355: result <= 12'b100010101001;
   13356: result <= 12'b100010101001;
   13357: result <= 12'b100010101010;
   13358: result <= 12'b100010101010;
   13359: result <= 12'b100010101010;
   13360: result <= 12'b100010101011;
   13361: result <= 12'b100010101011;
   13362: result <= 12'b100010101011;
   13363: result <= 12'b100010101100;
   13364: result <= 12'b100010101100;
   13365: result <= 12'b100010101100;
   13366: result <= 12'b100010101101;
   13367: result <= 12'b100010101101;
   13368: result <= 12'b100010101101;
   13369: result <= 12'b100010101101;
   13370: result <= 12'b100010101110;
   13371: result <= 12'b100010101110;
   13372: result <= 12'b100010101110;
   13373: result <= 12'b100010101111;
   13374: result <= 12'b100010101111;
   13375: result <= 12'b100010101111;
   13376: result <= 12'b100010110000;
   13377: result <= 12'b100010110000;
   13378: result <= 12'b100010110000;
   13379: result <= 12'b100010110001;
   13380: result <= 12'b100010110001;
   13381: result <= 12'b100010110001;
   13382: result <= 12'b100010110010;
   13383: result <= 12'b100010110010;
   13384: result <= 12'b100010110010;
   13385: result <= 12'b100010110011;
   13386: result <= 12'b100010110011;
   13387: result <= 12'b100010110011;
   13388: result <= 12'b100010110100;
   13389: result <= 12'b100010110100;
   13390: result <= 12'b100010110100;
   13391: result <= 12'b100010110101;
   13392: result <= 12'b100010110101;
   13393: result <= 12'b100010110101;
   13394: result <= 12'b100010110101;
   13395: result <= 12'b100010110110;
   13396: result <= 12'b100010110110;
   13397: result <= 12'b100010110110;
   13398: result <= 12'b100010110111;
   13399: result <= 12'b100010110111;
   13400: result <= 12'b100010110111;
   13401: result <= 12'b100010111000;
   13402: result <= 12'b100010111000;
   13403: result <= 12'b100010111000;
   13404: result <= 12'b100010111001;
   13405: result <= 12'b100010111001;
   13406: result <= 12'b100010111001;
   13407: result <= 12'b100010111010;
   13408: result <= 12'b100010111010;
   13409: result <= 12'b100010111010;
   13410: result <= 12'b100010111011;
   13411: result <= 12'b100010111011;
   13412: result <= 12'b100010111011;
   13413: result <= 12'b100010111100;
   13414: result <= 12'b100010111100;
   13415: result <= 12'b100010111100;
   13416: result <= 12'b100010111101;
   13417: result <= 12'b100010111101;
   13418: result <= 12'b100010111101;
   13419: result <= 12'b100010111110;
   13420: result <= 12'b100010111110;
   13421: result <= 12'b100010111110;
   13422: result <= 12'b100010111111;
   13423: result <= 12'b100010111111;
   13424: result <= 12'b100010111111;
   13425: result <= 12'b100011000000;
   13426: result <= 12'b100011000000;
   13427: result <= 12'b100011000000;
   13428: result <= 12'b100011000001;
   13429: result <= 12'b100011000001;
   13430: result <= 12'b100011000001;
   13431: result <= 12'b100011000010;
   13432: result <= 12'b100011000010;
   13433: result <= 12'b100011000010;
   13434: result <= 12'b100011000011;
   13435: result <= 12'b100011000011;
   13436: result <= 12'b100011000011;
   13437: result <= 12'b100011000100;
   13438: result <= 12'b100011000100;
   13439: result <= 12'b100011000100;
   13440: result <= 12'b100011000101;
   13441: result <= 12'b100011000101;
   13442: result <= 12'b100011000101;
   13443: result <= 12'b100011000110;
   13444: result <= 12'b100011000110;
   13445: result <= 12'b100011000110;
   13446: result <= 12'b100011000111;
   13447: result <= 12'b100011000111;
   13448: result <= 12'b100011000111;
   13449: result <= 12'b100011001000;
   13450: result <= 12'b100011001000;
   13451: result <= 12'b100011001000;
   13452: result <= 12'b100011001001;
   13453: result <= 12'b100011001001;
   13454: result <= 12'b100011001001;
   13455: result <= 12'b100011001010;
   13456: result <= 12'b100011001010;
   13457: result <= 12'b100011001010;
   13458: result <= 12'b100011001011;
   13459: result <= 12'b100011001011;
   13460: result <= 12'b100011001011;
   13461: result <= 12'b100011001100;
   13462: result <= 12'b100011001100;
   13463: result <= 12'b100011001100;
   13464: result <= 12'b100011001101;
   13465: result <= 12'b100011001101;
   13466: result <= 12'b100011001101;
   13467: result <= 12'b100011001110;
   13468: result <= 12'b100011001110;
   13469: result <= 12'b100011001110;
   13470: result <= 12'b100011001111;
   13471: result <= 12'b100011001111;
   13472: result <= 12'b100011010000;
   13473: result <= 12'b100011010000;
   13474: result <= 12'b100011010000;
   13475: result <= 12'b100011010001;
   13476: result <= 12'b100011010001;
   13477: result <= 12'b100011010001;
   13478: result <= 12'b100011010010;
   13479: result <= 12'b100011010010;
   13480: result <= 12'b100011010010;
   13481: result <= 12'b100011010011;
   13482: result <= 12'b100011010011;
   13483: result <= 12'b100011010011;
   13484: result <= 12'b100011010100;
   13485: result <= 12'b100011010100;
   13486: result <= 12'b100011010100;
   13487: result <= 12'b100011010101;
   13488: result <= 12'b100011010101;
   13489: result <= 12'b100011010101;
   13490: result <= 12'b100011010110;
   13491: result <= 12'b100011010110;
   13492: result <= 12'b100011010110;
   13493: result <= 12'b100011010111;
   13494: result <= 12'b100011010111;
   13495: result <= 12'b100011011000;
   13496: result <= 12'b100011011000;
   13497: result <= 12'b100011011000;
   13498: result <= 12'b100011011001;
   13499: result <= 12'b100011011001;
   13500: result <= 12'b100011011001;
   13501: result <= 12'b100011011010;
   13502: result <= 12'b100011011010;
   13503: result <= 12'b100011011010;
   13504: result <= 12'b100011011011;
   13505: result <= 12'b100011011011;
   13506: result <= 12'b100011011011;
   13507: result <= 12'b100011011100;
   13508: result <= 12'b100011011100;
   13509: result <= 12'b100011011100;
   13510: result <= 12'b100011011101;
   13511: result <= 12'b100011011101;
   13512: result <= 12'b100011011110;
   13513: result <= 12'b100011011110;
   13514: result <= 12'b100011011110;
   13515: result <= 12'b100011011111;
   13516: result <= 12'b100011011111;
   13517: result <= 12'b100011011111;
   13518: result <= 12'b100011100000;
   13519: result <= 12'b100011100000;
   13520: result <= 12'b100011100000;
   13521: result <= 12'b100011100001;
   13522: result <= 12'b100011100001;
   13523: result <= 12'b100011100001;
   13524: result <= 12'b100011100010;
   13525: result <= 12'b100011100010;
   13526: result <= 12'b100011100011;
   13527: result <= 12'b100011100011;
   13528: result <= 12'b100011100011;
   13529: result <= 12'b100011100100;
   13530: result <= 12'b100011100100;
   13531: result <= 12'b100011100100;
   13532: result <= 12'b100011100101;
   13533: result <= 12'b100011100101;
   13534: result <= 12'b100011100101;
   13535: result <= 12'b100011100110;
   13536: result <= 12'b100011100110;
   13537: result <= 12'b100011100110;
   13538: result <= 12'b100011100111;
   13539: result <= 12'b100011100111;
   13540: result <= 12'b100011101000;
   13541: result <= 12'b100011101000;
   13542: result <= 12'b100011101000;
   13543: result <= 12'b100011101001;
   13544: result <= 12'b100011101001;
   13545: result <= 12'b100011101001;
   13546: result <= 12'b100011101010;
   13547: result <= 12'b100011101010;
   13548: result <= 12'b100011101010;
   13549: result <= 12'b100011101011;
   13550: result <= 12'b100011101011;
   13551: result <= 12'b100011101100;
   13552: result <= 12'b100011101100;
   13553: result <= 12'b100011101100;
   13554: result <= 12'b100011101101;
   13555: result <= 12'b100011101101;
   13556: result <= 12'b100011101101;
   13557: result <= 12'b100011101110;
   13558: result <= 12'b100011101110;
   13559: result <= 12'b100011101111;
   13560: result <= 12'b100011101111;
   13561: result <= 12'b100011101111;
   13562: result <= 12'b100011110000;
   13563: result <= 12'b100011110000;
   13564: result <= 12'b100011110000;
   13565: result <= 12'b100011110001;
   13566: result <= 12'b100011110001;
   13567: result <= 12'b100011110001;
   13568: result <= 12'b100011110010;
   13569: result <= 12'b100011110010;
   13570: result <= 12'b100011110011;
   13571: result <= 12'b100011110011;
   13572: result <= 12'b100011110011;
   13573: result <= 12'b100011110100;
   13574: result <= 12'b100011110100;
   13575: result <= 12'b100011110100;
   13576: result <= 12'b100011110101;
   13577: result <= 12'b100011110101;
   13578: result <= 12'b100011110110;
   13579: result <= 12'b100011110110;
   13580: result <= 12'b100011110110;
   13581: result <= 12'b100011110111;
   13582: result <= 12'b100011110111;
   13583: result <= 12'b100011110111;
   13584: result <= 12'b100011111000;
   13585: result <= 12'b100011111000;
   13586: result <= 12'b100011111001;
   13587: result <= 12'b100011111001;
   13588: result <= 12'b100011111001;
   13589: result <= 12'b100011111010;
   13590: result <= 12'b100011111010;
   13591: result <= 12'b100011111010;
   13592: result <= 12'b100011111011;
   13593: result <= 12'b100011111011;
   13594: result <= 12'b100011111100;
   13595: result <= 12'b100011111100;
   13596: result <= 12'b100011111100;
   13597: result <= 12'b100011111101;
   13598: result <= 12'b100011111101;
   13599: result <= 12'b100011111101;
   13600: result <= 12'b100011111110;
   13601: result <= 12'b100011111110;
   13602: result <= 12'b100011111111;
   13603: result <= 12'b100011111111;
   13604: result <= 12'b100011111111;
   13605: result <= 12'b100100000000;
   13606: result <= 12'b100100000000;
   13607: result <= 12'b100100000000;
   13608: result <= 12'b100100000001;
   13609: result <= 12'b100100000001;
   13610: result <= 12'b100100000010;
   13611: result <= 12'b100100000010;
   13612: result <= 12'b100100000010;
   13613: result <= 12'b100100000011;
   13614: result <= 12'b100100000011;
   13615: result <= 12'b100100000100;
   13616: result <= 12'b100100000100;
   13617: result <= 12'b100100000100;
   13618: result <= 12'b100100000101;
   13619: result <= 12'b100100000101;
   13620: result <= 12'b100100000101;
   13621: result <= 12'b100100000110;
   13622: result <= 12'b100100000110;
   13623: result <= 12'b100100000111;
   13624: result <= 12'b100100000111;
   13625: result <= 12'b100100000111;
   13626: result <= 12'b100100001000;
   13627: result <= 12'b100100001000;
   13628: result <= 12'b100100001001;
   13629: result <= 12'b100100001001;
   13630: result <= 12'b100100001001;
   13631: result <= 12'b100100001010;
   13632: result <= 12'b100100001010;
   13633: result <= 12'b100100001010;
   13634: result <= 12'b100100001011;
   13635: result <= 12'b100100001011;
   13636: result <= 12'b100100001100;
   13637: result <= 12'b100100001100;
   13638: result <= 12'b100100001100;
   13639: result <= 12'b100100001101;
   13640: result <= 12'b100100001101;
   13641: result <= 12'b100100001110;
   13642: result <= 12'b100100001110;
   13643: result <= 12'b100100001110;
   13644: result <= 12'b100100001111;
   13645: result <= 12'b100100001111;
   13646: result <= 12'b100100010000;
   13647: result <= 12'b100100010000;
   13648: result <= 12'b100100010000;
   13649: result <= 12'b100100010001;
   13650: result <= 12'b100100010001;
   13651: result <= 12'b100100010001;
   13652: result <= 12'b100100010010;
   13653: result <= 12'b100100010010;
   13654: result <= 12'b100100010011;
   13655: result <= 12'b100100010011;
   13656: result <= 12'b100100010011;
   13657: result <= 12'b100100010100;
   13658: result <= 12'b100100010100;
   13659: result <= 12'b100100010101;
   13660: result <= 12'b100100010101;
   13661: result <= 12'b100100010101;
   13662: result <= 12'b100100010110;
   13663: result <= 12'b100100010110;
   13664: result <= 12'b100100010111;
   13665: result <= 12'b100100010111;
   13666: result <= 12'b100100010111;
   13667: result <= 12'b100100011000;
   13668: result <= 12'b100100011000;
   13669: result <= 12'b100100011001;
   13670: result <= 12'b100100011001;
   13671: result <= 12'b100100011001;
   13672: result <= 12'b100100011010;
   13673: result <= 12'b100100011010;
   13674: result <= 12'b100100011011;
   13675: result <= 12'b100100011011;
   13676: result <= 12'b100100011011;
   13677: result <= 12'b100100011100;
   13678: result <= 12'b100100011100;
   13679: result <= 12'b100100011101;
   13680: result <= 12'b100100011101;
   13681: result <= 12'b100100011101;
   13682: result <= 12'b100100011110;
   13683: result <= 12'b100100011110;
   13684: result <= 12'b100100011111;
   13685: result <= 12'b100100011111;
   13686: result <= 12'b100100011111;
   13687: result <= 12'b100100100000;
   13688: result <= 12'b100100100000;
   13689: result <= 12'b100100100001;
   13690: result <= 12'b100100100001;
   13691: result <= 12'b100100100001;
   13692: result <= 12'b100100100010;
   13693: result <= 12'b100100100010;
   13694: result <= 12'b100100100011;
   13695: result <= 12'b100100100011;
   13696: result <= 12'b100100100011;
   13697: result <= 12'b100100100100;
   13698: result <= 12'b100100100100;
   13699: result <= 12'b100100100101;
   13700: result <= 12'b100100100101;
   13701: result <= 12'b100100100101;
   13702: result <= 12'b100100100110;
   13703: result <= 12'b100100100110;
   13704: result <= 12'b100100100111;
   13705: result <= 12'b100100100111;
   13706: result <= 12'b100100100111;
   13707: result <= 12'b100100101000;
   13708: result <= 12'b100100101000;
   13709: result <= 12'b100100101001;
   13710: result <= 12'b100100101001;
   13711: result <= 12'b100100101001;
   13712: result <= 12'b100100101010;
   13713: result <= 12'b100100101010;
   13714: result <= 12'b100100101011;
   13715: result <= 12'b100100101011;
   13716: result <= 12'b100100101011;
   13717: result <= 12'b100100101100;
   13718: result <= 12'b100100101100;
   13719: result <= 12'b100100101101;
   13720: result <= 12'b100100101101;
   13721: result <= 12'b100100101110;
   13722: result <= 12'b100100101110;
   13723: result <= 12'b100100101110;
   13724: result <= 12'b100100101111;
   13725: result <= 12'b100100101111;
   13726: result <= 12'b100100110000;
   13727: result <= 12'b100100110000;
   13728: result <= 12'b100100110000;
   13729: result <= 12'b100100110001;
   13730: result <= 12'b100100110001;
   13731: result <= 12'b100100110010;
   13732: result <= 12'b100100110010;
   13733: result <= 12'b100100110010;
   13734: result <= 12'b100100110011;
   13735: result <= 12'b100100110011;
   13736: result <= 12'b100100110100;
   13737: result <= 12'b100100110100;
   13738: result <= 12'b100100110101;
   13739: result <= 12'b100100110101;
   13740: result <= 12'b100100110101;
   13741: result <= 12'b100100110110;
   13742: result <= 12'b100100110110;
   13743: result <= 12'b100100110111;
   13744: result <= 12'b100100110111;
   13745: result <= 12'b100100110111;
   13746: result <= 12'b100100111000;
   13747: result <= 12'b100100111000;
   13748: result <= 12'b100100111001;
   13749: result <= 12'b100100111001;
   13750: result <= 12'b100100111010;
   13751: result <= 12'b100100111010;
   13752: result <= 12'b100100111010;
   13753: result <= 12'b100100111011;
   13754: result <= 12'b100100111011;
   13755: result <= 12'b100100111100;
   13756: result <= 12'b100100111100;
   13757: result <= 12'b100100111100;
   13758: result <= 12'b100100111101;
   13759: result <= 12'b100100111101;
   13760: result <= 12'b100100111110;
   13761: result <= 12'b100100111110;
   13762: result <= 12'b100100111111;
   13763: result <= 12'b100100111111;
   13764: result <= 12'b100100111111;
   13765: result <= 12'b100101000000;
   13766: result <= 12'b100101000000;
   13767: result <= 12'b100101000001;
   13768: result <= 12'b100101000001;
   13769: result <= 12'b100101000010;
   13770: result <= 12'b100101000010;
   13771: result <= 12'b100101000010;
   13772: result <= 12'b100101000011;
   13773: result <= 12'b100101000011;
   13774: result <= 12'b100101000100;
   13775: result <= 12'b100101000100;
   13776: result <= 12'b100101000100;
   13777: result <= 12'b100101000101;
   13778: result <= 12'b100101000101;
   13779: result <= 12'b100101000110;
   13780: result <= 12'b100101000110;
   13781: result <= 12'b100101000111;
   13782: result <= 12'b100101000111;
   13783: result <= 12'b100101000111;
   13784: result <= 12'b100101001000;
   13785: result <= 12'b100101001000;
   13786: result <= 12'b100101001001;
   13787: result <= 12'b100101001001;
   13788: result <= 12'b100101001010;
   13789: result <= 12'b100101001010;
   13790: result <= 12'b100101001010;
   13791: result <= 12'b100101001011;
   13792: result <= 12'b100101001011;
   13793: result <= 12'b100101001100;
   13794: result <= 12'b100101001100;
   13795: result <= 12'b100101001101;
   13796: result <= 12'b100101001101;
   13797: result <= 12'b100101001101;
   13798: result <= 12'b100101001110;
   13799: result <= 12'b100101001110;
   13800: result <= 12'b100101001111;
   13801: result <= 12'b100101001111;
   13802: result <= 12'b100101010000;
   13803: result <= 12'b100101010000;
   13804: result <= 12'b100101010000;
   13805: result <= 12'b100101010001;
   13806: result <= 12'b100101010001;
   13807: result <= 12'b100101010010;
   13808: result <= 12'b100101010010;
   13809: result <= 12'b100101010011;
   13810: result <= 12'b100101010011;
   13811: result <= 12'b100101010011;
   13812: result <= 12'b100101010100;
   13813: result <= 12'b100101010100;
   13814: result <= 12'b100101010101;
   13815: result <= 12'b100101010101;
   13816: result <= 12'b100101010110;
   13817: result <= 12'b100101010110;
   13818: result <= 12'b100101010111;
   13819: result <= 12'b100101010111;
   13820: result <= 12'b100101010111;
   13821: result <= 12'b100101011000;
   13822: result <= 12'b100101011000;
   13823: result <= 12'b100101011001;
   13824: result <= 12'b100101011001;
   13825: result <= 12'b100101011010;
   13826: result <= 12'b100101011010;
   13827: result <= 12'b100101011010;
   13828: result <= 12'b100101011011;
   13829: result <= 12'b100101011011;
   13830: result <= 12'b100101011100;
   13831: result <= 12'b100101011100;
   13832: result <= 12'b100101011101;
   13833: result <= 12'b100101011101;
   13834: result <= 12'b100101011110;
   13835: result <= 12'b100101011110;
   13836: result <= 12'b100101011110;
   13837: result <= 12'b100101011111;
   13838: result <= 12'b100101011111;
   13839: result <= 12'b100101100000;
   13840: result <= 12'b100101100000;
   13841: result <= 12'b100101100001;
   13842: result <= 12'b100101100001;
   13843: result <= 12'b100101100001;
   13844: result <= 12'b100101100010;
   13845: result <= 12'b100101100010;
   13846: result <= 12'b100101100011;
   13847: result <= 12'b100101100011;
   13848: result <= 12'b100101100100;
   13849: result <= 12'b100101100100;
   13850: result <= 12'b100101100101;
   13851: result <= 12'b100101100101;
   13852: result <= 12'b100101100101;
   13853: result <= 12'b100101100110;
   13854: result <= 12'b100101100110;
   13855: result <= 12'b100101100111;
   13856: result <= 12'b100101100111;
   13857: result <= 12'b100101101000;
   13858: result <= 12'b100101101000;
   13859: result <= 12'b100101101001;
   13860: result <= 12'b100101101001;
   13861: result <= 12'b100101101001;
   13862: result <= 12'b100101101010;
   13863: result <= 12'b100101101010;
   13864: result <= 12'b100101101011;
   13865: result <= 12'b100101101011;
   13866: result <= 12'b100101101100;
   13867: result <= 12'b100101101100;
   13868: result <= 12'b100101101101;
   13869: result <= 12'b100101101101;
   13870: result <= 12'b100101101101;
   13871: result <= 12'b100101101110;
   13872: result <= 12'b100101101110;
   13873: result <= 12'b100101101111;
   13874: result <= 12'b100101101111;
   13875: result <= 12'b100101110000;
   13876: result <= 12'b100101110000;
   13877: result <= 12'b100101110001;
   13878: result <= 12'b100101110001;
   13879: result <= 12'b100101110010;
   13880: result <= 12'b100101110010;
   13881: result <= 12'b100101110010;
   13882: result <= 12'b100101110011;
   13883: result <= 12'b100101110011;
   13884: result <= 12'b100101110100;
   13885: result <= 12'b100101110100;
   13886: result <= 12'b100101110101;
   13887: result <= 12'b100101110101;
   13888: result <= 12'b100101110110;
   13889: result <= 12'b100101110110;
   13890: result <= 12'b100101110110;
   13891: result <= 12'b100101110111;
   13892: result <= 12'b100101110111;
   13893: result <= 12'b100101111000;
   13894: result <= 12'b100101111000;
   13895: result <= 12'b100101111001;
   13896: result <= 12'b100101111001;
   13897: result <= 12'b100101111010;
   13898: result <= 12'b100101111010;
   13899: result <= 12'b100101111011;
   13900: result <= 12'b100101111011;
   13901: result <= 12'b100101111011;
   13902: result <= 12'b100101111100;
   13903: result <= 12'b100101111100;
   13904: result <= 12'b100101111101;
   13905: result <= 12'b100101111101;
   13906: result <= 12'b100101111110;
   13907: result <= 12'b100101111110;
   13908: result <= 12'b100101111111;
   13909: result <= 12'b100101111111;
   13910: result <= 12'b100110000000;
   13911: result <= 12'b100110000000;
   13912: result <= 12'b100110000001;
   13913: result <= 12'b100110000001;
   13914: result <= 12'b100110000001;
   13915: result <= 12'b100110000010;
   13916: result <= 12'b100110000010;
   13917: result <= 12'b100110000011;
   13918: result <= 12'b100110000011;
   13919: result <= 12'b100110000100;
   13920: result <= 12'b100110000100;
   13921: result <= 12'b100110000101;
   13922: result <= 12'b100110000101;
   13923: result <= 12'b100110000110;
   13924: result <= 12'b100110000110;
   13925: result <= 12'b100110000110;
   13926: result <= 12'b100110000111;
   13927: result <= 12'b100110000111;
   13928: result <= 12'b100110001000;
   13929: result <= 12'b100110001000;
   13930: result <= 12'b100110001001;
   13931: result <= 12'b100110001001;
   13932: result <= 12'b100110001010;
   13933: result <= 12'b100110001010;
   13934: result <= 12'b100110001011;
   13935: result <= 12'b100110001011;
   13936: result <= 12'b100110001100;
   13937: result <= 12'b100110001100;
   13938: result <= 12'b100110001101;
   13939: result <= 12'b100110001101;
   13940: result <= 12'b100110001101;
   13941: result <= 12'b100110001110;
   13942: result <= 12'b100110001110;
   13943: result <= 12'b100110001111;
   13944: result <= 12'b100110001111;
   13945: result <= 12'b100110010000;
   13946: result <= 12'b100110010000;
   13947: result <= 12'b100110010001;
   13948: result <= 12'b100110010001;
   13949: result <= 12'b100110010010;
   13950: result <= 12'b100110010010;
   13951: result <= 12'b100110010011;
   13952: result <= 12'b100110010011;
   13953: result <= 12'b100110010011;
   13954: result <= 12'b100110010100;
   13955: result <= 12'b100110010100;
   13956: result <= 12'b100110010101;
   13957: result <= 12'b100110010101;
   13958: result <= 12'b100110010110;
   13959: result <= 12'b100110010110;
   13960: result <= 12'b100110010111;
   13961: result <= 12'b100110010111;
   13962: result <= 12'b100110011000;
   13963: result <= 12'b100110011000;
   13964: result <= 12'b100110011001;
   13965: result <= 12'b100110011001;
   13966: result <= 12'b100110011010;
   13967: result <= 12'b100110011010;
   13968: result <= 12'b100110011011;
   13969: result <= 12'b100110011011;
   13970: result <= 12'b100110011011;
   13971: result <= 12'b100110011100;
   13972: result <= 12'b100110011100;
   13973: result <= 12'b100110011101;
   13974: result <= 12'b100110011101;
   13975: result <= 12'b100110011110;
   13976: result <= 12'b100110011110;
   13977: result <= 12'b100110011111;
   13978: result <= 12'b100110011111;
   13979: result <= 12'b100110100000;
   13980: result <= 12'b100110100000;
   13981: result <= 12'b100110100001;
   13982: result <= 12'b100110100001;
   13983: result <= 12'b100110100010;
   13984: result <= 12'b100110100010;
   13985: result <= 12'b100110100011;
   13986: result <= 12'b100110100011;
   13987: result <= 12'b100110100100;
   13988: result <= 12'b100110100100;
   13989: result <= 12'b100110100101;
   13990: result <= 12'b100110100101;
   13991: result <= 12'b100110100101;
   13992: result <= 12'b100110100110;
   13993: result <= 12'b100110100110;
   13994: result <= 12'b100110100111;
   13995: result <= 12'b100110100111;
   13996: result <= 12'b100110101000;
   13997: result <= 12'b100110101000;
   13998: result <= 12'b100110101001;
   13999: result <= 12'b100110101001;
   14000: result <= 12'b100110101010;
   14001: result <= 12'b100110101010;
   14002: result <= 12'b100110101011;
   14003: result <= 12'b100110101011;
   14004: result <= 12'b100110101100;
   14005: result <= 12'b100110101100;
   14006: result <= 12'b100110101101;
   14007: result <= 12'b100110101101;
   14008: result <= 12'b100110101110;
   14009: result <= 12'b100110101110;
   14010: result <= 12'b100110101111;
   14011: result <= 12'b100110101111;
   14012: result <= 12'b100110110000;
   14013: result <= 12'b100110110000;
   14014: result <= 12'b100110110001;
   14015: result <= 12'b100110110001;
   14016: result <= 12'b100110110001;
   14017: result <= 12'b100110110010;
   14018: result <= 12'b100110110010;
   14019: result <= 12'b100110110011;
   14020: result <= 12'b100110110011;
   14021: result <= 12'b100110110100;
   14022: result <= 12'b100110110100;
   14023: result <= 12'b100110110101;
   14024: result <= 12'b100110110101;
   14025: result <= 12'b100110110110;
   14026: result <= 12'b100110110110;
   14027: result <= 12'b100110110111;
   14028: result <= 12'b100110110111;
   14029: result <= 12'b100110111000;
   14030: result <= 12'b100110111000;
   14031: result <= 12'b100110111001;
   14032: result <= 12'b100110111001;
   14033: result <= 12'b100110111010;
   14034: result <= 12'b100110111010;
   14035: result <= 12'b100110111011;
   14036: result <= 12'b100110111011;
   14037: result <= 12'b100110111100;
   14038: result <= 12'b100110111100;
   14039: result <= 12'b100110111101;
   14040: result <= 12'b100110111101;
   14041: result <= 12'b100110111110;
   14042: result <= 12'b100110111110;
   14043: result <= 12'b100110111111;
   14044: result <= 12'b100110111111;
   14045: result <= 12'b100111000000;
   14046: result <= 12'b100111000000;
   14047: result <= 12'b100111000001;
   14048: result <= 12'b100111000001;
   14049: result <= 12'b100111000010;
   14050: result <= 12'b100111000010;
   14051: result <= 12'b100111000011;
   14052: result <= 12'b100111000011;
   14053: result <= 12'b100111000100;
   14054: result <= 12'b100111000100;
   14055: result <= 12'b100111000100;
   14056: result <= 12'b100111000101;
   14057: result <= 12'b100111000101;
   14058: result <= 12'b100111000110;
   14059: result <= 12'b100111000110;
   14060: result <= 12'b100111000111;
   14061: result <= 12'b100111000111;
   14062: result <= 12'b100111001000;
   14063: result <= 12'b100111001000;
   14064: result <= 12'b100111001001;
   14065: result <= 12'b100111001001;
   14066: result <= 12'b100111001010;
   14067: result <= 12'b100111001010;
   14068: result <= 12'b100111001011;
   14069: result <= 12'b100111001011;
   14070: result <= 12'b100111001100;
   14071: result <= 12'b100111001100;
   14072: result <= 12'b100111001101;
   14073: result <= 12'b100111001101;
   14074: result <= 12'b100111001110;
   14075: result <= 12'b100111001110;
   14076: result <= 12'b100111001111;
   14077: result <= 12'b100111001111;
   14078: result <= 12'b100111010000;
   14079: result <= 12'b100111010000;
   14080: result <= 12'b100111010001;
   14081: result <= 12'b100111010001;
   14082: result <= 12'b100111010010;
   14083: result <= 12'b100111010010;
   14084: result <= 12'b100111010011;
   14085: result <= 12'b100111010011;
   14086: result <= 12'b100111010100;
   14087: result <= 12'b100111010100;
   14088: result <= 12'b100111010101;
   14089: result <= 12'b100111010101;
   14090: result <= 12'b100111010110;
   14091: result <= 12'b100111010110;
   14092: result <= 12'b100111010111;
   14093: result <= 12'b100111010111;
   14094: result <= 12'b100111011000;
   14095: result <= 12'b100111011000;
   14096: result <= 12'b100111011001;
   14097: result <= 12'b100111011001;
   14098: result <= 12'b100111011010;
   14099: result <= 12'b100111011010;
   14100: result <= 12'b100111011011;
   14101: result <= 12'b100111011011;
   14102: result <= 12'b100111011100;
   14103: result <= 12'b100111011100;
   14104: result <= 12'b100111011101;
   14105: result <= 12'b100111011101;
   14106: result <= 12'b100111011110;
   14107: result <= 12'b100111011110;
   14108: result <= 12'b100111011111;
   14109: result <= 12'b100111011111;
   14110: result <= 12'b100111100000;
   14111: result <= 12'b100111100000;
   14112: result <= 12'b100111100001;
   14113: result <= 12'b100111100001;
   14114: result <= 12'b100111100010;
   14115: result <= 12'b100111100010;
   14116: result <= 12'b100111100011;
   14117: result <= 12'b100111100011;
   14118: result <= 12'b100111100100;
   14119: result <= 12'b100111100100;
   14120: result <= 12'b100111100101;
   14121: result <= 12'b100111100101;
   14122: result <= 12'b100111100110;
   14123: result <= 12'b100111100111;
   14124: result <= 12'b100111100111;
   14125: result <= 12'b100111101000;
   14126: result <= 12'b100111101000;
   14127: result <= 12'b100111101001;
   14128: result <= 12'b100111101001;
   14129: result <= 12'b100111101010;
   14130: result <= 12'b100111101010;
   14131: result <= 12'b100111101011;
   14132: result <= 12'b100111101011;
   14133: result <= 12'b100111101100;
   14134: result <= 12'b100111101100;
   14135: result <= 12'b100111101101;
   14136: result <= 12'b100111101101;
   14137: result <= 12'b100111101110;
   14138: result <= 12'b100111101110;
   14139: result <= 12'b100111101111;
   14140: result <= 12'b100111101111;
   14141: result <= 12'b100111110000;
   14142: result <= 12'b100111110000;
   14143: result <= 12'b100111110001;
   14144: result <= 12'b100111110001;
   14145: result <= 12'b100111110010;
   14146: result <= 12'b100111110010;
   14147: result <= 12'b100111110011;
   14148: result <= 12'b100111110011;
   14149: result <= 12'b100111110100;
   14150: result <= 12'b100111110100;
   14151: result <= 12'b100111110101;
   14152: result <= 12'b100111110101;
   14153: result <= 12'b100111110110;
   14154: result <= 12'b100111110110;
   14155: result <= 12'b100111110111;
   14156: result <= 12'b100111110111;
   14157: result <= 12'b100111111000;
   14158: result <= 12'b100111111000;
   14159: result <= 12'b100111111001;
   14160: result <= 12'b100111111001;
   14161: result <= 12'b100111111010;
   14162: result <= 12'b100111111011;
   14163: result <= 12'b100111111011;
   14164: result <= 12'b100111111100;
   14165: result <= 12'b100111111100;
   14166: result <= 12'b100111111101;
   14167: result <= 12'b100111111101;
   14168: result <= 12'b100111111110;
   14169: result <= 12'b100111111110;
   14170: result <= 12'b100111111111;
   14171: result <= 12'b100111111111;
   14172: result <= 12'b101000000000;
   14173: result <= 12'b101000000000;
   14174: result <= 12'b101000000001;
   14175: result <= 12'b101000000001;
   14176: result <= 12'b101000000010;
   14177: result <= 12'b101000000010;
   14178: result <= 12'b101000000011;
   14179: result <= 12'b101000000011;
   14180: result <= 12'b101000000100;
   14181: result <= 12'b101000000100;
   14182: result <= 12'b101000000101;
   14183: result <= 12'b101000000101;
   14184: result <= 12'b101000000110;
   14185: result <= 12'b101000000110;
   14186: result <= 12'b101000000111;
   14187: result <= 12'b101000001000;
   14188: result <= 12'b101000001000;
   14189: result <= 12'b101000001001;
   14190: result <= 12'b101000001001;
   14191: result <= 12'b101000001010;
   14192: result <= 12'b101000001010;
   14193: result <= 12'b101000001011;
   14194: result <= 12'b101000001011;
   14195: result <= 12'b101000001100;
   14196: result <= 12'b101000001100;
   14197: result <= 12'b101000001101;
   14198: result <= 12'b101000001101;
   14199: result <= 12'b101000001110;
   14200: result <= 12'b101000001110;
   14201: result <= 12'b101000001111;
   14202: result <= 12'b101000001111;
   14203: result <= 12'b101000010000;
   14204: result <= 12'b101000010000;
   14205: result <= 12'b101000010001;
   14206: result <= 12'b101000010001;
   14207: result <= 12'b101000010010;
   14208: result <= 12'b101000010011;
   14209: result <= 12'b101000010011;
   14210: result <= 12'b101000010100;
   14211: result <= 12'b101000010100;
   14212: result <= 12'b101000010101;
   14213: result <= 12'b101000010101;
   14214: result <= 12'b101000010110;
   14215: result <= 12'b101000010110;
   14216: result <= 12'b101000010111;
   14217: result <= 12'b101000010111;
   14218: result <= 12'b101000011000;
   14219: result <= 12'b101000011000;
   14220: result <= 12'b101000011001;
   14221: result <= 12'b101000011001;
   14222: result <= 12'b101000011010;
   14223: result <= 12'b101000011010;
   14224: result <= 12'b101000011011;
   14225: result <= 12'b101000011100;
   14226: result <= 12'b101000011100;
   14227: result <= 12'b101000011101;
   14228: result <= 12'b101000011101;
   14229: result <= 12'b101000011110;
   14230: result <= 12'b101000011110;
   14231: result <= 12'b101000011111;
   14232: result <= 12'b101000011111;
   14233: result <= 12'b101000100000;
   14234: result <= 12'b101000100000;
   14235: result <= 12'b101000100001;
   14236: result <= 12'b101000100001;
   14237: result <= 12'b101000100010;
   14238: result <= 12'b101000100010;
   14239: result <= 12'b101000100011;
   14240: result <= 12'b101000100100;
   14241: result <= 12'b101000100100;
   14242: result <= 12'b101000100101;
   14243: result <= 12'b101000100101;
   14244: result <= 12'b101000100110;
   14245: result <= 12'b101000100110;
   14246: result <= 12'b101000100111;
   14247: result <= 12'b101000100111;
   14248: result <= 12'b101000101000;
   14249: result <= 12'b101000101000;
   14250: result <= 12'b101000101001;
   14251: result <= 12'b101000101001;
   14252: result <= 12'b101000101010;
   14253: result <= 12'b101000101010;
   14254: result <= 12'b101000101011;
   14255: result <= 12'b101000101100;
   14256: result <= 12'b101000101100;
   14257: result <= 12'b101000101101;
   14258: result <= 12'b101000101101;
   14259: result <= 12'b101000101110;
   14260: result <= 12'b101000101110;
   14261: result <= 12'b101000101111;
   14262: result <= 12'b101000101111;
   14263: result <= 12'b101000110000;
   14264: result <= 12'b101000110000;
   14265: result <= 12'b101000110001;
   14266: result <= 12'b101000110001;
   14267: result <= 12'b101000110010;
   14268: result <= 12'b101000110011;
   14269: result <= 12'b101000110011;
   14270: result <= 12'b101000110100;
   14271: result <= 12'b101000110100;
   14272: result <= 12'b101000110101;
   14273: result <= 12'b101000110101;
   14274: result <= 12'b101000110110;
   14275: result <= 12'b101000110110;
   14276: result <= 12'b101000110111;
   14277: result <= 12'b101000110111;
   14278: result <= 12'b101000111000;
   14279: result <= 12'b101000111001;
   14280: result <= 12'b101000111001;
   14281: result <= 12'b101000111010;
   14282: result <= 12'b101000111010;
   14283: result <= 12'b101000111011;
   14284: result <= 12'b101000111011;
   14285: result <= 12'b101000111100;
   14286: result <= 12'b101000111100;
   14287: result <= 12'b101000111101;
   14288: result <= 12'b101000111101;
   14289: result <= 12'b101000111110;
   14290: result <= 12'b101000111111;
   14291: result <= 12'b101000111111;
   14292: result <= 12'b101001000000;
   14293: result <= 12'b101001000000;
   14294: result <= 12'b101001000001;
   14295: result <= 12'b101001000001;
   14296: result <= 12'b101001000010;
   14297: result <= 12'b101001000010;
   14298: result <= 12'b101001000011;
   14299: result <= 12'b101001000011;
   14300: result <= 12'b101001000100;
   14301: result <= 12'b101001000101;
   14302: result <= 12'b101001000101;
   14303: result <= 12'b101001000110;
   14304: result <= 12'b101001000110;
   14305: result <= 12'b101001000111;
   14306: result <= 12'b101001000111;
   14307: result <= 12'b101001001000;
   14308: result <= 12'b101001001000;
   14309: result <= 12'b101001001001;
   14310: result <= 12'b101001001001;
   14311: result <= 12'b101001001010;
   14312: result <= 12'b101001001011;
   14313: result <= 12'b101001001011;
   14314: result <= 12'b101001001100;
   14315: result <= 12'b101001001100;
   14316: result <= 12'b101001001101;
   14317: result <= 12'b101001001101;
   14318: result <= 12'b101001001110;
   14319: result <= 12'b101001001110;
   14320: result <= 12'b101001001111;
   14321: result <= 12'b101001010000;
   14322: result <= 12'b101001010000;
   14323: result <= 12'b101001010001;
   14324: result <= 12'b101001010001;
   14325: result <= 12'b101001010010;
   14326: result <= 12'b101001010010;
   14327: result <= 12'b101001010011;
   14328: result <= 12'b101001010011;
   14329: result <= 12'b101001010100;
   14330: result <= 12'b101001010101;
   14331: result <= 12'b101001010101;
   14332: result <= 12'b101001010110;
   14333: result <= 12'b101001010110;
   14334: result <= 12'b101001010111;
   14335: result <= 12'b101001010111;
   14336: result <= 12'b101001011000;
   14337: result <= 12'b101001011000;
   14338: result <= 12'b101001011001;
   14339: result <= 12'b101001011010;
   14340: result <= 12'b101001011010;
   14341: result <= 12'b101001011011;
   14342: result <= 12'b101001011011;
   14343: result <= 12'b101001011100;
   14344: result <= 12'b101001011100;
   14345: result <= 12'b101001011101;
   14346: result <= 12'b101001011101;
   14347: result <= 12'b101001011110;
   14348: result <= 12'b101001011111;
   14349: result <= 12'b101001011111;
   14350: result <= 12'b101001100000;
   14351: result <= 12'b101001100000;
   14352: result <= 12'b101001100001;
   14353: result <= 12'b101001100001;
   14354: result <= 12'b101001100010;
   14355: result <= 12'b101001100010;
   14356: result <= 12'b101001100011;
   14357: result <= 12'b101001100100;
   14358: result <= 12'b101001100100;
   14359: result <= 12'b101001100101;
   14360: result <= 12'b101001100101;
   14361: result <= 12'b101001100110;
   14362: result <= 12'b101001100110;
   14363: result <= 12'b101001100111;
   14364: result <= 12'b101001100111;
   14365: result <= 12'b101001101000;
   14366: result <= 12'b101001101001;
   14367: result <= 12'b101001101001;
   14368: result <= 12'b101001101010;
   14369: result <= 12'b101001101010;
   14370: result <= 12'b101001101011;
   14371: result <= 12'b101001101011;
   14372: result <= 12'b101001101100;
   14373: result <= 12'b101001101101;
   14374: result <= 12'b101001101101;
   14375: result <= 12'b101001101110;
   14376: result <= 12'b101001101110;
   14377: result <= 12'b101001101111;
   14378: result <= 12'b101001101111;
   14379: result <= 12'b101001110000;
   14380: result <= 12'b101001110000;
   14381: result <= 12'b101001110001;
   14382: result <= 12'b101001110010;
   14383: result <= 12'b101001110010;
   14384: result <= 12'b101001110011;
   14385: result <= 12'b101001110011;
   14386: result <= 12'b101001110100;
   14387: result <= 12'b101001110100;
   14388: result <= 12'b101001110101;
   14389: result <= 12'b101001110110;
   14390: result <= 12'b101001110110;
   14391: result <= 12'b101001110111;
   14392: result <= 12'b101001110111;
   14393: result <= 12'b101001111000;
   14394: result <= 12'b101001111000;
   14395: result <= 12'b101001111001;
   14396: result <= 12'b101001111010;
   14397: result <= 12'b101001111010;
   14398: result <= 12'b101001111011;
   14399: result <= 12'b101001111011;
   14400: result <= 12'b101001111100;
   14401: result <= 12'b101001111100;
   14402: result <= 12'b101001111101;
   14403: result <= 12'b101001111110;
   14404: result <= 12'b101001111110;
   14405: result <= 12'b101001111111;
   14406: result <= 12'b101001111111;
   14407: result <= 12'b101010000000;
   14408: result <= 12'b101010000000;
   14409: result <= 12'b101010000001;
   14410: result <= 12'b101010000010;
   14411: result <= 12'b101010000010;
   14412: result <= 12'b101010000011;
   14413: result <= 12'b101010000011;
   14414: result <= 12'b101010000100;
   14415: result <= 12'b101010000100;
   14416: result <= 12'b101010000101;
   14417: result <= 12'b101010000110;
   14418: result <= 12'b101010000110;
   14419: result <= 12'b101010000111;
   14420: result <= 12'b101010000111;
   14421: result <= 12'b101010001000;
   14422: result <= 12'b101010001000;
   14423: result <= 12'b101010001001;
   14424: result <= 12'b101010001010;
   14425: result <= 12'b101010001010;
   14426: result <= 12'b101010001011;
   14427: result <= 12'b101010001011;
   14428: result <= 12'b101010001100;
   14429: result <= 12'b101010001100;
   14430: result <= 12'b101010001101;
   14431: result <= 12'b101010001110;
   14432: result <= 12'b101010001110;
   14433: result <= 12'b101010001111;
   14434: result <= 12'b101010001111;
   14435: result <= 12'b101010010000;
   14436: result <= 12'b101010010000;
   14437: result <= 12'b101010010001;
   14438: result <= 12'b101010010010;
   14439: result <= 12'b101010010010;
   14440: result <= 12'b101010010011;
   14441: result <= 12'b101010010011;
   14442: result <= 12'b101010010100;
   14443: result <= 12'b101010010100;
   14444: result <= 12'b101010010101;
   14445: result <= 12'b101010010110;
   14446: result <= 12'b101010010110;
   14447: result <= 12'b101010010111;
   14448: result <= 12'b101010010111;
   14449: result <= 12'b101010011000;
   14450: result <= 12'b101010011001;
   14451: result <= 12'b101010011001;
   14452: result <= 12'b101010011010;
   14453: result <= 12'b101010011010;
   14454: result <= 12'b101010011011;
   14455: result <= 12'b101010011011;
   14456: result <= 12'b101010011100;
   14457: result <= 12'b101010011101;
   14458: result <= 12'b101010011101;
   14459: result <= 12'b101010011110;
   14460: result <= 12'b101010011110;
   14461: result <= 12'b101010011111;
   14462: result <= 12'b101010011111;
   14463: result <= 12'b101010100000;
   14464: result <= 12'b101010100001;
   14465: result <= 12'b101010100001;
   14466: result <= 12'b101010100010;
   14467: result <= 12'b101010100010;
   14468: result <= 12'b101010100011;
   14469: result <= 12'b101010100100;
   14470: result <= 12'b101010100100;
   14471: result <= 12'b101010100101;
   14472: result <= 12'b101010100101;
   14473: result <= 12'b101010100110;
   14474: result <= 12'b101010100110;
   14475: result <= 12'b101010100111;
   14476: result <= 12'b101010101000;
   14477: result <= 12'b101010101000;
   14478: result <= 12'b101010101001;
   14479: result <= 12'b101010101001;
   14480: result <= 12'b101010101010;
   14481: result <= 12'b101010101011;
   14482: result <= 12'b101010101011;
   14483: result <= 12'b101010101100;
   14484: result <= 12'b101010101100;
   14485: result <= 12'b101010101101;
   14486: result <= 12'b101010101101;
   14487: result <= 12'b101010101110;
   14488: result <= 12'b101010101111;
   14489: result <= 12'b101010101111;
   14490: result <= 12'b101010110000;
   14491: result <= 12'b101010110000;
   14492: result <= 12'b101010110001;
   14493: result <= 12'b101010110010;
   14494: result <= 12'b101010110010;
   14495: result <= 12'b101010110011;
   14496: result <= 12'b101010110011;
   14497: result <= 12'b101010110100;
   14498: result <= 12'b101010110101;
   14499: result <= 12'b101010110101;
   14500: result <= 12'b101010110110;
   14501: result <= 12'b101010110110;
   14502: result <= 12'b101010110111;
   14503: result <= 12'b101010110111;
   14504: result <= 12'b101010111000;
   14505: result <= 12'b101010111001;
   14506: result <= 12'b101010111001;
   14507: result <= 12'b101010111010;
   14508: result <= 12'b101010111010;
   14509: result <= 12'b101010111011;
   14510: result <= 12'b101010111100;
   14511: result <= 12'b101010111100;
   14512: result <= 12'b101010111101;
   14513: result <= 12'b101010111101;
   14514: result <= 12'b101010111110;
   14515: result <= 12'b101010111111;
   14516: result <= 12'b101010111111;
   14517: result <= 12'b101011000000;
   14518: result <= 12'b101011000000;
   14519: result <= 12'b101011000001;
   14520: result <= 12'b101011000010;
   14521: result <= 12'b101011000010;
   14522: result <= 12'b101011000011;
   14523: result <= 12'b101011000011;
   14524: result <= 12'b101011000100;
   14525: result <= 12'b101011000101;
   14526: result <= 12'b101011000101;
   14527: result <= 12'b101011000110;
   14528: result <= 12'b101011000110;
   14529: result <= 12'b101011000111;
   14530: result <= 12'b101011000111;
   14531: result <= 12'b101011001000;
   14532: result <= 12'b101011001001;
   14533: result <= 12'b101011001001;
   14534: result <= 12'b101011001010;
   14535: result <= 12'b101011001010;
   14536: result <= 12'b101011001011;
   14537: result <= 12'b101011001100;
   14538: result <= 12'b101011001100;
   14539: result <= 12'b101011001101;
   14540: result <= 12'b101011001101;
   14541: result <= 12'b101011001110;
   14542: result <= 12'b101011001111;
   14543: result <= 12'b101011001111;
   14544: result <= 12'b101011010000;
   14545: result <= 12'b101011010000;
   14546: result <= 12'b101011010001;
   14547: result <= 12'b101011010010;
   14548: result <= 12'b101011010010;
   14549: result <= 12'b101011010011;
   14550: result <= 12'b101011010011;
   14551: result <= 12'b101011010100;
   14552: result <= 12'b101011010101;
   14553: result <= 12'b101011010101;
   14554: result <= 12'b101011010110;
   14555: result <= 12'b101011010110;
   14556: result <= 12'b101011010111;
   14557: result <= 12'b101011011000;
   14558: result <= 12'b101011011000;
   14559: result <= 12'b101011011001;
   14560: result <= 12'b101011011001;
   14561: result <= 12'b101011011010;
   14562: result <= 12'b101011011011;
   14563: result <= 12'b101011011011;
   14564: result <= 12'b101011011100;
   14565: result <= 12'b101011011100;
   14566: result <= 12'b101011011101;
   14567: result <= 12'b101011011110;
   14568: result <= 12'b101011011110;
   14569: result <= 12'b101011011111;
   14570: result <= 12'b101011011111;
   14571: result <= 12'b101011100000;
   14572: result <= 12'b101011100001;
   14573: result <= 12'b101011100001;
   14574: result <= 12'b101011100010;
   14575: result <= 12'b101011100010;
   14576: result <= 12'b101011100011;
   14577: result <= 12'b101011100100;
   14578: result <= 12'b101011100100;
   14579: result <= 12'b101011100101;
   14580: result <= 12'b101011100101;
   14581: result <= 12'b101011100110;
   14582: result <= 12'b101011100111;
   14583: result <= 12'b101011100111;
   14584: result <= 12'b101011101000;
   14585: result <= 12'b101011101001;
   14586: result <= 12'b101011101001;
   14587: result <= 12'b101011101010;
   14588: result <= 12'b101011101010;
   14589: result <= 12'b101011101011;
   14590: result <= 12'b101011101100;
   14591: result <= 12'b101011101100;
   14592: result <= 12'b101011101101;
   14593: result <= 12'b101011101101;
   14594: result <= 12'b101011101110;
   14595: result <= 12'b101011101111;
   14596: result <= 12'b101011101111;
   14597: result <= 12'b101011110000;
   14598: result <= 12'b101011110000;
   14599: result <= 12'b101011110001;
   14600: result <= 12'b101011110010;
   14601: result <= 12'b101011110010;
   14602: result <= 12'b101011110011;
   14603: result <= 12'b101011110011;
   14604: result <= 12'b101011110100;
   14605: result <= 12'b101011110101;
   14606: result <= 12'b101011110101;
   14607: result <= 12'b101011110110;
   14608: result <= 12'b101011110111;
   14609: result <= 12'b101011110111;
   14610: result <= 12'b101011111000;
   14611: result <= 12'b101011111000;
   14612: result <= 12'b101011111001;
   14613: result <= 12'b101011111010;
   14614: result <= 12'b101011111010;
   14615: result <= 12'b101011111011;
   14616: result <= 12'b101011111011;
   14617: result <= 12'b101011111100;
   14618: result <= 12'b101011111101;
   14619: result <= 12'b101011111101;
   14620: result <= 12'b101011111110;
   14621: result <= 12'b101011111110;
   14622: result <= 12'b101011111111;
   14623: result <= 12'b101100000000;
   14624: result <= 12'b101100000000;
   14625: result <= 12'b101100000001;
   14626: result <= 12'b101100000010;
   14627: result <= 12'b101100000010;
   14628: result <= 12'b101100000011;
   14629: result <= 12'b101100000011;
   14630: result <= 12'b101100000100;
   14631: result <= 12'b101100000101;
   14632: result <= 12'b101100000101;
   14633: result <= 12'b101100000110;
   14634: result <= 12'b101100000110;
   14635: result <= 12'b101100000111;
   14636: result <= 12'b101100001000;
   14637: result <= 12'b101100001000;
   14638: result <= 12'b101100001001;
   14639: result <= 12'b101100001010;
   14640: result <= 12'b101100001010;
   14641: result <= 12'b101100001011;
   14642: result <= 12'b101100001011;
   14643: result <= 12'b101100001100;
   14644: result <= 12'b101100001101;
   14645: result <= 12'b101100001101;
   14646: result <= 12'b101100001110;
   14647: result <= 12'b101100001110;
   14648: result <= 12'b101100001111;
   14649: result <= 12'b101100010000;
   14650: result <= 12'b101100010000;
   14651: result <= 12'b101100010001;
   14652: result <= 12'b101100010010;
   14653: result <= 12'b101100010010;
   14654: result <= 12'b101100010011;
   14655: result <= 12'b101100010011;
   14656: result <= 12'b101100010100;
   14657: result <= 12'b101100010101;
   14658: result <= 12'b101100010101;
   14659: result <= 12'b101100010110;
   14660: result <= 12'b101100010110;
   14661: result <= 12'b101100010111;
   14662: result <= 12'b101100011000;
   14663: result <= 12'b101100011000;
   14664: result <= 12'b101100011001;
   14665: result <= 12'b101100011010;
   14666: result <= 12'b101100011010;
   14667: result <= 12'b101100011011;
   14668: result <= 12'b101100011011;
   14669: result <= 12'b101100011100;
   14670: result <= 12'b101100011101;
   14671: result <= 12'b101100011101;
   14672: result <= 12'b101100011110;
   14673: result <= 12'b101100011111;
   14674: result <= 12'b101100011111;
   14675: result <= 12'b101100100000;
   14676: result <= 12'b101100100000;
   14677: result <= 12'b101100100001;
   14678: result <= 12'b101100100010;
   14679: result <= 12'b101100100010;
   14680: result <= 12'b101100100011;
   14681: result <= 12'b101100100100;
   14682: result <= 12'b101100100100;
   14683: result <= 12'b101100100101;
   14684: result <= 12'b101100100101;
   14685: result <= 12'b101100100110;
   14686: result <= 12'b101100100111;
   14687: result <= 12'b101100100111;
   14688: result <= 12'b101100101000;
   14689: result <= 12'b101100101001;
   14690: result <= 12'b101100101001;
   14691: result <= 12'b101100101010;
   14692: result <= 12'b101100101010;
   14693: result <= 12'b101100101011;
   14694: result <= 12'b101100101100;
   14695: result <= 12'b101100101100;
   14696: result <= 12'b101100101101;
   14697: result <= 12'b101100101110;
   14698: result <= 12'b101100101110;
   14699: result <= 12'b101100101111;
   14700: result <= 12'b101100101111;
   14701: result <= 12'b101100110000;
   14702: result <= 12'b101100110001;
   14703: result <= 12'b101100110001;
   14704: result <= 12'b101100110010;
   14705: result <= 12'b101100110011;
   14706: result <= 12'b101100110011;
   14707: result <= 12'b101100110100;
   14708: result <= 12'b101100110100;
   14709: result <= 12'b101100110101;
   14710: result <= 12'b101100110110;
   14711: result <= 12'b101100110110;
   14712: result <= 12'b101100110111;
   14713: result <= 12'b101100111000;
   14714: result <= 12'b101100111000;
   14715: result <= 12'b101100111001;
   14716: result <= 12'b101100111001;
   14717: result <= 12'b101100111010;
   14718: result <= 12'b101100111011;
   14719: result <= 12'b101100111011;
   14720: result <= 12'b101100111100;
   14721: result <= 12'b101100111101;
   14722: result <= 12'b101100111101;
   14723: result <= 12'b101100111110;
   14724: result <= 12'b101100111111;
   14725: result <= 12'b101100111111;
   14726: result <= 12'b101101000000;
   14727: result <= 12'b101101000000;
   14728: result <= 12'b101101000001;
   14729: result <= 12'b101101000010;
   14730: result <= 12'b101101000010;
   14731: result <= 12'b101101000011;
   14732: result <= 12'b101101000100;
   14733: result <= 12'b101101000100;
   14734: result <= 12'b101101000101;
   14735: result <= 12'b101101000101;
   14736: result <= 12'b101101000110;
   14737: result <= 12'b101101000111;
   14738: result <= 12'b101101000111;
   14739: result <= 12'b101101001000;
   14740: result <= 12'b101101001001;
   14741: result <= 12'b101101001001;
   14742: result <= 12'b101101001010;
   14743: result <= 12'b101101001011;
   14744: result <= 12'b101101001011;
   14745: result <= 12'b101101001100;
   14746: result <= 12'b101101001100;
   14747: result <= 12'b101101001101;
   14748: result <= 12'b101101001110;
   14749: result <= 12'b101101001110;
   14750: result <= 12'b101101001111;
   14751: result <= 12'b101101010000;
   14752: result <= 12'b101101010000;
   14753: result <= 12'b101101010001;
   14754: result <= 12'b101101010010;
   14755: result <= 12'b101101010010;
   14756: result <= 12'b101101010011;
   14757: result <= 12'b101101010011;
   14758: result <= 12'b101101010100;
   14759: result <= 12'b101101010101;
   14760: result <= 12'b101101010101;
   14761: result <= 12'b101101010110;
   14762: result <= 12'b101101010111;
   14763: result <= 12'b101101010111;
   14764: result <= 12'b101101011000;
   14765: result <= 12'b101101011001;
   14766: result <= 12'b101101011001;
   14767: result <= 12'b101101011010;
   14768: result <= 12'b101101011010;
   14769: result <= 12'b101101011011;
   14770: result <= 12'b101101011100;
   14771: result <= 12'b101101011100;
   14772: result <= 12'b101101011101;
   14773: result <= 12'b101101011110;
   14774: result <= 12'b101101011110;
   14775: result <= 12'b101101011111;
   14776: result <= 12'b101101100000;
   14777: result <= 12'b101101100000;
   14778: result <= 12'b101101100001;
   14779: result <= 12'b101101100010;
   14780: result <= 12'b101101100010;
   14781: result <= 12'b101101100011;
   14782: result <= 12'b101101100011;
   14783: result <= 12'b101101100100;
   14784: result <= 12'b101101100101;
   14785: result <= 12'b101101100101;
   14786: result <= 12'b101101100110;
   14787: result <= 12'b101101100111;
   14788: result <= 12'b101101100111;
   14789: result <= 12'b101101101000;
   14790: result <= 12'b101101101001;
   14791: result <= 12'b101101101001;
   14792: result <= 12'b101101101010;
   14793: result <= 12'b101101101011;
   14794: result <= 12'b101101101011;
   14795: result <= 12'b101101101100;
   14796: result <= 12'b101101101100;
   14797: result <= 12'b101101101101;
   14798: result <= 12'b101101101110;
   14799: result <= 12'b101101101110;
   14800: result <= 12'b101101101111;
   14801: result <= 12'b101101110000;
   14802: result <= 12'b101101110000;
   14803: result <= 12'b101101110001;
   14804: result <= 12'b101101110010;
   14805: result <= 12'b101101110010;
   14806: result <= 12'b101101110011;
   14807: result <= 12'b101101110100;
   14808: result <= 12'b101101110100;
   14809: result <= 12'b101101110101;
   14810: result <= 12'b101101110101;
   14811: result <= 12'b101101110110;
   14812: result <= 12'b101101110111;
   14813: result <= 12'b101101110111;
   14814: result <= 12'b101101111000;
   14815: result <= 12'b101101111001;
   14816: result <= 12'b101101111001;
   14817: result <= 12'b101101111010;
   14818: result <= 12'b101101111011;
   14819: result <= 12'b101101111011;
   14820: result <= 12'b101101111100;
   14821: result <= 12'b101101111101;
   14822: result <= 12'b101101111101;
   14823: result <= 12'b101101111110;
   14824: result <= 12'b101101111111;
   14825: result <= 12'b101101111111;
   14826: result <= 12'b101110000000;
   14827: result <= 12'b101110000001;
   14828: result <= 12'b101110000001;
   14829: result <= 12'b101110000010;
   14830: result <= 12'b101110000010;
   14831: result <= 12'b101110000011;
   14832: result <= 12'b101110000100;
   14833: result <= 12'b101110000100;
   14834: result <= 12'b101110000101;
   14835: result <= 12'b101110000110;
   14836: result <= 12'b101110000110;
   14837: result <= 12'b101110000111;
   14838: result <= 12'b101110001000;
   14839: result <= 12'b101110001000;
   14840: result <= 12'b101110001001;
   14841: result <= 12'b101110001010;
   14842: result <= 12'b101110001010;
   14843: result <= 12'b101110001011;
   14844: result <= 12'b101110001100;
   14845: result <= 12'b101110001100;
   14846: result <= 12'b101110001101;
   14847: result <= 12'b101110001110;
   14848: result <= 12'b101110001110;
   14849: result <= 12'b101110001111;
   14850: result <= 12'b101110001111;
   14851: result <= 12'b101110010000;
   14852: result <= 12'b101110010001;
   14853: result <= 12'b101110010001;
   14854: result <= 12'b101110010010;
   14855: result <= 12'b101110010011;
   14856: result <= 12'b101110010011;
   14857: result <= 12'b101110010100;
   14858: result <= 12'b101110010101;
   14859: result <= 12'b101110010101;
   14860: result <= 12'b101110010110;
   14861: result <= 12'b101110010111;
   14862: result <= 12'b101110010111;
   14863: result <= 12'b101110011000;
   14864: result <= 12'b101110011001;
   14865: result <= 12'b101110011001;
   14866: result <= 12'b101110011010;
   14867: result <= 12'b101110011011;
   14868: result <= 12'b101110011011;
   14869: result <= 12'b101110011100;
   14870: result <= 12'b101110011101;
   14871: result <= 12'b101110011101;
   14872: result <= 12'b101110011110;
   14873: result <= 12'b101110011111;
   14874: result <= 12'b101110011111;
   14875: result <= 12'b101110100000;
   14876: result <= 12'b101110100001;
   14877: result <= 12'b101110100001;
   14878: result <= 12'b101110100010;
   14879: result <= 12'b101110100011;
   14880: result <= 12'b101110100011;
   14881: result <= 12'b101110100100;
   14882: result <= 12'b101110100100;
   14883: result <= 12'b101110100101;
   14884: result <= 12'b101110100110;
   14885: result <= 12'b101110100110;
   14886: result <= 12'b101110100111;
   14887: result <= 12'b101110101000;
   14888: result <= 12'b101110101000;
   14889: result <= 12'b101110101001;
   14890: result <= 12'b101110101010;
   14891: result <= 12'b101110101010;
   14892: result <= 12'b101110101011;
   14893: result <= 12'b101110101100;
   14894: result <= 12'b101110101100;
   14895: result <= 12'b101110101101;
   14896: result <= 12'b101110101110;
   14897: result <= 12'b101110101110;
   14898: result <= 12'b101110101111;
   14899: result <= 12'b101110110000;
   14900: result <= 12'b101110110000;
   14901: result <= 12'b101110110001;
   14902: result <= 12'b101110110010;
   14903: result <= 12'b101110110010;
   14904: result <= 12'b101110110011;
   14905: result <= 12'b101110110100;
   14906: result <= 12'b101110110100;
   14907: result <= 12'b101110110101;
   14908: result <= 12'b101110110110;
   14909: result <= 12'b101110110110;
   14910: result <= 12'b101110110111;
   14911: result <= 12'b101110111000;
   14912: result <= 12'b101110111000;
   14913: result <= 12'b101110111001;
   14914: result <= 12'b101110111010;
   14915: result <= 12'b101110111010;
   14916: result <= 12'b101110111011;
   14917: result <= 12'b101110111100;
   14918: result <= 12'b101110111100;
   14919: result <= 12'b101110111101;
   14920: result <= 12'b101110111110;
   14921: result <= 12'b101110111110;
   14922: result <= 12'b101110111111;
   14923: result <= 12'b101111000000;
   14924: result <= 12'b101111000000;
   14925: result <= 12'b101111000001;
   14926: result <= 12'b101111000010;
   14927: result <= 12'b101111000010;
   14928: result <= 12'b101111000011;
   14929: result <= 12'b101111000100;
   14930: result <= 12'b101111000100;
   14931: result <= 12'b101111000101;
   14932: result <= 12'b101111000110;
   14933: result <= 12'b101111000110;
   14934: result <= 12'b101111000111;
   14935: result <= 12'b101111001000;
   14936: result <= 12'b101111001000;
   14937: result <= 12'b101111001001;
   14938: result <= 12'b101111001010;
   14939: result <= 12'b101111001010;
   14940: result <= 12'b101111001011;
   14941: result <= 12'b101111001100;
   14942: result <= 12'b101111001100;
   14943: result <= 12'b101111001101;
   14944: result <= 12'b101111001110;
   14945: result <= 12'b101111001110;
   14946: result <= 12'b101111001111;
   14947: result <= 12'b101111010000;
   14948: result <= 12'b101111010000;
   14949: result <= 12'b101111010001;
   14950: result <= 12'b101111010010;
   14951: result <= 12'b101111010010;
   14952: result <= 12'b101111010011;
   14953: result <= 12'b101111010100;
   14954: result <= 12'b101111010100;
   14955: result <= 12'b101111010101;
   14956: result <= 12'b101111010110;
   14957: result <= 12'b101111010110;
   14958: result <= 12'b101111010111;
   14959: result <= 12'b101111011000;
   14960: result <= 12'b101111011000;
   14961: result <= 12'b101111011001;
   14962: result <= 12'b101111011010;
   14963: result <= 12'b101111011010;
   14964: result <= 12'b101111011011;
   14965: result <= 12'b101111011100;
   14966: result <= 12'b101111011100;
   14967: result <= 12'b101111011101;
   14968: result <= 12'b101111011110;
   14969: result <= 12'b101111011110;
   14970: result <= 12'b101111011111;
   14971: result <= 12'b101111100000;
   14972: result <= 12'b101111100000;
   14973: result <= 12'b101111100001;
   14974: result <= 12'b101111100010;
   14975: result <= 12'b101111100010;
   14976: result <= 12'b101111100011;
   14977: result <= 12'b101111100100;
   14978: result <= 12'b101111100100;
   14979: result <= 12'b101111100101;
   14980: result <= 12'b101111100110;
   14981: result <= 12'b101111100110;
   14982: result <= 12'b101111100111;
   14983: result <= 12'b101111101000;
   14984: result <= 12'b101111101001;
   14985: result <= 12'b101111101001;
   14986: result <= 12'b101111101010;
   14987: result <= 12'b101111101011;
   14988: result <= 12'b101111101011;
   14989: result <= 12'b101111101100;
   14990: result <= 12'b101111101101;
   14991: result <= 12'b101111101101;
   14992: result <= 12'b101111101110;
   14993: result <= 12'b101111101111;
   14994: result <= 12'b101111101111;
   14995: result <= 12'b101111110000;
   14996: result <= 12'b101111110001;
   14997: result <= 12'b101111110001;
   14998: result <= 12'b101111110010;
   14999: result <= 12'b101111110011;
   15000: result <= 12'b101111110011;
   15001: result <= 12'b101111110100;
   15002: result <= 12'b101111110101;
   15003: result <= 12'b101111110101;
   15004: result <= 12'b101111110110;
   15005: result <= 12'b101111110111;
   15006: result <= 12'b101111110111;
   15007: result <= 12'b101111111000;
   15008: result <= 12'b101111111001;
   15009: result <= 12'b101111111001;
   15010: result <= 12'b101111111010;
   15011: result <= 12'b101111111011;
   15012: result <= 12'b101111111011;
   15013: result <= 12'b101111111100;
   15014: result <= 12'b101111111101;
   15015: result <= 12'b101111111110;
   15016: result <= 12'b101111111110;
   15017: result <= 12'b101111111111;
   15018: result <= 12'b110000000000;
   15019: result <= 12'b110000000000;
   15020: result <= 12'b110000000001;
   15021: result <= 12'b110000000010;
   15022: result <= 12'b110000000010;
   15023: result <= 12'b110000000011;
   15024: result <= 12'b110000000100;
   15025: result <= 12'b110000000100;
   15026: result <= 12'b110000000101;
   15027: result <= 12'b110000000110;
   15028: result <= 12'b110000000110;
   15029: result <= 12'b110000000111;
   15030: result <= 12'b110000001000;
   15031: result <= 12'b110000001000;
   15032: result <= 12'b110000001001;
   15033: result <= 12'b110000001010;
   15034: result <= 12'b110000001010;
   15035: result <= 12'b110000001011;
   15036: result <= 12'b110000001100;
   15037: result <= 12'b110000001100;
   15038: result <= 12'b110000001101;
   15039: result <= 12'b110000001110;
   15040: result <= 12'b110000001111;
   15041: result <= 12'b110000001111;
   15042: result <= 12'b110000010000;
   15043: result <= 12'b110000010001;
   15044: result <= 12'b110000010001;
   15045: result <= 12'b110000010010;
   15046: result <= 12'b110000010011;
   15047: result <= 12'b110000010011;
   15048: result <= 12'b110000010100;
   15049: result <= 12'b110000010101;
   15050: result <= 12'b110000010101;
   15051: result <= 12'b110000010110;
   15052: result <= 12'b110000010111;
   15053: result <= 12'b110000010111;
   15054: result <= 12'b110000011000;
   15055: result <= 12'b110000011001;
   15056: result <= 12'b110000011001;
   15057: result <= 12'b110000011010;
   15058: result <= 12'b110000011011;
   15059: result <= 12'b110000011100;
   15060: result <= 12'b110000011100;
   15061: result <= 12'b110000011101;
   15062: result <= 12'b110000011110;
   15063: result <= 12'b110000011110;
   15064: result <= 12'b110000011111;
   15065: result <= 12'b110000100000;
   15066: result <= 12'b110000100000;
   15067: result <= 12'b110000100001;
   15068: result <= 12'b110000100010;
   15069: result <= 12'b110000100010;
   15070: result <= 12'b110000100011;
   15071: result <= 12'b110000100100;
   15072: result <= 12'b110000100100;
   15073: result <= 12'b110000100101;
   15074: result <= 12'b110000100110;
   15075: result <= 12'b110000100111;
   15076: result <= 12'b110000100111;
   15077: result <= 12'b110000101000;
   15078: result <= 12'b110000101001;
   15079: result <= 12'b110000101001;
   15080: result <= 12'b110000101010;
   15081: result <= 12'b110000101011;
   15082: result <= 12'b110000101011;
   15083: result <= 12'b110000101100;
   15084: result <= 12'b110000101101;
   15085: result <= 12'b110000101101;
   15086: result <= 12'b110000101110;
   15087: result <= 12'b110000101111;
   15088: result <= 12'b110000110000;
   15089: result <= 12'b110000110000;
   15090: result <= 12'b110000110001;
   15091: result <= 12'b110000110010;
   15092: result <= 12'b110000110010;
   15093: result <= 12'b110000110011;
   15094: result <= 12'b110000110100;
   15095: result <= 12'b110000110100;
   15096: result <= 12'b110000110101;
   15097: result <= 12'b110000110110;
   15098: result <= 12'b110000110110;
   15099: result <= 12'b110000110111;
   15100: result <= 12'b110000111000;
   15101: result <= 12'b110000111001;
   15102: result <= 12'b110000111001;
   15103: result <= 12'b110000111010;
   15104: result <= 12'b110000111011;
   15105: result <= 12'b110000111011;
   15106: result <= 12'b110000111100;
   15107: result <= 12'b110000111101;
   15108: result <= 12'b110000111101;
   15109: result <= 12'b110000111110;
   15110: result <= 12'b110000111111;
   15111: result <= 12'b110000111111;
   15112: result <= 12'b110001000000;
   15113: result <= 12'b110001000001;
   15114: result <= 12'b110001000010;
   15115: result <= 12'b110001000010;
   15116: result <= 12'b110001000011;
   15117: result <= 12'b110001000100;
   15118: result <= 12'b110001000100;
   15119: result <= 12'b110001000101;
   15120: result <= 12'b110001000110;
   15121: result <= 12'b110001000110;
   15122: result <= 12'b110001000111;
   15123: result <= 12'b110001001000;
   15124: result <= 12'b110001001000;
   15125: result <= 12'b110001001001;
   15126: result <= 12'b110001001010;
   15127: result <= 12'b110001001011;
   15128: result <= 12'b110001001011;
   15129: result <= 12'b110001001100;
   15130: result <= 12'b110001001101;
   15131: result <= 12'b110001001101;
   15132: result <= 12'b110001001110;
   15133: result <= 12'b110001001111;
   15134: result <= 12'b110001001111;
   15135: result <= 12'b110001010000;
   15136: result <= 12'b110001010001;
   15137: result <= 12'b110001010010;
   15138: result <= 12'b110001010010;
   15139: result <= 12'b110001010011;
   15140: result <= 12'b110001010100;
   15141: result <= 12'b110001010100;
   15142: result <= 12'b110001010101;
   15143: result <= 12'b110001010110;
   15144: result <= 12'b110001010110;
   15145: result <= 12'b110001010111;
   15146: result <= 12'b110001011000;
   15147: result <= 12'b110001011000;
   15148: result <= 12'b110001011001;
   15149: result <= 12'b110001011010;
   15150: result <= 12'b110001011011;
   15151: result <= 12'b110001011011;
   15152: result <= 12'b110001011100;
   15153: result <= 12'b110001011101;
   15154: result <= 12'b110001011101;
   15155: result <= 12'b110001011110;
   15156: result <= 12'b110001011111;
   15157: result <= 12'b110001011111;
   15158: result <= 12'b110001100000;
   15159: result <= 12'b110001100001;
   15160: result <= 12'b110001100010;
   15161: result <= 12'b110001100010;
   15162: result <= 12'b110001100011;
   15163: result <= 12'b110001100100;
   15164: result <= 12'b110001100100;
   15165: result <= 12'b110001100101;
   15166: result <= 12'b110001100110;
   15167: result <= 12'b110001100110;
   15168: result <= 12'b110001100111;
   15169: result <= 12'b110001101000;
   15170: result <= 12'b110001101001;
   15171: result <= 12'b110001101001;
   15172: result <= 12'b110001101010;
   15173: result <= 12'b110001101011;
   15174: result <= 12'b110001101011;
   15175: result <= 12'b110001101100;
   15176: result <= 12'b110001101101;
   15177: result <= 12'b110001101110;
   15178: result <= 12'b110001101110;
   15179: result <= 12'b110001101111;
   15180: result <= 12'b110001110000;
   15181: result <= 12'b110001110000;
   15182: result <= 12'b110001110001;
   15183: result <= 12'b110001110010;
   15184: result <= 12'b110001110010;
   15185: result <= 12'b110001110011;
   15186: result <= 12'b110001110100;
   15187: result <= 12'b110001110101;
   15188: result <= 12'b110001110101;
   15189: result <= 12'b110001110110;
   15190: result <= 12'b110001110111;
   15191: result <= 12'b110001110111;
   15192: result <= 12'b110001111000;
   15193: result <= 12'b110001111001;
   15194: result <= 12'b110001111001;
   15195: result <= 12'b110001111010;
   15196: result <= 12'b110001111011;
   15197: result <= 12'b110001111100;
   15198: result <= 12'b110001111100;
   15199: result <= 12'b110001111101;
   15200: result <= 12'b110001111110;
   15201: result <= 12'b110001111110;
   15202: result <= 12'b110001111111;
   15203: result <= 12'b110010000000;
   15204: result <= 12'b110010000001;
   15205: result <= 12'b110010000001;
   15206: result <= 12'b110010000010;
   15207: result <= 12'b110010000011;
   15208: result <= 12'b110010000011;
   15209: result <= 12'b110010000100;
   15210: result <= 12'b110010000101;
   15211: result <= 12'b110010000101;
   15212: result <= 12'b110010000110;
   15213: result <= 12'b110010000111;
   15214: result <= 12'b110010001000;
   15215: result <= 12'b110010001000;
   15216: result <= 12'b110010001001;
   15217: result <= 12'b110010001010;
   15218: result <= 12'b110010001010;
   15219: result <= 12'b110010001011;
   15220: result <= 12'b110010001100;
   15221: result <= 12'b110010001101;
   15222: result <= 12'b110010001101;
   15223: result <= 12'b110010001110;
   15224: result <= 12'b110010001111;
   15225: result <= 12'b110010001111;
   15226: result <= 12'b110010010000;
   15227: result <= 12'b110010010001;
   15228: result <= 12'b110010010010;
   15229: result <= 12'b110010010010;
   15230: result <= 12'b110010010011;
   15231: result <= 12'b110010010100;
   15232: result <= 12'b110010010100;
   15233: result <= 12'b110010010101;
   15234: result <= 12'b110010010110;
   15235: result <= 12'b110010010110;
   15236: result <= 12'b110010010111;
   15237: result <= 12'b110010011000;
   15238: result <= 12'b110010011001;
   15239: result <= 12'b110010011001;
   15240: result <= 12'b110010011010;
   15241: result <= 12'b110010011011;
   15242: result <= 12'b110010011011;
   15243: result <= 12'b110010011100;
   15244: result <= 12'b110010011101;
   15245: result <= 12'b110010011110;
   15246: result <= 12'b110010011110;
   15247: result <= 12'b110010011111;
   15248: result <= 12'b110010100000;
   15249: result <= 12'b110010100000;
   15250: result <= 12'b110010100001;
   15251: result <= 12'b110010100010;
   15252: result <= 12'b110010100011;
   15253: result <= 12'b110010100011;
   15254: result <= 12'b110010100100;
   15255: result <= 12'b110010100101;
   15256: result <= 12'b110010100101;
   15257: result <= 12'b110010100110;
   15258: result <= 12'b110010100111;
   15259: result <= 12'b110010101000;
   15260: result <= 12'b110010101000;
   15261: result <= 12'b110010101001;
   15262: result <= 12'b110010101010;
   15263: result <= 12'b110010101010;
   15264: result <= 12'b110010101011;
   15265: result <= 12'b110010101100;
   15266: result <= 12'b110010101101;
   15267: result <= 12'b110010101101;
   15268: result <= 12'b110010101110;
   15269: result <= 12'b110010101111;
   15270: result <= 12'b110010101111;
   15271: result <= 12'b110010110000;
   15272: result <= 12'b110010110001;
   15273: result <= 12'b110010110010;
   15274: result <= 12'b110010110010;
   15275: result <= 12'b110010110011;
   15276: result <= 12'b110010110100;
   15277: result <= 12'b110010110100;
   15278: result <= 12'b110010110101;
   15279: result <= 12'b110010110110;
   15280: result <= 12'b110010110111;
   15281: result <= 12'b110010110111;
   15282: result <= 12'b110010111000;
   15283: result <= 12'b110010111001;
   15284: result <= 12'b110010111001;
   15285: result <= 12'b110010111010;
   15286: result <= 12'b110010111011;
   15287: result <= 12'b110010111100;
   15288: result <= 12'b110010111100;
   15289: result <= 12'b110010111101;
   15290: result <= 12'b110010111110;
   15291: result <= 12'b110010111110;
   15292: result <= 12'b110010111111;
   15293: result <= 12'b110011000000;
   15294: result <= 12'b110011000001;
   15295: result <= 12'b110011000001;
   15296: result <= 12'b110011000010;
   15297: result <= 12'b110011000011;
   15298: result <= 12'b110011000100;
   15299: result <= 12'b110011000100;
   15300: result <= 12'b110011000101;
   15301: result <= 12'b110011000110;
   15302: result <= 12'b110011000110;
   15303: result <= 12'b110011000111;
   15304: result <= 12'b110011001000;
   15305: result <= 12'b110011001001;
   15306: result <= 12'b110011001001;
   15307: result <= 12'b110011001010;
   15308: result <= 12'b110011001011;
   15309: result <= 12'b110011001011;
   15310: result <= 12'b110011001100;
   15311: result <= 12'b110011001101;
   15312: result <= 12'b110011001110;
   15313: result <= 12'b110011001110;
   15314: result <= 12'b110011001111;
   15315: result <= 12'b110011010000;
   15316: result <= 12'b110011010000;
   15317: result <= 12'b110011010001;
   15318: result <= 12'b110011010010;
   15319: result <= 12'b110011010011;
   15320: result <= 12'b110011010011;
   15321: result <= 12'b110011010100;
   15322: result <= 12'b110011010101;
   15323: result <= 12'b110011010101;
   15324: result <= 12'b110011010110;
   15325: result <= 12'b110011010111;
   15326: result <= 12'b110011011000;
   15327: result <= 12'b110011011000;
   15328: result <= 12'b110011011001;
   15329: result <= 12'b110011011010;
   15330: result <= 12'b110011011011;
   15331: result <= 12'b110011011011;
   15332: result <= 12'b110011011100;
   15333: result <= 12'b110011011101;
   15334: result <= 12'b110011011101;
   15335: result <= 12'b110011011110;
   15336: result <= 12'b110011011111;
   15337: result <= 12'b110011100000;
   15338: result <= 12'b110011100000;
   15339: result <= 12'b110011100001;
   15340: result <= 12'b110011100010;
   15341: result <= 12'b110011100010;
   15342: result <= 12'b110011100011;
   15343: result <= 12'b110011100100;
   15344: result <= 12'b110011100101;
   15345: result <= 12'b110011100101;
   15346: result <= 12'b110011100110;
   15347: result <= 12'b110011100111;
   15348: result <= 12'b110011101000;
   15349: result <= 12'b110011101000;
   15350: result <= 12'b110011101001;
   15351: result <= 12'b110011101010;
   15352: result <= 12'b110011101010;
   15353: result <= 12'b110011101011;
   15354: result <= 12'b110011101100;
   15355: result <= 12'b110011101101;
   15356: result <= 12'b110011101101;
   15357: result <= 12'b110011101110;
   15358: result <= 12'b110011101111;
   15359: result <= 12'b110011110000;
   15360: result <= 12'b110011110000;
   15361: result <= 12'b110011110001;
   15362: result <= 12'b110011110010;
   15363: result <= 12'b110011110010;
   15364: result <= 12'b110011110011;
   15365: result <= 12'b110011110100;
   15366: result <= 12'b110011110101;
   15367: result <= 12'b110011110101;
   15368: result <= 12'b110011110110;
   15369: result <= 12'b110011110111;
   15370: result <= 12'b110011111000;
   15371: result <= 12'b110011111000;
   15372: result <= 12'b110011111001;
   15373: result <= 12'b110011111010;
   15374: result <= 12'b110011111010;
   15375: result <= 12'b110011111011;
   15376: result <= 12'b110011111100;
   15377: result <= 12'b110011111101;
   15378: result <= 12'b110011111101;
   15379: result <= 12'b110011111110;
   15380: result <= 12'b110011111111;
   15381: result <= 12'b110100000000;
   15382: result <= 12'b110100000000;
   15383: result <= 12'b110100000001;
   15384: result <= 12'b110100000010;
   15385: result <= 12'b110100000010;
   15386: result <= 12'b110100000011;
   15387: result <= 12'b110100000100;
   15388: result <= 12'b110100000101;
   15389: result <= 12'b110100000101;
   15390: result <= 12'b110100000110;
   15391: result <= 12'b110100000111;
   15392: result <= 12'b110100001000;
   15393: result <= 12'b110100001000;
   15394: result <= 12'b110100001001;
   15395: result <= 12'b110100001010;
   15396: result <= 12'b110100001010;
   15397: result <= 12'b110100001011;
   15398: result <= 12'b110100001100;
   15399: result <= 12'b110100001101;
   15400: result <= 12'b110100001101;
   15401: result <= 12'b110100001110;
   15402: result <= 12'b110100001111;
   15403: result <= 12'b110100010000;
   15404: result <= 12'b110100010000;
   15405: result <= 12'b110100010001;
   15406: result <= 12'b110100010010;
   15407: result <= 12'b110100010010;
   15408: result <= 12'b110100010011;
   15409: result <= 12'b110100010100;
   15410: result <= 12'b110100010101;
   15411: result <= 12'b110100010101;
   15412: result <= 12'b110100010110;
   15413: result <= 12'b110100010111;
   15414: result <= 12'b110100011000;
   15415: result <= 12'b110100011000;
   15416: result <= 12'b110100011001;
   15417: result <= 12'b110100011010;
   15418: result <= 12'b110100011011;
   15419: result <= 12'b110100011011;
   15420: result <= 12'b110100011100;
   15421: result <= 12'b110100011101;
   15422: result <= 12'b110100011101;
   15423: result <= 12'b110100011110;
   15424: result <= 12'b110100011111;
   15425: result <= 12'b110100100000;
   15426: result <= 12'b110100100000;
   15427: result <= 12'b110100100001;
   15428: result <= 12'b110100100010;
   15429: result <= 12'b110100100011;
   15430: result <= 12'b110100100011;
   15431: result <= 12'b110100100100;
   15432: result <= 12'b110100100101;
   15433: result <= 12'b110100100110;
   15434: result <= 12'b110100100110;
   15435: result <= 12'b110100100111;
   15436: result <= 12'b110100101000;
   15437: result <= 12'b110100101000;
   15438: result <= 12'b110100101001;
   15439: result <= 12'b110100101010;
   15440: result <= 12'b110100101011;
   15441: result <= 12'b110100101011;
   15442: result <= 12'b110100101100;
   15443: result <= 12'b110100101101;
   15444: result <= 12'b110100101110;
   15445: result <= 12'b110100101110;
   15446: result <= 12'b110100101111;
   15447: result <= 12'b110100110000;
   15448: result <= 12'b110100110001;
   15449: result <= 12'b110100110001;
   15450: result <= 12'b110100110010;
   15451: result <= 12'b110100110011;
   15452: result <= 12'b110100110011;
   15453: result <= 12'b110100110100;
   15454: result <= 12'b110100110101;
   15455: result <= 12'b110100110110;
   15456: result <= 12'b110100110110;
   15457: result <= 12'b110100110111;
   15458: result <= 12'b110100111000;
   15459: result <= 12'b110100111001;
   15460: result <= 12'b110100111001;
   15461: result <= 12'b110100111010;
   15462: result <= 12'b110100111011;
   15463: result <= 12'b110100111100;
   15464: result <= 12'b110100111100;
   15465: result <= 12'b110100111101;
   15466: result <= 12'b110100111110;
   15467: result <= 12'b110100111111;
   15468: result <= 12'b110100111111;
   15469: result <= 12'b110101000000;
   15470: result <= 12'b110101000001;
   15471: result <= 12'b110101000001;
   15472: result <= 12'b110101000010;
   15473: result <= 12'b110101000011;
   15474: result <= 12'b110101000100;
   15475: result <= 12'b110101000100;
   15476: result <= 12'b110101000101;
   15477: result <= 12'b110101000110;
   15478: result <= 12'b110101000111;
   15479: result <= 12'b110101000111;
   15480: result <= 12'b110101001000;
   15481: result <= 12'b110101001001;
   15482: result <= 12'b110101001010;
   15483: result <= 12'b110101001010;
   15484: result <= 12'b110101001011;
   15485: result <= 12'b110101001100;
   15486: result <= 12'b110101001101;
   15487: result <= 12'b110101001101;
   15488: result <= 12'b110101001110;
   15489: result <= 12'b110101001111;
   15490: result <= 12'b110101010000;
   15491: result <= 12'b110101010000;
   15492: result <= 12'b110101010001;
   15493: result <= 12'b110101010010;
   15494: result <= 12'b110101010010;
   15495: result <= 12'b110101010011;
   15496: result <= 12'b110101010100;
   15497: result <= 12'b110101010101;
   15498: result <= 12'b110101010101;
   15499: result <= 12'b110101010110;
   15500: result <= 12'b110101010111;
   15501: result <= 12'b110101011000;
   15502: result <= 12'b110101011000;
   15503: result <= 12'b110101011001;
   15504: result <= 12'b110101011010;
   15505: result <= 12'b110101011011;
   15506: result <= 12'b110101011011;
   15507: result <= 12'b110101011100;
   15508: result <= 12'b110101011101;
   15509: result <= 12'b110101011110;
   15510: result <= 12'b110101011110;
   15511: result <= 12'b110101011111;
   15512: result <= 12'b110101100000;
   15513: result <= 12'b110101100001;
   15514: result <= 12'b110101100001;
   15515: result <= 12'b110101100010;
   15516: result <= 12'b110101100011;
   15517: result <= 12'b110101100100;
   15518: result <= 12'b110101100100;
   15519: result <= 12'b110101100101;
   15520: result <= 12'b110101100110;
   15521: result <= 12'b110101100111;
   15522: result <= 12'b110101100111;
   15523: result <= 12'b110101101000;
   15524: result <= 12'b110101101001;
   15525: result <= 12'b110101101001;
   15526: result <= 12'b110101101010;
   15527: result <= 12'b110101101011;
   15528: result <= 12'b110101101100;
   15529: result <= 12'b110101101100;
   15530: result <= 12'b110101101101;
   15531: result <= 12'b110101101110;
   15532: result <= 12'b110101101111;
   15533: result <= 12'b110101101111;
   15534: result <= 12'b110101110000;
   15535: result <= 12'b110101110001;
   15536: result <= 12'b110101110010;
   15537: result <= 12'b110101110010;
   15538: result <= 12'b110101110011;
   15539: result <= 12'b110101110100;
   15540: result <= 12'b110101110101;
   15541: result <= 12'b110101110101;
   15542: result <= 12'b110101110110;
   15543: result <= 12'b110101110111;
   15544: result <= 12'b110101111000;
   15545: result <= 12'b110101111000;
   15546: result <= 12'b110101111001;
   15547: result <= 12'b110101111010;
   15548: result <= 12'b110101111011;
   15549: result <= 12'b110101111011;
   15550: result <= 12'b110101111100;
   15551: result <= 12'b110101111101;
   15552: result <= 12'b110101111110;
   15553: result <= 12'b110101111110;
   15554: result <= 12'b110101111111;
   15555: result <= 12'b110110000000;
   15556: result <= 12'b110110000001;
   15557: result <= 12'b110110000001;
   15558: result <= 12'b110110000010;
   15559: result <= 12'b110110000011;
   15560: result <= 12'b110110000100;
   15561: result <= 12'b110110000100;
   15562: result <= 12'b110110000101;
   15563: result <= 12'b110110000110;
   15564: result <= 12'b110110000111;
   15565: result <= 12'b110110000111;
   15566: result <= 12'b110110001000;
   15567: result <= 12'b110110001001;
   15568: result <= 12'b110110001010;
   15569: result <= 12'b110110001010;
   15570: result <= 12'b110110001011;
   15571: result <= 12'b110110001100;
   15572: result <= 12'b110110001101;
   15573: result <= 12'b110110001101;
   15574: result <= 12'b110110001110;
   15575: result <= 12'b110110001111;
   15576: result <= 12'b110110010000;
   15577: result <= 12'b110110010000;
   15578: result <= 12'b110110010001;
   15579: result <= 12'b110110010010;
   15580: result <= 12'b110110010010;
   15581: result <= 12'b110110010011;
   15582: result <= 12'b110110010100;
   15583: result <= 12'b110110010101;
   15584: result <= 12'b110110010101;
   15585: result <= 12'b110110010110;
   15586: result <= 12'b110110010111;
   15587: result <= 12'b110110011000;
   15588: result <= 12'b110110011000;
   15589: result <= 12'b110110011001;
   15590: result <= 12'b110110011010;
   15591: result <= 12'b110110011011;
   15592: result <= 12'b110110011011;
   15593: result <= 12'b110110011100;
   15594: result <= 12'b110110011101;
   15595: result <= 12'b110110011110;
   15596: result <= 12'b110110011110;
   15597: result <= 12'b110110011111;
   15598: result <= 12'b110110100000;
   15599: result <= 12'b110110100001;
   15600: result <= 12'b110110100001;
   15601: result <= 12'b110110100010;
   15602: result <= 12'b110110100011;
   15603: result <= 12'b110110100100;
   15604: result <= 12'b110110100100;
   15605: result <= 12'b110110100101;
   15606: result <= 12'b110110100110;
   15607: result <= 12'b110110100111;
   15608: result <= 12'b110110100111;
   15609: result <= 12'b110110101000;
   15610: result <= 12'b110110101001;
   15611: result <= 12'b110110101010;
   15612: result <= 12'b110110101010;
   15613: result <= 12'b110110101011;
   15614: result <= 12'b110110101100;
   15615: result <= 12'b110110101101;
   15616: result <= 12'b110110101101;
   15617: result <= 12'b110110101110;
   15618: result <= 12'b110110101111;
   15619: result <= 12'b110110110000;
   15620: result <= 12'b110110110001;
   15621: result <= 12'b110110110001;
   15622: result <= 12'b110110110010;
   15623: result <= 12'b110110110011;
   15624: result <= 12'b110110110100;
   15625: result <= 12'b110110110100;
   15626: result <= 12'b110110110101;
   15627: result <= 12'b110110110110;
   15628: result <= 12'b110110110111;
   15629: result <= 12'b110110110111;
   15630: result <= 12'b110110111000;
   15631: result <= 12'b110110111001;
   15632: result <= 12'b110110111010;
   15633: result <= 12'b110110111010;
   15634: result <= 12'b110110111011;
   15635: result <= 12'b110110111100;
   15636: result <= 12'b110110111101;
   15637: result <= 12'b110110111101;
   15638: result <= 12'b110110111110;
   15639: result <= 12'b110110111111;
   15640: result <= 12'b110111000000;
   15641: result <= 12'b110111000000;
   15642: result <= 12'b110111000001;
   15643: result <= 12'b110111000010;
   15644: result <= 12'b110111000011;
   15645: result <= 12'b110111000011;
   15646: result <= 12'b110111000100;
   15647: result <= 12'b110111000101;
   15648: result <= 12'b110111000110;
   15649: result <= 12'b110111000110;
   15650: result <= 12'b110111000111;
   15651: result <= 12'b110111001000;
   15652: result <= 12'b110111001001;
   15653: result <= 12'b110111001001;
   15654: result <= 12'b110111001010;
   15655: result <= 12'b110111001011;
   15656: result <= 12'b110111001100;
   15657: result <= 12'b110111001100;
   15658: result <= 12'b110111001101;
   15659: result <= 12'b110111001110;
   15660: result <= 12'b110111001111;
   15661: result <= 12'b110111001111;
   15662: result <= 12'b110111010000;
   15663: result <= 12'b110111010001;
   15664: result <= 12'b110111010010;
   15665: result <= 12'b110111010010;
   15666: result <= 12'b110111010011;
   15667: result <= 12'b110111010100;
   15668: result <= 12'b110111010101;
   15669: result <= 12'b110111010101;
   15670: result <= 12'b110111010110;
   15671: result <= 12'b110111010111;
   15672: result <= 12'b110111011000;
   15673: result <= 12'b110111011000;
   15674: result <= 12'b110111011001;
   15675: result <= 12'b110111011010;
   15676: result <= 12'b110111011011;
   15677: result <= 12'b110111011100;
   15678: result <= 12'b110111011100;
   15679: result <= 12'b110111011101;
   15680: result <= 12'b110111011110;
   15681: result <= 12'b110111011111;
   15682: result <= 12'b110111011111;
   15683: result <= 12'b110111100000;
   15684: result <= 12'b110111100001;
   15685: result <= 12'b110111100010;
   15686: result <= 12'b110111100010;
   15687: result <= 12'b110111100011;
   15688: result <= 12'b110111100100;
   15689: result <= 12'b110111100101;
   15690: result <= 12'b110111100101;
   15691: result <= 12'b110111100110;
   15692: result <= 12'b110111100111;
   15693: result <= 12'b110111101000;
   15694: result <= 12'b110111101000;
   15695: result <= 12'b110111101001;
   15696: result <= 12'b110111101010;
   15697: result <= 12'b110111101011;
   15698: result <= 12'b110111101011;
   15699: result <= 12'b110111101100;
   15700: result <= 12'b110111101101;
   15701: result <= 12'b110111101110;
   15702: result <= 12'b110111101110;
   15703: result <= 12'b110111101111;
   15704: result <= 12'b110111110000;
   15705: result <= 12'b110111110001;
   15706: result <= 12'b110111110001;
   15707: result <= 12'b110111110010;
   15708: result <= 12'b110111110011;
   15709: result <= 12'b110111110100;
   15710: result <= 12'b110111110101;
   15711: result <= 12'b110111110101;
   15712: result <= 12'b110111110110;
   15713: result <= 12'b110111110111;
   15714: result <= 12'b110111111000;
   15715: result <= 12'b110111111000;
   15716: result <= 12'b110111111001;
   15717: result <= 12'b110111111010;
   15718: result <= 12'b110111111011;
   15719: result <= 12'b110111111011;
   15720: result <= 12'b110111111100;
   15721: result <= 12'b110111111101;
   15722: result <= 12'b110111111110;
   15723: result <= 12'b110111111110;
   15724: result <= 12'b110111111111;
   15725: result <= 12'b111000000000;
   15726: result <= 12'b111000000001;
   15727: result <= 12'b111000000001;
   15728: result <= 12'b111000000010;
   15729: result <= 12'b111000000011;
   15730: result <= 12'b111000000100;
   15731: result <= 12'b111000000100;
   15732: result <= 12'b111000000101;
   15733: result <= 12'b111000000110;
   15734: result <= 12'b111000000111;
   15735: result <= 12'b111000001000;
   15736: result <= 12'b111000001000;
   15737: result <= 12'b111000001001;
   15738: result <= 12'b111000001010;
   15739: result <= 12'b111000001011;
   15740: result <= 12'b111000001011;
   15741: result <= 12'b111000001100;
   15742: result <= 12'b111000001101;
   15743: result <= 12'b111000001110;
   15744: result <= 12'b111000001110;
   15745: result <= 12'b111000001111;
   15746: result <= 12'b111000010000;
   15747: result <= 12'b111000010001;
   15748: result <= 12'b111000010001;
   15749: result <= 12'b111000010010;
   15750: result <= 12'b111000010011;
   15751: result <= 12'b111000010100;
   15752: result <= 12'b111000010100;
   15753: result <= 12'b111000010101;
   15754: result <= 12'b111000010110;
   15755: result <= 12'b111000010111;
   15756: result <= 12'b111000011000;
   15757: result <= 12'b111000011000;
   15758: result <= 12'b111000011001;
   15759: result <= 12'b111000011010;
   15760: result <= 12'b111000011011;
   15761: result <= 12'b111000011011;
   15762: result <= 12'b111000011100;
   15763: result <= 12'b111000011101;
   15764: result <= 12'b111000011110;
   15765: result <= 12'b111000011110;
   15766: result <= 12'b111000011111;
   15767: result <= 12'b111000100000;
   15768: result <= 12'b111000100001;
   15769: result <= 12'b111000100001;
   15770: result <= 12'b111000100010;
   15771: result <= 12'b111000100011;
   15772: result <= 12'b111000100100;
   15773: result <= 12'b111000100101;
   15774: result <= 12'b111000100101;
   15775: result <= 12'b111000100110;
   15776: result <= 12'b111000100111;
   15777: result <= 12'b111000101000;
   15778: result <= 12'b111000101000;
   15779: result <= 12'b111000101001;
   15780: result <= 12'b111000101010;
   15781: result <= 12'b111000101011;
   15782: result <= 12'b111000101011;
   15783: result <= 12'b111000101100;
   15784: result <= 12'b111000101101;
   15785: result <= 12'b111000101110;
   15786: result <= 12'b111000101110;
   15787: result <= 12'b111000101111;
   15788: result <= 12'b111000110000;
   15789: result <= 12'b111000110001;
   15790: result <= 12'b111000110001;
   15791: result <= 12'b111000110010;
   15792: result <= 12'b111000110011;
   15793: result <= 12'b111000110100;
   15794: result <= 12'b111000110101;
   15795: result <= 12'b111000110101;
   15796: result <= 12'b111000110110;
   15797: result <= 12'b111000110111;
   15798: result <= 12'b111000111000;
   15799: result <= 12'b111000111000;
   15800: result <= 12'b111000111001;
   15801: result <= 12'b111000111010;
   15802: result <= 12'b111000111011;
   15803: result <= 12'b111000111011;
   15804: result <= 12'b111000111100;
   15805: result <= 12'b111000111101;
   15806: result <= 12'b111000111110;
   15807: result <= 12'b111000111111;
   15808: result <= 12'b111000111111;
   15809: result <= 12'b111001000000;
   15810: result <= 12'b111001000001;
   15811: result <= 12'b111001000010;
   15812: result <= 12'b111001000010;
   15813: result <= 12'b111001000011;
   15814: result <= 12'b111001000100;
   15815: result <= 12'b111001000101;
   15816: result <= 12'b111001000101;
   15817: result <= 12'b111001000110;
   15818: result <= 12'b111001000111;
   15819: result <= 12'b111001001000;
   15820: result <= 12'b111001001000;
   15821: result <= 12'b111001001001;
   15822: result <= 12'b111001001010;
   15823: result <= 12'b111001001011;
   15824: result <= 12'b111001001100;
   15825: result <= 12'b111001001100;
   15826: result <= 12'b111001001101;
   15827: result <= 12'b111001001110;
   15828: result <= 12'b111001001111;
   15829: result <= 12'b111001001111;
   15830: result <= 12'b111001010000;
   15831: result <= 12'b111001010001;
   15832: result <= 12'b111001010010;
   15833: result <= 12'b111001010010;
   15834: result <= 12'b111001010011;
   15835: result <= 12'b111001010100;
   15836: result <= 12'b111001010101;
   15837: result <= 12'b111001010110;
   15838: result <= 12'b111001010110;
   15839: result <= 12'b111001010111;
   15840: result <= 12'b111001011000;
   15841: result <= 12'b111001011001;
   15842: result <= 12'b111001011001;
   15843: result <= 12'b111001011010;
   15844: result <= 12'b111001011011;
   15845: result <= 12'b111001011100;
   15846: result <= 12'b111001011100;
   15847: result <= 12'b111001011101;
   15848: result <= 12'b111001011110;
   15849: result <= 12'b111001011111;
   15850: result <= 12'b111001100000;
   15851: result <= 12'b111001100000;
   15852: result <= 12'b111001100001;
   15853: result <= 12'b111001100010;
   15854: result <= 12'b111001100011;
   15855: result <= 12'b111001100011;
   15856: result <= 12'b111001100100;
   15857: result <= 12'b111001100101;
   15858: result <= 12'b111001100110;
   15859: result <= 12'b111001100110;
   15860: result <= 12'b111001100111;
   15861: result <= 12'b111001101000;
   15862: result <= 12'b111001101001;
   15863: result <= 12'b111001101010;
   15864: result <= 12'b111001101010;
   15865: result <= 12'b111001101011;
   15866: result <= 12'b111001101100;
   15867: result <= 12'b111001101101;
   15868: result <= 12'b111001101101;
   15869: result <= 12'b111001101110;
   15870: result <= 12'b111001101111;
   15871: result <= 12'b111001110000;
   15872: result <= 12'b111001110000;
   15873: result <= 12'b111001110001;
   15874: result <= 12'b111001110010;
   15875: result <= 12'b111001110011;
   15876: result <= 12'b111001110100;
   15877: result <= 12'b111001110100;
   15878: result <= 12'b111001110101;
   15879: result <= 12'b111001110110;
   15880: result <= 12'b111001110111;
   15881: result <= 12'b111001110111;
   15882: result <= 12'b111001111000;
   15883: result <= 12'b111001111001;
   15884: result <= 12'b111001111010;
   15885: result <= 12'b111001111010;
   15886: result <= 12'b111001111011;
   15887: result <= 12'b111001111100;
   15888: result <= 12'b111001111101;
   15889: result <= 12'b111001111110;
   15890: result <= 12'b111001111110;
   15891: result <= 12'b111001111111;
   15892: result <= 12'b111010000000;
   15893: result <= 12'b111010000001;
   15894: result <= 12'b111010000001;
   15895: result <= 12'b111010000010;
   15896: result <= 12'b111010000011;
   15897: result <= 12'b111010000100;
   15898: result <= 12'b111010000101;
   15899: result <= 12'b111010000101;
   15900: result <= 12'b111010000110;
   15901: result <= 12'b111010000111;
   15902: result <= 12'b111010001000;
   15903: result <= 12'b111010001000;
   15904: result <= 12'b111010001001;
   15905: result <= 12'b111010001010;
   15906: result <= 12'b111010001011;
   15907: result <= 12'b111010001011;
   15908: result <= 12'b111010001100;
   15909: result <= 12'b111010001101;
   15910: result <= 12'b111010001110;
   15911: result <= 12'b111010001111;
   15912: result <= 12'b111010001111;
   15913: result <= 12'b111010010000;
   15914: result <= 12'b111010010001;
   15915: result <= 12'b111010010010;
   15916: result <= 12'b111010010010;
   15917: result <= 12'b111010010011;
   15918: result <= 12'b111010010100;
   15919: result <= 12'b111010010101;
   15920: result <= 12'b111010010101;
   15921: result <= 12'b111010010110;
   15922: result <= 12'b111010010111;
   15923: result <= 12'b111010011000;
   15924: result <= 12'b111010011001;
   15925: result <= 12'b111010011001;
   15926: result <= 12'b111010011010;
   15927: result <= 12'b111010011011;
   15928: result <= 12'b111010011100;
   15929: result <= 12'b111010011100;
   15930: result <= 12'b111010011101;
   15931: result <= 12'b111010011110;
   15932: result <= 12'b111010011111;
   15933: result <= 12'b111010100000;
   15934: result <= 12'b111010100000;
   15935: result <= 12'b111010100001;
   15936: result <= 12'b111010100010;
   15937: result <= 12'b111010100011;
   15938: result <= 12'b111010100011;
   15939: result <= 12'b111010100100;
   15940: result <= 12'b111010100101;
   15941: result <= 12'b111010100110;
   15942: result <= 12'b111010100111;
   15943: result <= 12'b111010100111;
   15944: result <= 12'b111010101000;
   15945: result <= 12'b111010101001;
   15946: result <= 12'b111010101010;
   15947: result <= 12'b111010101010;
   15948: result <= 12'b111010101011;
   15949: result <= 12'b111010101100;
   15950: result <= 12'b111010101101;
   15951: result <= 12'b111010101101;
   15952: result <= 12'b111010101110;
   15953: result <= 12'b111010101111;
   15954: result <= 12'b111010110000;
   15955: result <= 12'b111010110001;
   15956: result <= 12'b111010110001;
   15957: result <= 12'b111010110010;
   15958: result <= 12'b111010110011;
   15959: result <= 12'b111010110100;
   15960: result <= 12'b111010110100;
   15961: result <= 12'b111010110101;
   15962: result <= 12'b111010110110;
   15963: result <= 12'b111010110111;
   15964: result <= 12'b111010111000;
   15965: result <= 12'b111010111000;
   15966: result <= 12'b111010111001;
   15967: result <= 12'b111010111010;
   15968: result <= 12'b111010111011;
   15969: result <= 12'b111010111011;
   15970: result <= 12'b111010111100;
   15971: result <= 12'b111010111101;
   15972: result <= 12'b111010111110;
   15973: result <= 12'b111010111111;
   15974: result <= 12'b111010111111;
   15975: result <= 12'b111011000000;
   15976: result <= 12'b111011000001;
   15977: result <= 12'b111011000010;
   15978: result <= 12'b111011000010;
   15979: result <= 12'b111011000011;
   15980: result <= 12'b111011000100;
   15981: result <= 12'b111011000101;
   15982: result <= 12'b111011000110;
   15983: result <= 12'b111011000110;
   15984: result <= 12'b111011000111;
   15985: result <= 12'b111011001000;
   15986: result <= 12'b111011001001;
   15987: result <= 12'b111011001001;
   15988: result <= 12'b111011001010;
   15989: result <= 12'b111011001011;
   15990: result <= 12'b111011001100;
   15991: result <= 12'b111011001101;
   15992: result <= 12'b111011001101;
   15993: result <= 12'b111011001110;
   15994: result <= 12'b111011001111;
   15995: result <= 12'b111011010000;
   15996: result <= 12'b111011010000;
   15997: result <= 12'b111011010001;
   15998: result <= 12'b111011010010;
   15999: result <= 12'b111011010011;
   16000: result <= 12'b111011010011;
   16001: result <= 12'b111011010100;
   16002: result <= 12'b111011010101;
   16003: result <= 12'b111011010110;
   16004: result <= 12'b111011010111;
   16005: result <= 12'b111011010111;
   16006: result <= 12'b111011011000;
   16007: result <= 12'b111011011001;
   16008: result <= 12'b111011011010;
   16009: result <= 12'b111011011010;
   16010: result <= 12'b111011011011;
   16011: result <= 12'b111011011100;
   16012: result <= 12'b111011011101;
   16013: result <= 12'b111011011110;
   16014: result <= 12'b111011011110;
   16015: result <= 12'b111011011111;
   16016: result <= 12'b111011100000;
   16017: result <= 12'b111011100001;
   16018: result <= 12'b111011100001;
   16019: result <= 12'b111011100010;
   16020: result <= 12'b111011100011;
   16021: result <= 12'b111011100100;
   16022: result <= 12'b111011100101;
   16023: result <= 12'b111011100101;
   16024: result <= 12'b111011100110;
   16025: result <= 12'b111011100111;
   16026: result <= 12'b111011101000;
   16027: result <= 12'b111011101000;
   16028: result <= 12'b111011101001;
   16029: result <= 12'b111011101010;
   16030: result <= 12'b111011101011;
   16031: result <= 12'b111011101100;
   16032: result <= 12'b111011101100;
   16033: result <= 12'b111011101101;
   16034: result <= 12'b111011101110;
   16035: result <= 12'b111011101111;
   16036: result <= 12'b111011101111;
   16037: result <= 12'b111011110000;
   16038: result <= 12'b111011110001;
   16039: result <= 12'b111011110010;
   16040: result <= 12'b111011110011;
   16041: result <= 12'b111011110011;
   16042: result <= 12'b111011110100;
   16043: result <= 12'b111011110101;
   16044: result <= 12'b111011110110;
   16045: result <= 12'b111011110110;
   16046: result <= 12'b111011110111;
   16047: result <= 12'b111011111000;
   16048: result <= 12'b111011111001;
   16049: result <= 12'b111011111010;
   16050: result <= 12'b111011111010;
   16051: result <= 12'b111011111011;
   16052: result <= 12'b111011111100;
   16053: result <= 12'b111011111101;
   16054: result <= 12'b111011111110;
   16055: result <= 12'b111011111110;
   16056: result <= 12'b111011111111;
   16057: result <= 12'b111100000000;
   16058: result <= 12'b111100000001;
   16059: result <= 12'b111100000001;
   16060: result <= 12'b111100000010;
   16061: result <= 12'b111100000011;
   16062: result <= 12'b111100000100;
   16063: result <= 12'b111100000101;
   16064: result <= 12'b111100000101;
   16065: result <= 12'b111100000110;
   16066: result <= 12'b111100000111;
   16067: result <= 12'b111100001000;
   16068: result <= 12'b111100001000;
   16069: result <= 12'b111100001001;
   16070: result <= 12'b111100001010;
   16071: result <= 12'b111100001011;
   16072: result <= 12'b111100001100;
   16073: result <= 12'b111100001100;
   16074: result <= 12'b111100001101;
   16075: result <= 12'b111100001110;
   16076: result <= 12'b111100001111;
   16077: result <= 12'b111100001111;
   16078: result <= 12'b111100010000;
   16079: result <= 12'b111100010001;
   16080: result <= 12'b111100010010;
   16081: result <= 12'b111100010011;
   16082: result <= 12'b111100010011;
   16083: result <= 12'b111100010100;
   16084: result <= 12'b111100010101;
   16085: result <= 12'b111100010110;
   16086: result <= 12'b111100010110;
   16087: result <= 12'b111100010111;
   16088: result <= 12'b111100011000;
   16089: result <= 12'b111100011001;
   16090: result <= 12'b111100011010;
   16091: result <= 12'b111100011010;
   16092: result <= 12'b111100011011;
   16093: result <= 12'b111100011100;
   16094: result <= 12'b111100011101;
   16095: result <= 12'b111100011101;
   16096: result <= 12'b111100011110;
   16097: result <= 12'b111100011111;
   16098: result <= 12'b111100100000;
   16099: result <= 12'b111100100001;
   16100: result <= 12'b111100100001;
   16101: result <= 12'b111100100010;
   16102: result <= 12'b111100100011;
   16103: result <= 12'b111100100100;
   16104: result <= 12'b111100100101;
   16105: result <= 12'b111100100101;
   16106: result <= 12'b111100100110;
   16107: result <= 12'b111100100111;
   16108: result <= 12'b111100101000;
   16109: result <= 12'b111100101000;
   16110: result <= 12'b111100101001;
   16111: result <= 12'b111100101010;
   16112: result <= 12'b111100101011;
   16113: result <= 12'b111100101100;
   16114: result <= 12'b111100101100;
   16115: result <= 12'b111100101101;
   16116: result <= 12'b111100101110;
   16117: result <= 12'b111100101111;
   16118: result <= 12'b111100101111;
   16119: result <= 12'b111100110000;
   16120: result <= 12'b111100110001;
   16121: result <= 12'b111100110010;
   16122: result <= 12'b111100110011;
   16123: result <= 12'b111100110011;
   16124: result <= 12'b111100110100;
   16125: result <= 12'b111100110101;
   16126: result <= 12'b111100110110;
   16127: result <= 12'b111100110110;
   16128: result <= 12'b111100110111;
   16129: result <= 12'b111100111000;
   16130: result <= 12'b111100111001;
   16131: result <= 12'b111100111010;
   16132: result <= 12'b111100111010;
   16133: result <= 12'b111100111011;
   16134: result <= 12'b111100111100;
   16135: result <= 12'b111100111101;
   16136: result <= 12'b111100111110;
   16137: result <= 12'b111100111110;
   16138: result <= 12'b111100111111;
   16139: result <= 12'b111101000000;
   16140: result <= 12'b111101000001;
   16141: result <= 12'b111101000001;
   16142: result <= 12'b111101000010;
   16143: result <= 12'b111101000011;
   16144: result <= 12'b111101000100;
   16145: result <= 12'b111101000101;
   16146: result <= 12'b111101000101;
   16147: result <= 12'b111101000110;
   16148: result <= 12'b111101000111;
   16149: result <= 12'b111101001000;
   16150: result <= 12'b111101001000;
   16151: result <= 12'b111101001001;
   16152: result <= 12'b111101001010;
   16153: result <= 12'b111101001011;
   16154: result <= 12'b111101001100;
   16155: result <= 12'b111101001100;
   16156: result <= 12'b111101001101;
   16157: result <= 12'b111101001110;
   16158: result <= 12'b111101001111;
   16159: result <= 12'b111101010000;
   16160: result <= 12'b111101010000;
   16161: result <= 12'b111101010001;
   16162: result <= 12'b111101010010;
   16163: result <= 12'b111101010011;
   16164: result <= 12'b111101010011;
   16165: result <= 12'b111101010100;
   16166: result <= 12'b111101010101;
   16167: result <= 12'b111101010110;
   16168: result <= 12'b111101010111;
   16169: result <= 12'b111101010111;
   16170: result <= 12'b111101011000;
   16171: result <= 12'b111101011001;
   16172: result <= 12'b111101011010;
   16173: result <= 12'b111101011010;
   16174: result <= 12'b111101011011;
   16175: result <= 12'b111101011100;
   16176: result <= 12'b111101011101;
   16177: result <= 12'b111101011110;
   16178: result <= 12'b111101011110;
   16179: result <= 12'b111101011111;
   16180: result <= 12'b111101100000;
   16181: result <= 12'b111101100001;
   16182: result <= 12'b111101100010;
   16183: result <= 12'b111101100010;
   16184: result <= 12'b111101100011;
   16185: result <= 12'b111101100100;
   16186: result <= 12'b111101100101;
   16187: result <= 12'b111101100101;
   16188: result <= 12'b111101100110;
   16189: result <= 12'b111101100111;
   16190: result <= 12'b111101101000;
   16191: result <= 12'b111101101001;
   16192: result <= 12'b111101101001;
   16193: result <= 12'b111101101010;
   16194: result <= 12'b111101101011;
   16195: result <= 12'b111101101100;
   16196: result <= 12'b111101101100;
   16197: result <= 12'b111101101101;
   16198: result <= 12'b111101101110;
   16199: result <= 12'b111101101111;
   16200: result <= 12'b111101110000;
   16201: result <= 12'b111101110000;
   16202: result <= 12'b111101110001;
   16203: result <= 12'b111101110010;
   16204: result <= 12'b111101110011;
   16205: result <= 12'b111101110100;
   16206: result <= 12'b111101110100;
   16207: result <= 12'b111101110101;
   16208: result <= 12'b111101110110;
   16209: result <= 12'b111101110111;
   16210: result <= 12'b111101110111;
   16211: result <= 12'b111101111000;
   16212: result <= 12'b111101111001;
   16213: result <= 12'b111101111010;
   16214: result <= 12'b111101111011;
   16215: result <= 12'b111101111011;
   16216: result <= 12'b111101111100;
   16217: result <= 12'b111101111101;
   16218: result <= 12'b111101111110;
   16219: result <= 12'b111101111110;
   16220: result <= 12'b111101111111;
   16221: result <= 12'b111110000000;
   16222: result <= 12'b111110000001;
   16223: result <= 12'b111110000010;
   16224: result <= 12'b111110000010;
   16225: result <= 12'b111110000011;
   16226: result <= 12'b111110000100;
   16227: result <= 12'b111110000101;
   16228: result <= 12'b111110000110;
   16229: result <= 12'b111110000110;
   16230: result <= 12'b111110000111;
   16231: result <= 12'b111110001000;
   16232: result <= 12'b111110001001;
   16233: result <= 12'b111110001001;
   16234: result <= 12'b111110001010;
   16235: result <= 12'b111110001011;
   16236: result <= 12'b111110001100;
   16237: result <= 12'b111110001101;
   16238: result <= 12'b111110001101;
   16239: result <= 12'b111110001110;
   16240: result <= 12'b111110001111;
   16241: result <= 12'b111110010000;
   16242: result <= 12'b111110010001;
   16243: result <= 12'b111110010001;
   16244: result <= 12'b111110010010;
   16245: result <= 12'b111110010011;
   16246: result <= 12'b111110010100;
   16247: result <= 12'b111110010100;
   16248: result <= 12'b111110010101;
   16249: result <= 12'b111110010110;
   16250: result <= 12'b111110010111;
   16251: result <= 12'b111110011000;
   16252: result <= 12'b111110011000;
   16253: result <= 12'b111110011001;
   16254: result <= 12'b111110011010;
   16255: result <= 12'b111110011011;
   16256: result <= 12'b111110011100;
   16257: result <= 12'b111110011100;
   16258: result <= 12'b111110011101;
   16259: result <= 12'b111110011110;
   16260: result <= 12'b111110011111;
   16261: result <= 12'b111110011111;
   16262: result <= 12'b111110100000;
   16263: result <= 12'b111110100001;
   16264: result <= 12'b111110100010;
   16265: result <= 12'b111110100011;
   16266: result <= 12'b111110100011;
   16267: result <= 12'b111110100100;
   16268: result <= 12'b111110100101;
   16269: result <= 12'b111110100110;
   16270: result <= 12'b111110100110;
   16271: result <= 12'b111110100111;
   16272: result <= 12'b111110101000;
   16273: result <= 12'b111110101001;
   16274: result <= 12'b111110101010;
   16275: result <= 12'b111110101010;
   16276: result <= 12'b111110101011;
   16277: result <= 12'b111110101100;
   16278: result <= 12'b111110101101;
   16279: result <= 12'b111110101110;
   16280: result <= 12'b111110101110;
   16281: result <= 12'b111110101111;
   16282: result <= 12'b111110110000;
   16283: result <= 12'b111110110001;
   16284: result <= 12'b111110110001;
   16285: result <= 12'b111110110010;
   16286: result <= 12'b111110110011;
   16287: result <= 12'b111110110100;
   16288: result <= 12'b111110110101;
   16289: result <= 12'b111110110101;
   16290: result <= 12'b111110110110;
   16291: result <= 12'b111110110111;
   16292: result <= 12'b111110111000;
   16293: result <= 12'b111110111001;
   16294: result <= 12'b111110111001;
   16295: result <= 12'b111110111010;
   16296: result <= 12'b111110111011;
   16297: result <= 12'b111110111100;
   16298: result <= 12'b111110111100;
   16299: result <= 12'b111110111101;
   16300: result <= 12'b111110111110;
   16301: result <= 12'b111110111111;
   16302: result <= 12'b111111000000;
   16303: result <= 12'b111111000000;
   16304: result <= 12'b111111000001;
   16305: result <= 12'b111111000010;
   16306: result <= 12'b111111000011;
   16307: result <= 12'b111111000100;
   16308: result <= 12'b111111000100;
   16309: result <= 12'b111111000101;
   16310: result <= 12'b111111000110;
   16311: result <= 12'b111111000111;
   16312: result <= 12'b111111000111;
   16313: result <= 12'b111111001000;
   16314: result <= 12'b111111001001;
   16315: result <= 12'b111111001010;
   16316: result <= 12'b111111001011;
   16317: result <= 12'b111111001011;
   16318: result <= 12'b111111001100;
   16319: result <= 12'b111111001101;
   16320: result <= 12'b111111001110;
   16321: result <= 12'b111111001111;
   16322: result <= 12'b111111001111;
   16323: result <= 12'b111111010000;
   16324: result <= 12'b111111010001;
   16325: result <= 12'b111111010010;
   16326: result <= 12'b111111010010;
   16327: result <= 12'b111111010011;
   16328: result <= 12'b111111010100;
   16329: result <= 12'b111111010101;
   16330: result <= 12'b111111010110;
   16331: result <= 12'b111111010110;
   16332: result <= 12'b111111010111;
   16333: result <= 12'b111111011000;
   16334: result <= 12'b111111011001;
   16335: result <= 12'b111111011010;
   16336: result <= 12'b111111011010;
   16337: result <= 12'b111111011011;
   16338: result <= 12'b111111011100;
   16339: result <= 12'b111111011101;
   16340: result <= 12'b111111011101;
   16341: result <= 12'b111111011110;
   16342: result <= 12'b111111011111;
   16343: result <= 12'b111111100000;
   16344: result <= 12'b111111100001;
   16345: result <= 12'b111111100001;
   16346: result <= 12'b111111100010;
   16347: result <= 12'b111111100011;
   16348: result <= 12'b111111100100;
   16349: result <= 12'b111111100101;
   16350: result <= 12'b111111100101;
   16351: result <= 12'b111111100110;
   16352: result <= 12'b111111100111;
   16353: result <= 12'b111111101000;
   16354: result <= 12'b111111101000;
   16355: result <= 12'b111111101001;
   16356: result <= 12'b111111101010;
   16357: result <= 12'b111111101011;
   16358: result <= 12'b111111101100;
   16359: result <= 12'b111111101100;
   16360: result <= 12'b111111101101;
   16361: result <= 12'b111111101110;
   16362: result <= 12'b111111101111;
   16363: result <= 12'b111111110000;
   16364: result <= 12'b111111110000;
   16365: result <= 12'b111111110001;
   16366: result <= 12'b111111110010;
   16367: result <= 12'b111111110011;
   16368: result <= 12'b111111110011;
   16369: result <= 12'b111111110100;
   16370: result <= 12'b111111110101;
   16371: result <= 12'b111111110110;
   16372: result <= 12'b111111110111;
   16373: result <= 12'b111111110111;
   16374: result <= 12'b111111111000;
   16375: result <= 12'b111111111001;
   16376: result <= 12'b111111111010;
   16377: result <= 12'b111111111011;
   16378: result <= 12'b111111111011;
   16379: result <= 12'b111111111100;
   16380: result <= 12'b111111111101;
   16381: result <= 12'b111111111110;
   16382: result <= 12'b111111111110;
   16383: result <= 12'b111111111111;
   endcase
endmodule
