`timescale 1ns / 1ps
`default_nettype none


//Created by script createsinelookup.py
module sinetable(input wire [11:0] phase, input wire clk, output reg [7:0] result);

always @(posedge clk)
  case(phase)
   0: result <= 8'b00000000;
   1: result <= 8'b00000000;
   2: result <= 8'b00000000;
   3: result <= 8'b00000001;
   4: result <= 8'b00000001;
   5: result <= 8'b00000001;
   6: result <= 8'b00000001;
   7: result <= 8'b00000001;
   8: result <= 8'b00000010;
   9: result <= 8'b00000010;
   10: result <= 8'b00000010;
   11: result <= 8'b00000010;
   12: result <= 8'b00000010;
   13: result <= 8'b00000011;
   14: result <= 8'b00000011;
   15: result <= 8'b00000011;
   16: result <= 8'b00000011;
   17: result <= 8'b00000011;
   18: result <= 8'b00000100;
   19: result <= 8'b00000100;
   20: result <= 8'b00000100;
   21: result <= 8'b00000100;
   22: result <= 8'b00000100;
   23: result <= 8'b00000101;
   24: result <= 8'b00000101;
   25: result <= 8'b00000101;
   26: result <= 8'b00000101;
   27: result <= 8'b00000101;
   28: result <= 8'b00000101;
   29: result <= 8'b00000110;
   30: result <= 8'b00000110;
   31: result <= 8'b00000110;
   32: result <= 8'b00000110;
   33: result <= 8'b00000110;
   34: result <= 8'b00000111;
   35: result <= 8'b00000111;
   36: result <= 8'b00000111;
   37: result <= 8'b00000111;
   38: result <= 8'b00000111;
   39: result <= 8'b00001000;
   40: result <= 8'b00001000;
   41: result <= 8'b00001000;
   42: result <= 8'b00001000;
   43: result <= 8'b00001000;
   44: result <= 8'b00001001;
   45: result <= 8'b00001001;
   46: result <= 8'b00001001;
   47: result <= 8'b00001001;
   48: result <= 8'b00001001;
   49: result <= 8'b00001010;
   50: result <= 8'b00001010;
   51: result <= 8'b00001010;
   52: result <= 8'b00001010;
   53: result <= 8'b00001010;
   54: result <= 8'b00001011;
   55: result <= 8'b00001011;
   56: result <= 8'b00001011;
   57: result <= 8'b00001011;
   58: result <= 8'b00001011;
   59: result <= 8'b00001100;
   60: result <= 8'b00001100;
   61: result <= 8'b00001100;
   62: result <= 8'b00001100;
   63: result <= 8'b00001100;
   64: result <= 8'b00001101;
   65: result <= 8'b00001101;
   66: result <= 8'b00001101;
   67: result <= 8'b00001101;
   68: result <= 8'b00001101;
   69: result <= 8'b00001110;
   70: result <= 8'b00001110;
   71: result <= 8'b00001110;
   72: result <= 8'b00001110;
   73: result <= 8'b00001110;
   74: result <= 8'b00001110;
   75: result <= 8'b00001111;
   76: result <= 8'b00001111;
   77: result <= 8'b00001111;
   78: result <= 8'b00001111;
   79: result <= 8'b00001111;
   80: result <= 8'b00010000;
   81: result <= 8'b00010000;
   82: result <= 8'b00010000;
   83: result <= 8'b00010000;
   84: result <= 8'b00010000;
   85: result <= 8'b00010001;
   86: result <= 8'b00010001;
   87: result <= 8'b00010001;
   88: result <= 8'b00010001;
   89: result <= 8'b00010001;
   90: result <= 8'b00010010;
   91: result <= 8'b00010010;
   92: result <= 8'b00010010;
   93: result <= 8'b00010010;
   94: result <= 8'b00010010;
   95: result <= 8'b00010011;
   96: result <= 8'b00010011;
   97: result <= 8'b00010011;
   98: result <= 8'b00010011;
   99: result <= 8'b00010011;
   100: result <= 8'b00010100;
   101: result <= 8'b00010100;
   102: result <= 8'b00010100;
   103: result <= 8'b00010100;
   104: result <= 8'b00010100;
   105: result <= 8'b00010101;
   106: result <= 8'b00010101;
   107: result <= 8'b00010101;
   108: result <= 8'b00010101;
   109: result <= 8'b00010101;
   110: result <= 8'b00010101;
   111: result <= 8'b00010110;
   112: result <= 8'b00010110;
   113: result <= 8'b00010110;
   114: result <= 8'b00010110;
   115: result <= 8'b00010110;
   116: result <= 8'b00010111;
   117: result <= 8'b00010111;
   118: result <= 8'b00010111;
   119: result <= 8'b00010111;
   120: result <= 8'b00010111;
   121: result <= 8'b00011000;
   122: result <= 8'b00011000;
   123: result <= 8'b00011000;
   124: result <= 8'b00011000;
   125: result <= 8'b00011000;
   126: result <= 8'b00011001;
   127: result <= 8'b00011001;
   128: result <= 8'b00011001;
   129: result <= 8'b00011001;
   130: result <= 8'b00011001;
   131: result <= 8'b00011010;
   132: result <= 8'b00011010;
   133: result <= 8'b00011010;
   134: result <= 8'b00011010;
   135: result <= 8'b00011010;
   136: result <= 8'b00011011;
   137: result <= 8'b00011011;
   138: result <= 8'b00011011;
   139: result <= 8'b00011011;
   140: result <= 8'b00011011;
   141: result <= 8'b00011011;
   142: result <= 8'b00011100;
   143: result <= 8'b00011100;
   144: result <= 8'b00011100;
   145: result <= 8'b00011100;
   146: result <= 8'b00011100;
   147: result <= 8'b00011101;
   148: result <= 8'b00011101;
   149: result <= 8'b00011101;
   150: result <= 8'b00011101;
   151: result <= 8'b00011101;
   152: result <= 8'b00011110;
   153: result <= 8'b00011110;
   154: result <= 8'b00011110;
   155: result <= 8'b00011110;
   156: result <= 8'b00011110;
   157: result <= 8'b00011111;
   158: result <= 8'b00011111;
   159: result <= 8'b00011111;
   160: result <= 8'b00011111;
   161: result <= 8'b00011111;
   162: result <= 8'b00011111;
   163: result <= 8'b00100000;
   164: result <= 8'b00100000;
   165: result <= 8'b00100000;
   166: result <= 8'b00100000;
   167: result <= 8'b00100000;
   168: result <= 8'b00100001;
   169: result <= 8'b00100001;
   170: result <= 8'b00100001;
   171: result <= 8'b00100001;
   172: result <= 8'b00100001;
   173: result <= 8'b00100010;
   174: result <= 8'b00100010;
   175: result <= 8'b00100010;
   176: result <= 8'b00100010;
   177: result <= 8'b00100010;
   178: result <= 8'b00100011;
   179: result <= 8'b00100011;
   180: result <= 8'b00100011;
   181: result <= 8'b00100011;
   182: result <= 8'b00100011;
   183: result <= 8'b00100011;
   184: result <= 8'b00100100;
   185: result <= 8'b00100100;
   186: result <= 8'b00100100;
   187: result <= 8'b00100100;
   188: result <= 8'b00100100;
   189: result <= 8'b00100101;
   190: result <= 8'b00100101;
   191: result <= 8'b00100101;
   192: result <= 8'b00100101;
   193: result <= 8'b00100101;
   194: result <= 8'b00100110;
   195: result <= 8'b00100110;
   196: result <= 8'b00100110;
   197: result <= 8'b00100110;
   198: result <= 8'b00100110;
   199: result <= 8'b00100110;
   200: result <= 8'b00100111;
   201: result <= 8'b00100111;
   202: result <= 8'b00100111;
   203: result <= 8'b00100111;
   204: result <= 8'b00100111;
   205: result <= 8'b00101000;
   206: result <= 8'b00101000;
   207: result <= 8'b00101000;
   208: result <= 8'b00101000;
   209: result <= 8'b00101000;
   210: result <= 8'b00101001;
   211: result <= 8'b00101001;
   212: result <= 8'b00101001;
   213: result <= 8'b00101001;
   214: result <= 8'b00101001;
   215: result <= 8'b00101001;
   216: result <= 8'b00101010;
   217: result <= 8'b00101010;
   218: result <= 8'b00101010;
   219: result <= 8'b00101010;
   220: result <= 8'b00101010;
   221: result <= 8'b00101011;
   222: result <= 8'b00101011;
   223: result <= 8'b00101011;
   224: result <= 8'b00101011;
   225: result <= 8'b00101011;
   226: result <= 8'b00101011;
   227: result <= 8'b00101100;
   228: result <= 8'b00101100;
   229: result <= 8'b00101100;
   230: result <= 8'b00101100;
   231: result <= 8'b00101100;
   232: result <= 8'b00101101;
   233: result <= 8'b00101101;
   234: result <= 8'b00101101;
   235: result <= 8'b00101101;
   236: result <= 8'b00101101;
   237: result <= 8'b00101110;
   238: result <= 8'b00101110;
   239: result <= 8'b00101110;
   240: result <= 8'b00101110;
   241: result <= 8'b00101110;
   242: result <= 8'b00101110;
   243: result <= 8'b00101111;
   244: result <= 8'b00101111;
   245: result <= 8'b00101111;
   246: result <= 8'b00101111;
   247: result <= 8'b00101111;
   248: result <= 8'b00110000;
   249: result <= 8'b00110000;
   250: result <= 8'b00110000;
   251: result <= 8'b00110000;
   252: result <= 8'b00110000;
   253: result <= 8'b00110000;
   254: result <= 8'b00110001;
   255: result <= 8'b00110001;
   256: result <= 8'b00110001;
   257: result <= 8'b00110001;
   258: result <= 8'b00110001;
   259: result <= 8'b00110010;
   260: result <= 8'b00110010;
   261: result <= 8'b00110010;
   262: result <= 8'b00110010;
   263: result <= 8'b00110010;
   264: result <= 8'b00110010;
   265: result <= 8'b00110011;
   266: result <= 8'b00110011;
   267: result <= 8'b00110011;
   268: result <= 8'b00110011;
   269: result <= 8'b00110011;
   270: result <= 8'b00110100;
   271: result <= 8'b00110100;
   272: result <= 8'b00110100;
   273: result <= 8'b00110100;
   274: result <= 8'b00110100;
   275: result <= 8'b00110100;
   276: result <= 8'b00110101;
   277: result <= 8'b00110101;
   278: result <= 8'b00110101;
   279: result <= 8'b00110101;
   280: result <= 8'b00110101;
   281: result <= 8'b00110101;
   282: result <= 8'b00110110;
   283: result <= 8'b00110110;
   284: result <= 8'b00110110;
   285: result <= 8'b00110110;
   286: result <= 8'b00110110;
   287: result <= 8'b00110111;
   288: result <= 8'b00110111;
   289: result <= 8'b00110111;
   290: result <= 8'b00110111;
   291: result <= 8'b00110111;
   292: result <= 8'b00110111;
   293: result <= 8'b00111000;
   294: result <= 8'b00111000;
   295: result <= 8'b00111000;
   296: result <= 8'b00111000;
   297: result <= 8'b00111000;
   298: result <= 8'b00111000;
   299: result <= 8'b00111001;
   300: result <= 8'b00111001;
   301: result <= 8'b00111001;
   302: result <= 8'b00111001;
   303: result <= 8'b00111001;
   304: result <= 8'b00111010;
   305: result <= 8'b00111010;
   306: result <= 8'b00111010;
   307: result <= 8'b00111010;
   308: result <= 8'b00111010;
   309: result <= 8'b00111010;
   310: result <= 8'b00111011;
   311: result <= 8'b00111011;
   312: result <= 8'b00111011;
   313: result <= 8'b00111011;
   314: result <= 8'b00111011;
   315: result <= 8'b00111011;
   316: result <= 8'b00111100;
   317: result <= 8'b00111100;
   318: result <= 8'b00111100;
   319: result <= 8'b00111100;
   320: result <= 8'b00111100;
   321: result <= 8'b00111101;
   322: result <= 8'b00111101;
   323: result <= 8'b00111101;
   324: result <= 8'b00111101;
   325: result <= 8'b00111101;
   326: result <= 8'b00111101;
   327: result <= 8'b00111110;
   328: result <= 8'b00111110;
   329: result <= 8'b00111110;
   330: result <= 8'b00111110;
   331: result <= 8'b00111110;
   332: result <= 8'b00111110;
   333: result <= 8'b00111111;
   334: result <= 8'b00111111;
   335: result <= 8'b00111111;
   336: result <= 8'b00111111;
   337: result <= 8'b00111111;
   338: result <= 8'b00111111;
   339: result <= 8'b01000000;
   340: result <= 8'b01000000;
   341: result <= 8'b01000000;
   342: result <= 8'b01000000;
   343: result <= 8'b01000000;
   344: result <= 8'b01000000;
   345: result <= 8'b01000001;
   346: result <= 8'b01000001;
   347: result <= 8'b01000001;
   348: result <= 8'b01000001;
   349: result <= 8'b01000001;
   350: result <= 8'b01000001;
   351: result <= 8'b01000010;
   352: result <= 8'b01000010;
   353: result <= 8'b01000010;
   354: result <= 8'b01000010;
   355: result <= 8'b01000010;
   356: result <= 8'b01000010;
   357: result <= 8'b01000011;
   358: result <= 8'b01000011;
   359: result <= 8'b01000011;
   360: result <= 8'b01000011;
   361: result <= 8'b01000011;
   362: result <= 8'b01000011;
   363: result <= 8'b01000100;
   364: result <= 8'b01000100;
   365: result <= 8'b01000100;
   366: result <= 8'b01000100;
   367: result <= 8'b01000100;
   368: result <= 8'b01000100;
   369: result <= 8'b01000101;
   370: result <= 8'b01000101;
   371: result <= 8'b01000101;
   372: result <= 8'b01000101;
   373: result <= 8'b01000101;
   374: result <= 8'b01000101;
   375: result <= 8'b01000110;
   376: result <= 8'b01000110;
   377: result <= 8'b01000110;
   378: result <= 8'b01000110;
   379: result <= 8'b01000110;
   380: result <= 8'b01000110;
   381: result <= 8'b01000111;
   382: result <= 8'b01000111;
   383: result <= 8'b01000111;
   384: result <= 8'b01000111;
   385: result <= 8'b01000111;
   386: result <= 8'b01000111;
   387: result <= 8'b01001000;
   388: result <= 8'b01001000;
   389: result <= 8'b01001000;
   390: result <= 8'b01001000;
   391: result <= 8'b01001000;
   392: result <= 8'b01001000;
   393: result <= 8'b01001001;
   394: result <= 8'b01001001;
   395: result <= 8'b01001001;
   396: result <= 8'b01001001;
   397: result <= 8'b01001001;
   398: result <= 8'b01001001;
   399: result <= 8'b01001010;
   400: result <= 8'b01001010;
   401: result <= 8'b01001010;
   402: result <= 8'b01001010;
   403: result <= 8'b01001010;
   404: result <= 8'b01001010;
   405: result <= 8'b01001011;
   406: result <= 8'b01001011;
   407: result <= 8'b01001011;
   408: result <= 8'b01001011;
   409: result <= 8'b01001011;
   410: result <= 8'b01001011;
   411: result <= 8'b01001011;
   412: result <= 8'b01001100;
   413: result <= 8'b01001100;
   414: result <= 8'b01001100;
   415: result <= 8'b01001100;
   416: result <= 8'b01001100;
   417: result <= 8'b01001100;
   418: result <= 8'b01001101;
   419: result <= 8'b01001101;
   420: result <= 8'b01001101;
   421: result <= 8'b01001101;
   422: result <= 8'b01001101;
   423: result <= 8'b01001101;
   424: result <= 8'b01001110;
   425: result <= 8'b01001110;
   426: result <= 8'b01001110;
   427: result <= 8'b01001110;
   428: result <= 8'b01001110;
   429: result <= 8'b01001110;
   430: result <= 8'b01001110;
   431: result <= 8'b01001111;
   432: result <= 8'b01001111;
   433: result <= 8'b01001111;
   434: result <= 8'b01001111;
   435: result <= 8'b01001111;
   436: result <= 8'b01001111;
   437: result <= 8'b01010000;
   438: result <= 8'b01010000;
   439: result <= 8'b01010000;
   440: result <= 8'b01010000;
   441: result <= 8'b01010000;
   442: result <= 8'b01010000;
   443: result <= 8'b01010000;
   444: result <= 8'b01010001;
   445: result <= 8'b01010001;
   446: result <= 8'b01010001;
   447: result <= 8'b01010001;
   448: result <= 8'b01010001;
   449: result <= 8'b01010001;
   450: result <= 8'b01010010;
   451: result <= 8'b01010010;
   452: result <= 8'b01010010;
   453: result <= 8'b01010010;
   454: result <= 8'b01010010;
   455: result <= 8'b01010010;
   456: result <= 8'b01010010;
   457: result <= 8'b01010011;
   458: result <= 8'b01010011;
   459: result <= 8'b01010011;
   460: result <= 8'b01010011;
   461: result <= 8'b01010011;
   462: result <= 8'b01010011;
   463: result <= 8'b01010011;
   464: result <= 8'b01010100;
   465: result <= 8'b01010100;
   466: result <= 8'b01010100;
   467: result <= 8'b01010100;
   468: result <= 8'b01010100;
   469: result <= 8'b01010100;
   470: result <= 8'b01010100;
   471: result <= 8'b01010101;
   472: result <= 8'b01010101;
   473: result <= 8'b01010101;
   474: result <= 8'b01010101;
   475: result <= 8'b01010101;
   476: result <= 8'b01010101;
   477: result <= 8'b01010110;
   478: result <= 8'b01010110;
   479: result <= 8'b01010110;
   480: result <= 8'b01010110;
   481: result <= 8'b01010110;
   482: result <= 8'b01010110;
   483: result <= 8'b01010110;
   484: result <= 8'b01010111;
   485: result <= 8'b01010111;
   486: result <= 8'b01010111;
   487: result <= 8'b01010111;
   488: result <= 8'b01010111;
   489: result <= 8'b01010111;
   490: result <= 8'b01010111;
   491: result <= 8'b01011000;
   492: result <= 8'b01011000;
   493: result <= 8'b01011000;
   494: result <= 8'b01011000;
   495: result <= 8'b01011000;
   496: result <= 8'b01011000;
   497: result <= 8'b01011000;
   498: result <= 8'b01011001;
   499: result <= 8'b01011001;
   500: result <= 8'b01011001;
   501: result <= 8'b01011001;
   502: result <= 8'b01011001;
   503: result <= 8'b01011001;
   504: result <= 8'b01011001;
   505: result <= 8'b01011010;
   506: result <= 8'b01011010;
   507: result <= 8'b01011010;
   508: result <= 8'b01011010;
   509: result <= 8'b01011010;
   510: result <= 8'b01011010;
   511: result <= 8'b01011010;
   512: result <= 8'b01011011;
   513: result <= 8'b01011011;
   514: result <= 8'b01011011;
   515: result <= 8'b01011011;
   516: result <= 8'b01011011;
   517: result <= 8'b01011011;
   518: result <= 8'b01011011;
   519: result <= 8'b01011011;
   520: result <= 8'b01011100;
   521: result <= 8'b01011100;
   522: result <= 8'b01011100;
   523: result <= 8'b01011100;
   524: result <= 8'b01011100;
   525: result <= 8'b01011100;
   526: result <= 8'b01011100;
   527: result <= 8'b01011101;
   528: result <= 8'b01011101;
   529: result <= 8'b01011101;
   530: result <= 8'b01011101;
   531: result <= 8'b01011101;
   532: result <= 8'b01011101;
   533: result <= 8'b01011101;
   534: result <= 8'b01011110;
   535: result <= 8'b01011110;
   536: result <= 8'b01011110;
   537: result <= 8'b01011110;
   538: result <= 8'b01011110;
   539: result <= 8'b01011110;
   540: result <= 8'b01011110;
   541: result <= 8'b01011110;
   542: result <= 8'b01011111;
   543: result <= 8'b01011111;
   544: result <= 8'b01011111;
   545: result <= 8'b01011111;
   546: result <= 8'b01011111;
   547: result <= 8'b01011111;
   548: result <= 8'b01011111;
   549: result <= 8'b01011111;
   550: result <= 8'b01100000;
   551: result <= 8'b01100000;
   552: result <= 8'b01100000;
   553: result <= 8'b01100000;
   554: result <= 8'b01100000;
   555: result <= 8'b01100000;
   556: result <= 8'b01100000;
   557: result <= 8'b01100001;
   558: result <= 8'b01100001;
   559: result <= 8'b01100001;
   560: result <= 8'b01100001;
   561: result <= 8'b01100001;
   562: result <= 8'b01100001;
   563: result <= 8'b01100001;
   564: result <= 8'b01100001;
   565: result <= 8'b01100010;
   566: result <= 8'b01100010;
   567: result <= 8'b01100010;
   568: result <= 8'b01100010;
   569: result <= 8'b01100010;
   570: result <= 8'b01100010;
   571: result <= 8'b01100010;
   572: result <= 8'b01100010;
   573: result <= 8'b01100011;
   574: result <= 8'b01100011;
   575: result <= 8'b01100011;
   576: result <= 8'b01100011;
   577: result <= 8'b01100011;
   578: result <= 8'b01100011;
   579: result <= 8'b01100011;
   580: result <= 8'b01100011;
   581: result <= 8'b01100100;
   582: result <= 8'b01100100;
   583: result <= 8'b01100100;
   584: result <= 8'b01100100;
   585: result <= 8'b01100100;
   586: result <= 8'b01100100;
   587: result <= 8'b01100100;
   588: result <= 8'b01100100;
   589: result <= 8'b01100101;
   590: result <= 8'b01100101;
   591: result <= 8'b01100101;
   592: result <= 8'b01100101;
   593: result <= 8'b01100101;
   594: result <= 8'b01100101;
   595: result <= 8'b01100101;
   596: result <= 8'b01100101;
   597: result <= 8'b01100110;
   598: result <= 8'b01100110;
   599: result <= 8'b01100110;
   600: result <= 8'b01100110;
   601: result <= 8'b01100110;
   602: result <= 8'b01100110;
   603: result <= 8'b01100110;
   604: result <= 8'b01100110;
   605: result <= 8'b01100110;
   606: result <= 8'b01100111;
   607: result <= 8'b01100111;
   608: result <= 8'b01100111;
   609: result <= 8'b01100111;
   610: result <= 8'b01100111;
   611: result <= 8'b01100111;
   612: result <= 8'b01100111;
   613: result <= 8'b01100111;
   614: result <= 8'b01101000;
   615: result <= 8'b01101000;
   616: result <= 8'b01101000;
   617: result <= 8'b01101000;
   618: result <= 8'b01101000;
   619: result <= 8'b01101000;
   620: result <= 8'b01101000;
   621: result <= 8'b01101000;
   622: result <= 8'b01101000;
   623: result <= 8'b01101001;
   624: result <= 8'b01101001;
   625: result <= 8'b01101001;
   626: result <= 8'b01101001;
   627: result <= 8'b01101001;
   628: result <= 8'b01101001;
   629: result <= 8'b01101001;
   630: result <= 8'b01101001;
   631: result <= 8'b01101001;
   632: result <= 8'b01101010;
   633: result <= 8'b01101010;
   634: result <= 8'b01101010;
   635: result <= 8'b01101010;
   636: result <= 8'b01101010;
   637: result <= 8'b01101010;
   638: result <= 8'b01101010;
   639: result <= 8'b01101010;
   640: result <= 8'b01101010;
   641: result <= 8'b01101011;
   642: result <= 8'b01101011;
   643: result <= 8'b01101011;
   644: result <= 8'b01101011;
   645: result <= 8'b01101011;
   646: result <= 8'b01101011;
   647: result <= 8'b01101011;
   648: result <= 8'b01101011;
   649: result <= 8'b01101011;
   650: result <= 8'b01101100;
   651: result <= 8'b01101100;
   652: result <= 8'b01101100;
   653: result <= 8'b01101100;
   654: result <= 8'b01101100;
   655: result <= 8'b01101100;
   656: result <= 8'b01101100;
   657: result <= 8'b01101100;
   658: result <= 8'b01101100;
   659: result <= 8'b01101100;
   660: result <= 8'b01101101;
   661: result <= 8'b01101101;
   662: result <= 8'b01101101;
   663: result <= 8'b01101101;
   664: result <= 8'b01101101;
   665: result <= 8'b01101101;
   666: result <= 8'b01101101;
   667: result <= 8'b01101101;
   668: result <= 8'b01101101;
   669: result <= 8'b01101101;
   670: result <= 8'b01101110;
   671: result <= 8'b01101110;
   672: result <= 8'b01101110;
   673: result <= 8'b01101110;
   674: result <= 8'b01101110;
   675: result <= 8'b01101110;
   676: result <= 8'b01101110;
   677: result <= 8'b01101110;
   678: result <= 8'b01101110;
   679: result <= 8'b01101110;
   680: result <= 8'b01101111;
   681: result <= 8'b01101111;
   682: result <= 8'b01101111;
   683: result <= 8'b01101111;
   684: result <= 8'b01101111;
   685: result <= 8'b01101111;
   686: result <= 8'b01101111;
   687: result <= 8'b01101111;
   688: result <= 8'b01101111;
   689: result <= 8'b01101111;
   690: result <= 8'b01110000;
   691: result <= 8'b01110000;
   692: result <= 8'b01110000;
   693: result <= 8'b01110000;
   694: result <= 8'b01110000;
   695: result <= 8'b01110000;
   696: result <= 8'b01110000;
   697: result <= 8'b01110000;
   698: result <= 8'b01110000;
   699: result <= 8'b01110000;
   700: result <= 8'b01110001;
   701: result <= 8'b01110001;
   702: result <= 8'b01110001;
   703: result <= 8'b01110001;
   704: result <= 8'b01110001;
   705: result <= 8'b01110001;
   706: result <= 8'b01110001;
   707: result <= 8'b01110001;
   708: result <= 8'b01110001;
   709: result <= 8'b01110001;
   710: result <= 8'b01110001;
   711: result <= 8'b01110010;
   712: result <= 8'b01110010;
   713: result <= 8'b01110010;
   714: result <= 8'b01110010;
   715: result <= 8'b01110010;
   716: result <= 8'b01110010;
   717: result <= 8'b01110010;
   718: result <= 8'b01110010;
   719: result <= 8'b01110010;
   720: result <= 8'b01110010;
   721: result <= 8'b01110010;
   722: result <= 8'b01110011;
   723: result <= 8'b01110011;
   724: result <= 8'b01110011;
   725: result <= 8'b01110011;
   726: result <= 8'b01110011;
   727: result <= 8'b01110011;
   728: result <= 8'b01110011;
   729: result <= 8'b01110011;
   730: result <= 8'b01110011;
   731: result <= 8'b01110011;
   732: result <= 8'b01110011;
   733: result <= 8'b01110011;
   734: result <= 8'b01110100;
   735: result <= 8'b01110100;
   736: result <= 8'b01110100;
   737: result <= 8'b01110100;
   738: result <= 8'b01110100;
   739: result <= 8'b01110100;
   740: result <= 8'b01110100;
   741: result <= 8'b01110100;
   742: result <= 8'b01110100;
   743: result <= 8'b01110100;
   744: result <= 8'b01110100;
   745: result <= 8'b01110100;
   746: result <= 8'b01110101;
   747: result <= 8'b01110101;
   748: result <= 8'b01110101;
   749: result <= 8'b01110101;
   750: result <= 8'b01110101;
   751: result <= 8'b01110101;
   752: result <= 8'b01110101;
   753: result <= 8'b01110101;
   754: result <= 8'b01110101;
   755: result <= 8'b01110101;
   756: result <= 8'b01110101;
   757: result <= 8'b01110101;
   758: result <= 8'b01110101;
   759: result <= 8'b01110110;
   760: result <= 8'b01110110;
   761: result <= 8'b01110110;
   762: result <= 8'b01110110;
   763: result <= 8'b01110110;
   764: result <= 8'b01110110;
   765: result <= 8'b01110110;
   766: result <= 8'b01110110;
   767: result <= 8'b01110110;
   768: result <= 8'b01110110;
   769: result <= 8'b01110110;
   770: result <= 8'b01110110;
   771: result <= 8'b01110110;
   772: result <= 8'b01110111;
   773: result <= 8'b01110111;
   774: result <= 8'b01110111;
   775: result <= 8'b01110111;
   776: result <= 8'b01110111;
   777: result <= 8'b01110111;
   778: result <= 8'b01110111;
   779: result <= 8'b01110111;
   780: result <= 8'b01110111;
   781: result <= 8'b01110111;
   782: result <= 8'b01110111;
   783: result <= 8'b01110111;
   784: result <= 8'b01110111;
   785: result <= 8'b01110111;
   786: result <= 8'b01111000;
   787: result <= 8'b01111000;
   788: result <= 8'b01111000;
   789: result <= 8'b01111000;
   790: result <= 8'b01111000;
   791: result <= 8'b01111000;
   792: result <= 8'b01111000;
   793: result <= 8'b01111000;
   794: result <= 8'b01111000;
   795: result <= 8'b01111000;
   796: result <= 8'b01111000;
   797: result <= 8'b01111000;
   798: result <= 8'b01111000;
   799: result <= 8'b01111000;
   800: result <= 8'b01111001;
   801: result <= 8'b01111001;
   802: result <= 8'b01111001;
   803: result <= 8'b01111001;
   804: result <= 8'b01111001;
   805: result <= 8'b01111001;
   806: result <= 8'b01111001;
   807: result <= 8'b01111001;
   808: result <= 8'b01111001;
   809: result <= 8'b01111001;
   810: result <= 8'b01111001;
   811: result <= 8'b01111001;
   812: result <= 8'b01111001;
   813: result <= 8'b01111001;
   814: result <= 8'b01111001;
   815: result <= 8'b01111001;
   816: result <= 8'b01111010;
   817: result <= 8'b01111010;
   818: result <= 8'b01111010;
   819: result <= 8'b01111010;
   820: result <= 8'b01111010;
   821: result <= 8'b01111010;
   822: result <= 8'b01111010;
   823: result <= 8'b01111010;
   824: result <= 8'b01111010;
   825: result <= 8'b01111010;
   826: result <= 8'b01111010;
   827: result <= 8'b01111010;
   828: result <= 8'b01111010;
   829: result <= 8'b01111010;
   830: result <= 8'b01111010;
   831: result <= 8'b01111010;
   832: result <= 8'b01111010;
   833: result <= 8'b01111011;
   834: result <= 8'b01111011;
   835: result <= 8'b01111011;
   836: result <= 8'b01111011;
   837: result <= 8'b01111011;
   838: result <= 8'b01111011;
   839: result <= 8'b01111011;
   840: result <= 8'b01111011;
   841: result <= 8'b01111011;
   842: result <= 8'b01111011;
   843: result <= 8'b01111011;
   844: result <= 8'b01111011;
   845: result <= 8'b01111011;
   846: result <= 8'b01111011;
   847: result <= 8'b01111011;
   848: result <= 8'b01111011;
   849: result <= 8'b01111011;
   850: result <= 8'b01111011;
   851: result <= 8'b01111100;
   852: result <= 8'b01111100;
   853: result <= 8'b01111100;
   854: result <= 8'b01111100;
   855: result <= 8'b01111100;
   856: result <= 8'b01111100;
   857: result <= 8'b01111100;
   858: result <= 8'b01111100;
   859: result <= 8'b01111100;
   860: result <= 8'b01111100;
   861: result <= 8'b01111100;
   862: result <= 8'b01111100;
   863: result <= 8'b01111100;
   864: result <= 8'b01111100;
   865: result <= 8'b01111100;
   866: result <= 8'b01111100;
   867: result <= 8'b01111100;
   868: result <= 8'b01111100;
   869: result <= 8'b01111100;
   870: result <= 8'b01111100;
   871: result <= 8'b01111100;
   872: result <= 8'b01111101;
   873: result <= 8'b01111101;
   874: result <= 8'b01111101;
   875: result <= 8'b01111101;
   876: result <= 8'b01111101;
   877: result <= 8'b01111101;
   878: result <= 8'b01111101;
   879: result <= 8'b01111101;
   880: result <= 8'b01111101;
   881: result <= 8'b01111101;
   882: result <= 8'b01111101;
   883: result <= 8'b01111101;
   884: result <= 8'b01111101;
   885: result <= 8'b01111101;
   886: result <= 8'b01111101;
   887: result <= 8'b01111101;
   888: result <= 8'b01111101;
   889: result <= 8'b01111101;
   890: result <= 8'b01111101;
   891: result <= 8'b01111101;
   892: result <= 8'b01111101;
   893: result <= 8'b01111101;
   894: result <= 8'b01111101;
   895: result <= 8'b01111110;
   896: result <= 8'b01111110;
   897: result <= 8'b01111110;
   898: result <= 8'b01111110;
   899: result <= 8'b01111110;
   900: result <= 8'b01111110;
   901: result <= 8'b01111110;
   902: result <= 8'b01111110;
   903: result <= 8'b01111110;
   904: result <= 8'b01111110;
   905: result <= 8'b01111110;
   906: result <= 8'b01111110;
   907: result <= 8'b01111110;
   908: result <= 8'b01111110;
   909: result <= 8'b01111110;
   910: result <= 8'b01111110;
   911: result <= 8'b01111110;
   912: result <= 8'b01111110;
   913: result <= 8'b01111110;
   914: result <= 8'b01111110;
   915: result <= 8'b01111110;
   916: result <= 8'b01111110;
   917: result <= 8'b01111110;
   918: result <= 8'b01111110;
   919: result <= 8'b01111110;
   920: result <= 8'b01111110;
   921: result <= 8'b01111110;
   922: result <= 8'b01111110;
   923: result <= 8'b01111110;
   924: result <= 8'b01111110;
   925: result <= 8'b01111111;
   926: result <= 8'b01111111;
   927: result <= 8'b01111111;
   928: result <= 8'b01111111;
   929: result <= 8'b01111111;
   930: result <= 8'b01111111;
   931: result <= 8'b01111111;
   932: result <= 8'b01111111;
   933: result <= 8'b01111111;
   934: result <= 8'b01111111;
   935: result <= 8'b01111111;
   936: result <= 8'b01111111;
   937: result <= 8'b01111111;
   938: result <= 8'b01111111;
   939: result <= 8'b01111111;
   940: result <= 8'b01111111;
   941: result <= 8'b01111111;
   942: result <= 8'b01111111;
   943: result <= 8'b01111111;
   944: result <= 8'b01111111;
   945: result <= 8'b01111111;
   946: result <= 8'b01111111;
   947: result <= 8'b01111111;
   948: result <= 8'b01111111;
   949: result <= 8'b01111111;
   950: result <= 8'b01111111;
   951: result <= 8'b01111111;
   952: result <= 8'b01111111;
   953: result <= 8'b01111111;
   954: result <= 8'b01111111;
   955: result <= 8'b01111111;
   956: result <= 8'b01111111;
   957: result <= 8'b01111111;
   958: result <= 8'b01111111;
   959: result <= 8'b01111111;
   960: result <= 8'b01111111;
   961: result <= 8'b01111111;
   962: result <= 8'b01111111;
   963: result <= 8'b01111111;
   964: result <= 8'b01111111;
   965: result <= 8'b01111111;
   966: result <= 8'b01111111;
   967: result <= 8'b01111111;
   968: result <= 8'b01111111;
   969: result <= 8'b01111111;
   970: result <= 8'b01111111;
   971: result <= 8'b01111111;
   972: result <= 8'b01111111;
   973: result <= 8'b01111111;
   974: result <= 8'b01111111;
   975: result <= 8'b01111111;
   976: result <= 8'b01111111;
   977: result <= 8'b01111111;
   978: result <= 8'b01111111;
   979: result <= 8'b01111111;
   980: result <= 8'b01111111;
   981: result <= 8'b01111111;
   982: result <= 8'b01111111;
   983: result <= 8'b01111111;
   984: result <= 8'b01111111;
   985: result <= 8'b01111111;
   986: result <= 8'b01111111;
   987: result <= 8'b01111111;
   988: result <= 8'b01111111;
   989: result <= 8'b01111111;
   990: result <= 8'b01111111;
   991: result <= 8'b01111111;
   992: result <= 8'b01111111;
   993: result <= 8'b01111111;
   994: result <= 8'b01111111;
   995: result <= 8'b01111111;
   996: result <= 8'b01111111;
   997: result <= 8'b01111111;
   998: result <= 8'b01111111;
   999: result <= 8'b01111111;
   1000: result <= 8'b01111111;
   1001: result <= 8'b01111111;
   1002: result <= 8'b01111111;
   1003: result <= 8'b01111111;
   1004: result <= 8'b01111111;
   1005: result <= 8'b01111111;
   1006: result <= 8'b01111111;
   1007: result <= 8'b01111111;
   1008: result <= 8'b01111111;
   1009: result <= 8'b01111111;
   1010: result <= 8'b01111111;
   1011: result <= 8'b01111111;
   1012: result <= 8'b01111111;
   1013: result <= 8'b01111111;
   1014: result <= 8'b01111111;
   1015: result <= 8'b01111111;
   1016: result <= 8'b01111111;
   1017: result <= 8'b01111111;
   1018: result <= 8'b01111111;
   1019: result <= 8'b01111111;
   1020: result <= 8'b01111111;
   1021: result <= 8'b01111111;
   1022: result <= 8'b01111111;
   1023: result <= 8'b01111111;
   1024: result <= 8'b01111111;
   1025: result <= 8'b01111111;
   1026: result <= 8'b01111111;
   1027: result <= 8'b01111111;
   1028: result <= 8'b01111111;
   1029: result <= 8'b01111111;
   1030: result <= 8'b01111111;
   1031: result <= 8'b01111111;
   1032: result <= 8'b01111111;
   1033: result <= 8'b01111111;
   1034: result <= 8'b01111111;
   1035: result <= 8'b01111111;
   1036: result <= 8'b01111111;
   1037: result <= 8'b01111111;
   1038: result <= 8'b01111111;
   1039: result <= 8'b01111111;
   1040: result <= 8'b01111111;
   1041: result <= 8'b01111111;
   1042: result <= 8'b01111111;
   1043: result <= 8'b01111111;
   1044: result <= 8'b01111111;
   1045: result <= 8'b01111111;
   1046: result <= 8'b01111111;
   1047: result <= 8'b01111111;
   1048: result <= 8'b01111111;
   1049: result <= 8'b01111111;
   1050: result <= 8'b01111111;
   1051: result <= 8'b01111111;
   1052: result <= 8'b01111111;
   1053: result <= 8'b01111111;
   1054: result <= 8'b01111111;
   1055: result <= 8'b01111111;
   1056: result <= 8'b01111111;
   1057: result <= 8'b01111111;
   1058: result <= 8'b01111111;
   1059: result <= 8'b01111111;
   1060: result <= 8'b01111111;
   1061: result <= 8'b01111111;
   1062: result <= 8'b01111111;
   1063: result <= 8'b01111111;
   1064: result <= 8'b01111111;
   1065: result <= 8'b01111111;
   1066: result <= 8'b01111111;
   1067: result <= 8'b01111111;
   1068: result <= 8'b01111111;
   1069: result <= 8'b01111111;
   1070: result <= 8'b01111111;
   1071: result <= 8'b01111111;
   1072: result <= 8'b01111111;
   1073: result <= 8'b01111111;
   1074: result <= 8'b01111111;
   1075: result <= 8'b01111111;
   1076: result <= 8'b01111111;
   1077: result <= 8'b01111111;
   1078: result <= 8'b01111111;
   1079: result <= 8'b01111111;
   1080: result <= 8'b01111111;
   1081: result <= 8'b01111111;
   1082: result <= 8'b01111111;
   1083: result <= 8'b01111111;
   1084: result <= 8'b01111111;
   1085: result <= 8'b01111111;
   1086: result <= 8'b01111111;
   1087: result <= 8'b01111111;
   1088: result <= 8'b01111111;
   1089: result <= 8'b01111111;
   1090: result <= 8'b01111111;
   1091: result <= 8'b01111111;
   1092: result <= 8'b01111111;
   1093: result <= 8'b01111111;
   1094: result <= 8'b01111111;
   1095: result <= 8'b01111111;
   1096: result <= 8'b01111111;
   1097: result <= 8'b01111111;
   1098: result <= 8'b01111111;
   1099: result <= 8'b01111111;
   1100: result <= 8'b01111111;
   1101: result <= 8'b01111111;
   1102: result <= 8'b01111111;
   1103: result <= 8'b01111111;
   1104: result <= 8'b01111111;
   1105: result <= 8'b01111111;
   1106: result <= 8'b01111111;
   1107: result <= 8'b01111111;
   1108: result <= 8'b01111111;
   1109: result <= 8'b01111111;
   1110: result <= 8'b01111111;
   1111: result <= 8'b01111111;
   1112: result <= 8'b01111111;
   1113: result <= 8'b01111111;
   1114: result <= 8'b01111111;
   1115: result <= 8'b01111111;
   1116: result <= 8'b01111111;
   1117: result <= 8'b01111111;
   1118: result <= 8'b01111111;
   1119: result <= 8'b01111111;
   1120: result <= 8'b01111111;
   1121: result <= 8'b01111111;
   1122: result <= 8'b01111111;
   1123: result <= 8'b01111111;
   1124: result <= 8'b01111110;
   1125: result <= 8'b01111110;
   1126: result <= 8'b01111110;
   1127: result <= 8'b01111110;
   1128: result <= 8'b01111110;
   1129: result <= 8'b01111110;
   1130: result <= 8'b01111110;
   1131: result <= 8'b01111110;
   1132: result <= 8'b01111110;
   1133: result <= 8'b01111110;
   1134: result <= 8'b01111110;
   1135: result <= 8'b01111110;
   1136: result <= 8'b01111110;
   1137: result <= 8'b01111110;
   1138: result <= 8'b01111110;
   1139: result <= 8'b01111110;
   1140: result <= 8'b01111110;
   1141: result <= 8'b01111110;
   1142: result <= 8'b01111110;
   1143: result <= 8'b01111110;
   1144: result <= 8'b01111110;
   1145: result <= 8'b01111110;
   1146: result <= 8'b01111110;
   1147: result <= 8'b01111110;
   1148: result <= 8'b01111110;
   1149: result <= 8'b01111110;
   1150: result <= 8'b01111110;
   1151: result <= 8'b01111110;
   1152: result <= 8'b01111110;
   1153: result <= 8'b01111110;
   1154: result <= 8'b01111101;
   1155: result <= 8'b01111101;
   1156: result <= 8'b01111101;
   1157: result <= 8'b01111101;
   1158: result <= 8'b01111101;
   1159: result <= 8'b01111101;
   1160: result <= 8'b01111101;
   1161: result <= 8'b01111101;
   1162: result <= 8'b01111101;
   1163: result <= 8'b01111101;
   1164: result <= 8'b01111101;
   1165: result <= 8'b01111101;
   1166: result <= 8'b01111101;
   1167: result <= 8'b01111101;
   1168: result <= 8'b01111101;
   1169: result <= 8'b01111101;
   1170: result <= 8'b01111101;
   1171: result <= 8'b01111101;
   1172: result <= 8'b01111101;
   1173: result <= 8'b01111101;
   1174: result <= 8'b01111101;
   1175: result <= 8'b01111101;
   1176: result <= 8'b01111101;
   1177: result <= 8'b01111100;
   1178: result <= 8'b01111100;
   1179: result <= 8'b01111100;
   1180: result <= 8'b01111100;
   1181: result <= 8'b01111100;
   1182: result <= 8'b01111100;
   1183: result <= 8'b01111100;
   1184: result <= 8'b01111100;
   1185: result <= 8'b01111100;
   1186: result <= 8'b01111100;
   1187: result <= 8'b01111100;
   1188: result <= 8'b01111100;
   1189: result <= 8'b01111100;
   1190: result <= 8'b01111100;
   1191: result <= 8'b01111100;
   1192: result <= 8'b01111100;
   1193: result <= 8'b01111100;
   1194: result <= 8'b01111100;
   1195: result <= 8'b01111100;
   1196: result <= 8'b01111100;
   1197: result <= 8'b01111100;
   1198: result <= 8'b01111011;
   1199: result <= 8'b01111011;
   1200: result <= 8'b01111011;
   1201: result <= 8'b01111011;
   1202: result <= 8'b01111011;
   1203: result <= 8'b01111011;
   1204: result <= 8'b01111011;
   1205: result <= 8'b01111011;
   1206: result <= 8'b01111011;
   1207: result <= 8'b01111011;
   1208: result <= 8'b01111011;
   1209: result <= 8'b01111011;
   1210: result <= 8'b01111011;
   1211: result <= 8'b01111011;
   1212: result <= 8'b01111011;
   1213: result <= 8'b01111011;
   1214: result <= 8'b01111011;
   1215: result <= 8'b01111011;
   1216: result <= 8'b01111010;
   1217: result <= 8'b01111010;
   1218: result <= 8'b01111010;
   1219: result <= 8'b01111010;
   1220: result <= 8'b01111010;
   1221: result <= 8'b01111010;
   1222: result <= 8'b01111010;
   1223: result <= 8'b01111010;
   1224: result <= 8'b01111010;
   1225: result <= 8'b01111010;
   1226: result <= 8'b01111010;
   1227: result <= 8'b01111010;
   1228: result <= 8'b01111010;
   1229: result <= 8'b01111010;
   1230: result <= 8'b01111010;
   1231: result <= 8'b01111010;
   1232: result <= 8'b01111010;
   1233: result <= 8'b01111001;
   1234: result <= 8'b01111001;
   1235: result <= 8'b01111001;
   1236: result <= 8'b01111001;
   1237: result <= 8'b01111001;
   1238: result <= 8'b01111001;
   1239: result <= 8'b01111001;
   1240: result <= 8'b01111001;
   1241: result <= 8'b01111001;
   1242: result <= 8'b01111001;
   1243: result <= 8'b01111001;
   1244: result <= 8'b01111001;
   1245: result <= 8'b01111001;
   1246: result <= 8'b01111001;
   1247: result <= 8'b01111001;
   1248: result <= 8'b01111001;
   1249: result <= 8'b01111000;
   1250: result <= 8'b01111000;
   1251: result <= 8'b01111000;
   1252: result <= 8'b01111000;
   1253: result <= 8'b01111000;
   1254: result <= 8'b01111000;
   1255: result <= 8'b01111000;
   1256: result <= 8'b01111000;
   1257: result <= 8'b01111000;
   1258: result <= 8'b01111000;
   1259: result <= 8'b01111000;
   1260: result <= 8'b01111000;
   1261: result <= 8'b01111000;
   1262: result <= 8'b01111000;
   1263: result <= 8'b01110111;
   1264: result <= 8'b01110111;
   1265: result <= 8'b01110111;
   1266: result <= 8'b01110111;
   1267: result <= 8'b01110111;
   1268: result <= 8'b01110111;
   1269: result <= 8'b01110111;
   1270: result <= 8'b01110111;
   1271: result <= 8'b01110111;
   1272: result <= 8'b01110111;
   1273: result <= 8'b01110111;
   1274: result <= 8'b01110111;
   1275: result <= 8'b01110111;
   1276: result <= 8'b01110111;
   1277: result <= 8'b01110110;
   1278: result <= 8'b01110110;
   1279: result <= 8'b01110110;
   1280: result <= 8'b01110110;
   1281: result <= 8'b01110110;
   1282: result <= 8'b01110110;
   1283: result <= 8'b01110110;
   1284: result <= 8'b01110110;
   1285: result <= 8'b01110110;
   1286: result <= 8'b01110110;
   1287: result <= 8'b01110110;
   1288: result <= 8'b01110110;
   1289: result <= 8'b01110110;
   1290: result <= 8'b01110101;
   1291: result <= 8'b01110101;
   1292: result <= 8'b01110101;
   1293: result <= 8'b01110101;
   1294: result <= 8'b01110101;
   1295: result <= 8'b01110101;
   1296: result <= 8'b01110101;
   1297: result <= 8'b01110101;
   1298: result <= 8'b01110101;
   1299: result <= 8'b01110101;
   1300: result <= 8'b01110101;
   1301: result <= 8'b01110101;
   1302: result <= 8'b01110101;
   1303: result <= 8'b01110100;
   1304: result <= 8'b01110100;
   1305: result <= 8'b01110100;
   1306: result <= 8'b01110100;
   1307: result <= 8'b01110100;
   1308: result <= 8'b01110100;
   1309: result <= 8'b01110100;
   1310: result <= 8'b01110100;
   1311: result <= 8'b01110100;
   1312: result <= 8'b01110100;
   1313: result <= 8'b01110100;
   1314: result <= 8'b01110100;
   1315: result <= 8'b01110011;
   1316: result <= 8'b01110011;
   1317: result <= 8'b01110011;
   1318: result <= 8'b01110011;
   1319: result <= 8'b01110011;
   1320: result <= 8'b01110011;
   1321: result <= 8'b01110011;
   1322: result <= 8'b01110011;
   1323: result <= 8'b01110011;
   1324: result <= 8'b01110011;
   1325: result <= 8'b01110011;
   1326: result <= 8'b01110011;
   1327: result <= 8'b01110010;
   1328: result <= 8'b01110010;
   1329: result <= 8'b01110010;
   1330: result <= 8'b01110010;
   1331: result <= 8'b01110010;
   1332: result <= 8'b01110010;
   1333: result <= 8'b01110010;
   1334: result <= 8'b01110010;
   1335: result <= 8'b01110010;
   1336: result <= 8'b01110010;
   1337: result <= 8'b01110010;
   1338: result <= 8'b01110001;
   1339: result <= 8'b01110001;
   1340: result <= 8'b01110001;
   1341: result <= 8'b01110001;
   1342: result <= 8'b01110001;
   1343: result <= 8'b01110001;
   1344: result <= 8'b01110001;
   1345: result <= 8'b01110001;
   1346: result <= 8'b01110001;
   1347: result <= 8'b01110001;
   1348: result <= 8'b01110001;
   1349: result <= 8'b01110000;
   1350: result <= 8'b01110000;
   1351: result <= 8'b01110000;
   1352: result <= 8'b01110000;
   1353: result <= 8'b01110000;
   1354: result <= 8'b01110000;
   1355: result <= 8'b01110000;
   1356: result <= 8'b01110000;
   1357: result <= 8'b01110000;
   1358: result <= 8'b01110000;
   1359: result <= 8'b01101111;
   1360: result <= 8'b01101111;
   1361: result <= 8'b01101111;
   1362: result <= 8'b01101111;
   1363: result <= 8'b01101111;
   1364: result <= 8'b01101111;
   1365: result <= 8'b01101111;
   1366: result <= 8'b01101111;
   1367: result <= 8'b01101111;
   1368: result <= 8'b01101111;
   1369: result <= 8'b01101110;
   1370: result <= 8'b01101110;
   1371: result <= 8'b01101110;
   1372: result <= 8'b01101110;
   1373: result <= 8'b01101110;
   1374: result <= 8'b01101110;
   1375: result <= 8'b01101110;
   1376: result <= 8'b01101110;
   1377: result <= 8'b01101110;
   1378: result <= 8'b01101110;
   1379: result <= 8'b01101101;
   1380: result <= 8'b01101101;
   1381: result <= 8'b01101101;
   1382: result <= 8'b01101101;
   1383: result <= 8'b01101101;
   1384: result <= 8'b01101101;
   1385: result <= 8'b01101101;
   1386: result <= 8'b01101101;
   1387: result <= 8'b01101101;
   1388: result <= 8'b01101101;
   1389: result <= 8'b01101100;
   1390: result <= 8'b01101100;
   1391: result <= 8'b01101100;
   1392: result <= 8'b01101100;
   1393: result <= 8'b01101100;
   1394: result <= 8'b01101100;
   1395: result <= 8'b01101100;
   1396: result <= 8'b01101100;
   1397: result <= 8'b01101100;
   1398: result <= 8'b01101100;
   1399: result <= 8'b01101011;
   1400: result <= 8'b01101011;
   1401: result <= 8'b01101011;
   1402: result <= 8'b01101011;
   1403: result <= 8'b01101011;
   1404: result <= 8'b01101011;
   1405: result <= 8'b01101011;
   1406: result <= 8'b01101011;
   1407: result <= 8'b01101011;
   1408: result <= 8'b01101010;
   1409: result <= 8'b01101010;
   1410: result <= 8'b01101010;
   1411: result <= 8'b01101010;
   1412: result <= 8'b01101010;
   1413: result <= 8'b01101010;
   1414: result <= 8'b01101010;
   1415: result <= 8'b01101010;
   1416: result <= 8'b01101010;
   1417: result <= 8'b01101001;
   1418: result <= 8'b01101001;
   1419: result <= 8'b01101001;
   1420: result <= 8'b01101001;
   1421: result <= 8'b01101001;
   1422: result <= 8'b01101001;
   1423: result <= 8'b01101001;
   1424: result <= 8'b01101001;
   1425: result <= 8'b01101001;
   1426: result <= 8'b01101000;
   1427: result <= 8'b01101000;
   1428: result <= 8'b01101000;
   1429: result <= 8'b01101000;
   1430: result <= 8'b01101000;
   1431: result <= 8'b01101000;
   1432: result <= 8'b01101000;
   1433: result <= 8'b01101000;
   1434: result <= 8'b01101000;
   1435: result <= 8'b01100111;
   1436: result <= 8'b01100111;
   1437: result <= 8'b01100111;
   1438: result <= 8'b01100111;
   1439: result <= 8'b01100111;
   1440: result <= 8'b01100111;
   1441: result <= 8'b01100111;
   1442: result <= 8'b01100111;
   1443: result <= 8'b01100110;
   1444: result <= 8'b01100110;
   1445: result <= 8'b01100110;
   1446: result <= 8'b01100110;
   1447: result <= 8'b01100110;
   1448: result <= 8'b01100110;
   1449: result <= 8'b01100110;
   1450: result <= 8'b01100110;
   1451: result <= 8'b01100110;
   1452: result <= 8'b01100101;
   1453: result <= 8'b01100101;
   1454: result <= 8'b01100101;
   1455: result <= 8'b01100101;
   1456: result <= 8'b01100101;
   1457: result <= 8'b01100101;
   1458: result <= 8'b01100101;
   1459: result <= 8'b01100101;
   1460: result <= 8'b01100100;
   1461: result <= 8'b01100100;
   1462: result <= 8'b01100100;
   1463: result <= 8'b01100100;
   1464: result <= 8'b01100100;
   1465: result <= 8'b01100100;
   1466: result <= 8'b01100100;
   1467: result <= 8'b01100100;
   1468: result <= 8'b01100011;
   1469: result <= 8'b01100011;
   1470: result <= 8'b01100011;
   1471: result <= 8'b01100011;
   1472: result <= 8'b01100011;
   1473: result <= 8'b01100011;
   1474: result <= 8'b01100011;
   1475: result <= 8'b01100011;
   1476: result <= 8'b01100010;
   1477: result <= 8'b01100010;
   1478: result <= 8'b01100010;
   1479: result <= 8'b01100010;
   1480: result <= 8'b01100010;
   1481: result <= 8'b01100010;
   1482: result <= 8'b01100010;
   1483: result <= 8'b01100010;
   1484: result <= 8'b01100001;
   1485: result <= 8'b01100001;
   1486: result <= 8'b01100001;
   1487: result <= 8'b01100001;
   1488: result <= 8'b01100001;
   1489: result <= 8'b01100001;
   1490: result <= 8'b01100001;
   1491: result <= 8'b01100001;
   1492: result <= 8'b01100000;
   1493: result <= 8'b01100000;
   1494: result <= 8'b01100000;
   1495: result <= 8'b01100000;
   1496: result <= 8'b01100000;
   1497: result <= 8'b01100000;
   1498: result <= 8'b01100000;
   1499: result <= 8'b01011111;
   1500: result <= 8'b01011111;
   1501: result <= 8'b01011111;
   1502: result <= 8'b01011111;
   1503: result <= 8'b01011111;
   1504: result <= 8'b01011111;
   1505: result <= 8'b01011111;
   1506: result <= 8'b01011111;
   1507: result <= 8'b01011110;
   1508: result <= 8'b01011110;
   1509: result <= 8'b01011110;
   1510: result <= 8'b01011110;
   1511: result <= 8'b01011110;
   1512: result <= 8'b01011110;
   1513: result <= 8'b01011110;
   1514: result <= 8'b01011110;
   1515: result <= 8'b01011101;
   1516: result <= 8'b01011101;
   1517: result <= 8'b01011101;
   1518: result <= 8'b01011101;
   1519: result <= 8'b01011101;
   1520: result <= 8'b01011101;
   1521: result <= 8'b01011101;
   1522: result <= 8'b01011100;
   1523: result <= 8'b01011100;
   1524: result <= 8'b01011100;
   1525: result <= 8'b01011100;
   1526: result <= 8'b01011100;
   1527: result <= 8'b01011100;
   1528: result <= 8'b01011100;
   1529: result <= 8'b01011011;
   1530: result <= 8'b01011011;
   1531: result <= 8'b01011011;
   1532: result <= 8'b01011011;
   1533: result <= 8'b01011011;
   1534: result <= 8'b01011011;
   1535: result <= 8'b01011011;
   1536: result <= 8'b01011011;
   1537: result <= 8'b01011010;
   1538: result <= 8'b01011010;
   1539: result <= 8'b01011010;
   1540: result <= 8'b01011010;
   1541: result <= 8'b01011010;
   1542: result <= 8'b01011010;
   1543: result <= 8'b01011010;
   1544: result <= 8'b01011001;
   1545: result <= 8'b01011001;
   1546: result <= 8'b01011001;
   1547: result <= 8'b01011001;
   1548: result <= 8'b01011001;
   1549: result <= 8'b01011001;
   1550: result <= 8'b01011001;
   1551: result <= 8'b01011000;
   1552: result <= 8'b01011000;
   1553: result <= 8'b01011000;
   1554: result <= 8'b01011000;
   1555: result <= 8'b01011000;
   1556: result <= 8'b01011000;
   1557: result <= 8'b01011000;
   1558: result <= 8'b01010111;
   1559: result <= 8'b01010111;
   1560: result <= 8'b01010111;
   1561: result <= 8'b01010111;
   1562: result <= 8'b01010111;
   1563: result <= 8'b01010111;
   1564: result <= 8'b01010111;
   1565: result <= 8'b01010110;
   1566: result <= 8'b01010110;
   1567: result <= 8'b01010110;
   1568: result <= 8'b01010110;
   1569: result <= 8'b01010110;
   1570: result <= 8'b01010110;
   1571: result <= 8'b01010110;
   1572: result <= 8'b01010101;
   1573: result <= 8'b01010101;
   1574: result <= 8'b01010101;
   1575: result <= 8'b01010101;
   1576: result <= 8'b01010101;
   1577: result <= 8'b01010101;
   1578: result <= 8'b01010100;
   1579: result <= 8'b01010100;
   1580: result <= 8'b01010100;
   1581: result <= 8'b01010100;
   1582: result <= 8'b01010100;
   1583: result <= 8'b01010100;
   1584: result <= 8'b01010100;
   1585: result <= 8'b01010011;
   1586: result <= 8'b01010011;
   1587: result <= 8'b01010011;
   1588: result <= 8'b01010011;
   1589: result <= 8'b01010011;
   1590: result <= 8'b01010011;
   1591: result <= 8'b01010011;
   1592: result <= 8'b01010010;
   1593: result <= 8'b01010010;
   1594: result <= 8'b01010010;
   1595: result <= 8'b01010010;
   1596: result <= 8'b01010010;
   1597: result <= 8'b01010010;
   1598: result <= 8'b01010010;
   1599: result <= 8'b01010001;
   1600: result <= 8'b01010001;
   1601: result <= 8'b01010001;
   1602: result <= 8'b01010001;
   1603: result <= 8'b01010001;
   1604: result <= 8'b01010001;
   1605: result <= 8'b01010000;
   1606: result <= 8'b01010000;
   1607: result <= 8'b01010000;
   1608: result <= 8'b01010000;
   1609: result <= 8'b01010000;
   1610: result <= 8'b01010000;
   1611: result <= 8'b01010000;
   1612: result <= 8'b01001111;
   1613: result <= 8'b01001111;
   1614: result <= 8'b01001111;
   1615: result <= 8'b01001111;
   1616: result <= 8'b01001111;
   1617: result <= 8'b01001111;
   1618: result <= 8'b01001110;
   1619: result <= 8'b01001110;
   1620: result <= 8'b01001110;
   1621: result <= 8'b01001110;
   1622: result <= 8'b01001110;
   1623: result <= 8'b01001110;
   1624: result <= 8'b01001110;
   1625: result <= 8'b01001101;
   1626: result <= 8'b01001101;
   1627: result <= 8'b01001101;
   1628: result <= 8'b01001101;
   1629: result <= 8'b01001101;
   1630: result <= 8'b01001101;
   1631: result <= 8'b01001100;
   1632: result <= 8'b01001100;
   1633: result <= 8'b01001100;
   1634: result <= 8'b01001100;
   1635: result <= 8'b01001100;
   1636: result <= 8'b01001100;
   1637: result <= 8'b01001011;
   1638: result <= 8'b01001011;
   1639: result <= 8'b01001011;
   1640: result <= 8'b01001011;
   1641: result <= 8'b01001011;
   1642: result <= 8'b01001011;
   1643: result <= 8'b01001011;
   1644: result <= 8'b01001010;
   1645: result <= 8'b01001010;
   1646: result <= 8'b01001010;
   1647: result <= 8'b01001010;
   1648: result <= 8'b01001010;
   1649: result <= 8'b01001010;
   1650: result <= 8'b01001001;
   1651: result <= 8'b01001001;
   1652: result <= 8'b01001001;
   1653: result <= 8'b01001001;
   1654: result <= 8'b01001001;
   1655: result <= 8'b01001001;
   1656: result <= 8'b01001000;
   1657: result <= 8'b01001000;
   1658: result <= 8'b01001000;
   1659: result <= 8'b01001000;
   1660: result <= 8'b01001000;
   1661: result <= 8'b01001000;
   1662: result <= 8'b01000111;
   1663: result <= 8'b01000111;
   1664: result <= 8'b01000111;
   1665: result <= 8'b01000111;
   1666: result <= 8'b01000111;
   1667: result <= 8'b01000111;
   1668: result <= 8'b01000110;
   1669: result <= 8'b01000110;
   1670: result <= 8'b01000110;
   1671: result <= 8'b01000110;
   1672: result <= 8'b01000110;
   1673: result <= 8'b01000110;
   1674: result <= 8'b01000101;
   1675: result <= 8'b01000101;
   1676: result <= 8'b01000101;
   1677: result <= 8'b01000101;
   1678: result <= 8'b01000101;
   1679: result <= 8'b01000101;
   1680: result <= 8'b01000100;
   1681: result <= 8'b01000100;
   1682: result <= 8'b01000100;
   1683: result <= 8'b01000100;
   1684: result <= 8'b01000100;
   1685: result <= 8'b01000100;
   1686: result <= 8'b01000011;
   1687: result <= 8'b01000011;
   1688: result <= 8'b01000011;
   1689: result <= 8'b01000011;
   1690: result <= 8'b01000011;
   1691: result <= 8'b01000011;
   1692: result <= 8'b01000010;
   1693: result <= 8'b01000010;
   1694: result <= 8'b01000010;
   1695: result <= 8'b01000010;
   1696: result <= 8'b01000010;
   1697: result <= 8'b01000010;
   1698: result <= 8'b01000001;
   1699: result <= 8'b01000001;
   1700: result <= 8'b01000001;
   1701: result <= 8'b01000001;
   1702: result <= 8'b01000001;
   1703: result <= 8'b01000001;
   1704: result <= 8'b01000000;
   1705: result <= 8'b01000000;
   1706: result <= 8'b01000000;
   1707: result <= 8'b01000000;
   1708: result <= 8'b01000000;
   1709: result <= 8'b01000000;
   1710: result <= 8'b00111111;
   1711: result <= 8'b00111111;
   1712: result <= 8'b00111111;
   1713: result <= 8'b00111111;
   1714: result <= 8'b00111111;
   1715: result <= 8'b00111111;
   1716: result <= 8'b00111110;
   1717: result <= 8'b00111110;
   1718: result <= 8'b00111110;
   1719: result <= 8'b00111110;
   1720: result <= 8'b00111110;
   1721: result <= 8'b00111110;
   1722: result <= 8'b00111101;
   1723: result <= 8'b00111101;
   1724: result <= 8'b00111101;
   1725: result <= 8'b00111101;
   1726: result <= 8'b00111101;
   1727: result <= 8'b00111101;
   1728: result <= 8'b00111100;
   1729: result <= 8'b00111100;
   1730: result <= 8'b00111100;
   1731: result <= 8'b00111100;
   1732: result <= 8'b00111100;
   1733: result <= 8'b00111011;
   1734: result <= 8'b00111011;
   1735: result <= 8'b00111011;
   1736: result <= 8'b00111011;
   1737: result <= 8'b00111011;
   1738: result <= 8'b00111011;
   1739: result <= 8'b00111010;
   1740: result <= 8'b00111010;
   1741: result <= 8'b00111010;
   1742: result <= 8'b00111010;
   1743: result <= 8'b00111010;
   1744: result <= 8'b00111010;
   1745: result <= 8'b00111001;
   1746: result <= 8'b00111001;
   1747: result <= 8'b00111001;
   1748: result <= 8'b00111001;
   1749: result <= 8'b00111001;
   1750: result <= 8'b00111000;
   1751: result <= 8'b00111000;
   1752: result <= 8'b00111000;
   1753: result <= 8'b00111000;
   1754: result <= 8'b00111000;
   1755: result <= 8'b00111000;
   1756: result <= 8'b00110111;
   1757: result <= 8'b00110111;
   1758: result <= 8'b00110111;
   1759: result <= 8'b00110111;
   1760: result <= 8'b00110111;
   1761: result <= 8'b00110111;
   1762: result <= 8'b00110110;
   1763: result <= 8'b00110110;
   1764: result <= 8'b00110110;
   1765: result <= 8'b00110110;
   1766: result <= 8'b00110110;
   1767: result <= 8'b00110101;
   1768: result <= 8'b00110101;
   1769: result <= 8'b00110101;
   1770: result <= 8'b00110101;
   1771: result <= 8'b00110101;
   1772: result <= 8'b00110101;
   1773: result <= 8'b00110100;
   1774: result <= 8'b00110100;
   1775: result <= 8'b00110100;
   1776: result <= 8'b00110100;
   1777: result <= 8'b00110100;
   1778: result <= 8'b00110100;
   1779: result <= 8'b00110011;
   1780: result <= 8'b00110011;
   1781: result <= 8'b00110011;
   1782: result <= 8'b00110011;
   1783: result <= 8'b00110011;
   1784: result <= 8'b00110010;
   1785: result <= 8'b00110010;
   1786: result <= 8'b00110010;
   1787: result <= 8'b00110010;
   1788: result <= 8'b00110010;
   1789: result <= 8'b00110010;
   1790: result <= 8'b00110001;
   1791: result <= 8'b00110001;
   1792: result <= 8'b00110001;
   1793: result <= 8'b00110001;
   1794: result <= 8'b00110001;
   1795: result <= 8'b00110000;
   1796: result <= 8'b00110000;
   1797: result <= 8'b00110000;
   1798: result <= 8'b00110000;
   1799: result <= 8'b00110000;
   1800: result <= 8'b00110000;
   1801: result <= 8'b00101111;
   1802: result <= 8'b00101111;
   1803: result <= 8'b00101111;
   1804: result <= 8'b00101111;
   1805: result <= 8'b00101111;
   1806: result <= 8'b00101110;
   1807: result <= 8'b00101110;
   1808: result <= 8'b00101110;
   1809: result <= 8'b00101110;
   1810: result <= 8'b00101110;
   1811: result <= 8'b00101110;
   1812: result <= 8'b00101101;
   1813: result <= 8'b00101101;
   1814: result <= 8'b00101101;
   1815: result <= 8'b00101101;
   1816: result <= 8'b00101101;
   1817: result <= 8'b00101100;
   1818: result <= 8'b00101100;
   1819: result <= 8'b00101100;
   1820: result <= 8'b00101100;
   1821: result <= 8'b00101100;
   1822: result <= 8'b00101011;
   1823: result <= 8'b00101011;
   1824: result <= 8'b00101011;
   1825: result <= 8'b00101011;
   1826: result <= 8'b00101011;
   1827: result <= 8'b00101011;
   1828: result <= 8'b00101010;
   1829: result <= 8'b00101010;
   1830: result <= 8'b00101010;
   1831: result <= 8'b00101010;
   1832: result <= 8'b00101010;
   1833: result <= 8'b00101001;
   1834: result <= 8'b00101001;
   1835: result <= 8'b00101001;
   1836: result <= 8'b00101001;
   1837: result <= 8'b00101001;
   1838: result <= 8'b00101001;
   1839: result <= 8'b00101000;
   1840: result <= 8'b00101000;
   1841: result <= 8'b00101000;
   1842: result <= 8'b00101000;
   1843: result <= 8'b00101000;
   1844: result <= 8'b00100111;
   1845: result <= 8'b00100111;
   1846: result <= 8'b00100111;
   1847: result <= 8'b00100111;
   1848: result <= 8'b00100111;
   1849: result <= 8'b00100110;
   1850: result <= 8'b00100110;
   1851: result <= 8'b00100110;
   1852: result <= 8'b00100110;
   1853: result <= 8'b00100110;
   1854: result <= 8'b00100110;
   1855: result <= 8'b00100101;
   1856: result <= 8'b00100101;
   1857: result <= 8'b00100101;
   1858: result <= 8'b00100101;
   1859: result <= 8'b00100101;
   1860: result <= 8'b00100100;
   1861: result <= 8'b00100100;
   1862: result <= 8'b00100100;
   1863: result <= 8'b00100100;
   1864: result <= 8'b00100100;
   1865: result <= 8'b00100011;
   1866: result <= 8'b00100011;
   1867: result <= 8'b00100011;
   1868: result <= 8'b00100011;
   1869: result <= 8'b00100011;
   1870: result <= 8'b00100011;
   1871: result <= 8'b00100010;
   1872: result <= 8'b00100010;
   1873: result <= 8'b00100010;
   1874: result <= 8'b00100010;
   1875: result <= 8'b00100010;
   1876: result <= 8'b00100001;
   1877: result <= 8'b00100001;
   1878: result <= 8'b00100001;
   1879: result <= 8'b00100001;
   1880: result <= 8'b00100001;
   1881: result <= 8'b00100000;
   1882: result <= 8'b00100000;
   1883: result <= 8'b00100000;
   1884: result <= 8'b00100000;
   1885: result <= 8'b00100000;
   1886: result <= 8'b00011111;
   1887: result <= 8'b00011111;
   1888: result <= 8'b00011111;
   1889: result <= 8'b00011111;
   1890: result <= 8'b00011111;
   1891: result <= 8'b00011111;
   1892: result <= 8'b00011110;
   1893: result <= 8'b00011110;
   1894: result <= 8'b00011110;
   1895: result <= 8'b00011110;
   1896: result <= 8'b00011110;
   1897: result <= 8'b00011101;
   1898: result <= 8'b00011101;
   1899: result <= 8'b00011101;
   1900: result <= 8'b00011101;
   1901: result <= 8'b00011101;
   1902: result <= 8'b00011100;
   1903: result <= 8'b00011100;
   1904: result <= 8'b00011100;
   1905: result <= 8'b00011100;
   1906: result <= 8'b00011100;
   1907: result <= 8'b00011011;
   1908: result <= 8'b00011011;
   1909: result <= 8'b00011011;
   1910: result <= 8'b00011011;
   1911: result <= 8'b00011011;
   1912: result <= 8'b00011011;
   1913: result <= 8'b00011010;
   1914: result <= 8'b00011010;
   1915: result <= 8'b00011010;
   1916: result <= 8'b00011010;
   1917: result <= 8'b00011010;
   1918: result <= 8'b00011001;
   1919: result <= 8'b00011001;
   1920: result <= 8'b00011001;
   1921: result <= 8'b00011001;
   1922: result <= 8'b00011001;
   1923: result <= 8'b00011000;
   1924: result <= 8'b00011000;
   1925: result <= 8'b00011000;
   1926: result <= 8'b00011000;
   1927: result <= 8'b00011000;
   1928: result <= 8'b00010111;
   1929: result <= 8'b00010111;
   1930: result <= 8'b00010111;
   1931: result <= 8'b00010111;
   1932: result <= 8'b00010111;
   1933: result <= 8'b00010110;
   1934: result <= 8'b00010110;
   1935: result <= 8'b00010110;
   1936: result <= 8'b00010110;
   1937: result <= 8'b00010110;
   1938: result <= 8'b00010101;
   1939: result <= 8'b00010101;
   1940: result <= 8'b00010101;
   1941: result <= 8'b00010101;
   1942: result <= 8'b00010101;
   1943: result <= 8'b00010101;
   1944: result <= 8'b00010100;
   1945: result <= 8'b00010100;
   1946: result <= 8'b00010100;
   1947: result <= 8'b00010100;
   1948: result <= 8'b00010100;
   1949: result <= 8'b00010011;
   1950: result <= 8'b00010011;
   1951: result <= 8'b00010011;
   1952: result <= 8'b00010011;
   1953: result <= 8'b00010011;
   1954: result <= 8'b00010010;
   1955: result <= 8'b00010010;
   1956: result <= 8'b00010010;
   1957: result <= 8'b00010010;
   1958: result <= 8'b00010010;
   1959: result <= 8'b00010001;
   1960: result <= 8'b00010001;
   1961: result <= 8'b00010001;
   1962: result <= 8'b00010001;
   1963: result <= 8'b00010001;
   1964: result <= 8'b00010000;
   1965: result <= 8'b00010000;
   1966: result <= 8'b00010000;
   1967: result <= 8'b00010000;
   1968: result <= 8'b00010000;
   1969: result <= 8'b00001111;
   1970: result <= 8'b00001111;
   1971: result <= 8'b00001111;
   1972: result <= 8'b00001111;
   1973: result <= 8'b00001111;
   1974: result <= 8'b00001110;
   1975: result <= 8'b00001110;
   1976: result <= 8'b00001110;
   1977: result <= 8'b00001110;
   1978: result <= 8'b00001110;
   1979: result <= 8'b00001110;
   1980: result <= 8'b00001101;
   1981: result <= 8'b00001101;
   1982: result <= 8'b00001101;
   1983: result <= 8'b00001101;
   1984: result <= 8'b00001101;
   1985: result <= 8'b00001100;
   1986: result <= 8'b00001100;
   1987: result <= 8'b00001100;
   1988: result <= 8'b00001100;
   1989: result <= 8'b00001100;
   1990: result <= 8'b00001011;
   1991: result <= 8'b00001011;
   1992: result <= 8'b00001011;
   1993: result <= 8'b00001011;
   1994: result <= 8'b00001011;
   1995: result <= 8'b00001010;
   1996: result <= 8'b00001010;
   1997: result <= 8'b00001010;
   1998: result <= 8'b00001010;
   1999: result <= 8'b00001010;
   2000: result <= 8'b00001001;
   2001: result <= 8'b00001001;
   2002: result <= 8'b00001001;
   2003: result <= 8'b00001001;
   2004: result <= 8'b00001001;
   2005: result <= 8'b00001000;
   2006: result <= 8'b00001000;
   2007: result <= 8'b00001000;
   2008: result <= 8'b00001000;
   2009: result <= 8'b00001000;
   2010: result <= 8'b00000111;
   2011: result <= 8'b00000111;
   2012: result <= 8'b00000111;
   2013: result <= 8'b00000111;
   2014: result <= 8'b00000111;
   2015: result <= 8'b00000110;
   2016: result <= 8'b00000110;
   2017: result <= 8'b00000110;
   2018: result <= 8'b00000110;
   2019: result <= 8'b00000110;
   2020: result <= 8'b00000101;
   2021: result <= 8'b00000101;
   2022: result <= 8'b00000101;
   2023: result <= 8'b00000101;
   2024: result <= 8'b00000101;
   2025: result <= 8'b00000101;
   2026: result <= 8'b00000100;
   2027: result <= 8'b00000100;
   2028: result <= 8'b00000100;
   2029: result <= 8'b00000100;
   2030: result <= 8'b00000100;
   2031: result <= 8'b00000011;
   2032: result <= 8'b00000011;
   2033: result <= 8'b00000011;
   2034: result <= 8'b00000011;
   2035: result <= 8'b00000011;
   2036: result <= 8'b00000010;
   2037: result <= 8'b00000010;
   2038: result <= 8'b00000010;
   2039: result <= 8'b00000010;
   2040: result <= 8'b00000010;
   2041: result <= 8'b00000001;
   2042: result <= 8'b00000001;
   2043: result <= 8'b00000001;
   2044: result <= 8'b00000001;
   2045: result <= 8'b00000001;
   2046: result <= 8'b00000000;
   2047: result <= 8'b00000000;
   2048: result <= 8'b00000000;
   2049: result <= 8'b00000000;
   2050: result <= 8'b00000000;
   2051: result <= 8'b11111111;
   2052: result <= 8'b11111111;
   2053: result <= 8'b11111111;
   2054: result <= 8'b11111111;
   2055: result <= 8'b11111111;
   2056: result <= 8'b11111110;
   2057: result <= 8'b11111110;
   2058: result <= 8'b11111110;
   2059: result <= 8'b11111110;
   2060: result <= 8'b11111110;
   2061: result <= 8'b11111101;
   2062: result <= 8'b11111101;
   2063: result <= 8'b11111101;
   2064: result <= 8'b11111101;
   2065: result <= 8'b11111101;
   2066: result <= 8'b11111100;
   2067: result <= 8'b11111100;
   2068: result <= 8'b11111100;
   2069: result <= 8'b11111100;
   2070: result <= 8'b11111100;
   2071: result <= 8'b11111011;
   2072: result <= 8'b11111011;
   2073: result <= 8'b11111011;
   2074: result <= 8'b11111011;
   2075: result <= 8'b11111011;
   2076: result <= 8'b11111011;
   2077: result <= 8'b11111010;
   2078: result <= 8'b11111010;
   2079: result <= 8'b11111010;
   2080: result <= 8'b11111010;
   2081: result <= 8'b11111010;
   2082: result <= 8'b11111001;
   2083: result <= 8'b11111001;
   2084: result <= 8'b11111001;
   2085: result <= 8'b11111001;
   2086: result <= 8'b11111001;
   2087: result <= 8'b11111000;
   2088: result <= 8'b11111000;
   2089: result <= 8'b11111000;
   2090: result <= 8'b11111000;
   2091: result <= 8'b11111000;
   2092: result <= 8'b11110111;
   2093: result <= 8'b11110111;
   2094: result <= 8'b11110111;
   2095: result <= 8'b11110111;
   2096: result <= 8'b11110111;
   2097: result <= 8'b11110110;
   2098: result <= 8'b11110110;
   2099: result <= 8'b11110110;
   2100: result <= 8'b11110110;
   2101: result <= 8'b11110110;
   2102: result <= 8'b11110101;
   2103: result <= 8'b11110101;
   2104: result <= 8'b11110101;
   2105: result <= 8'b11110101;
   2106: result <= 8'b11110101;
   2107: result <= 8'b11110100;
   2108: result <= 8'b11110100;
   2109: result <= 8'b11110100;
   2110: result <= 8'b11110100;
   2111: result <= 8'b11110100;
   2112: result <= 8'b11110011;
   2113: result <= 8'b11110011;
   2114: result <= 8'b11110011;
   2115: result <= 8'b11110011;
   2116: result <= 8'b11110011;
   2117: result <= 8'b11110010;
   2118: result <= 8'b11110010;
   2119: result <= 8'b11110010;
   2120: result <= 8'b11110010;
   2121: result <= 8'b11110010;
   2122: result <= 8'b11110010;
   2123: result <= 8'b11110001;
   2124: result <= 8'b11110001;
   2125: result <= 8'b11110001;
   2126: result <= 8'b11110001;
   2127: result <= 8'b11110001;
   2128: result <= 8'b11110000;
   2129: result <= 8'b11110000;
   2130: result <= 8'b11110000;
   2131: result <= 8'b11110000;
   2132: result <= 8'b11110000;
   2133: result <= 8'b11101111;
   2134: result <= 8'b11101111;
   2135: result <= 8'b11101111;
   2136: result <= 8'b11101111;
   2137: result <= 8'b11101111;
   2138: result <= 8'b11101110;
   2139: result <= 8'b11101110;
   2140: result <= 8'b11101110;
   2141: result <= 8'b11101110;
   2142: result <= 8'b11101110;
   2143: result <= 8'b11101101;
   2144: result <= 8'b11101101;
   2145: result <= 8'b11101101;
   2146: result <= 8'b11101101;
   2147: result <= 8'b11101101;
   2148: result <= 8'b11101100;
   2149: result <= 8'b11101100;
   2150: result <= 8'b11101100;
   2151: result <= 8'b11101100;
   2152: result <= 8'b11101100;
   2153: result <= 8'b11101011;
   2154: result <= 8'b11101011;
   2155: result <= 8'b11101011;
   2156: result <= 8'b11101011;
   2157: result <= 8'b11101011;
   2158: result <= 8'b11101011;
   2159: result <= 8'b11101010;
   2160: result <= 8'b11101010;
   2161: result <= 8'b11101010;
   2162: result <= 8'b11101010;
   2163: result <= 8'b11101010;
   2164: result <= 8'b11101001;
   2165: result <= 8'b11101001;
   2166: result <= 8'b11101001;
   2167: result <= 8'b11101001;
   2168: result <= 8'b11101001;
   2169: result <= 8'b11101000;
   2170: result <= 8'b11101000;
   2171: result <= 8'b11101000;
   2172: result <= 8'b11101000;
   2173: result <= 8'b11101000;
   2174: result <= 8'b11100111;
   2175: result <= 8'b11100111;
   2176: result <= 8'b11100111;
   2177: result <= 8'b11100111;
   2178: result <= 8'b11100111;
   2179: result <= 8'b11100110;
   2180: result <= 8'b11100110;
   2181: result <= 8'b11100110;
   2182: result <= 8'b11100110;
   2183: result <= 8'b11100110;
   2184: result <= 8'b11100101;
   2185: result <= 8'b11100101;
   2186: result <= 8'b11100101;
   2187: result <= 8'b11100101;
   2188: result <= 8'b11100101;
   2189: result <= 8'b11100101;
   2190: result <= 8'b11100100;
   2191: result <= 8'b11100100;
   2192: result <= 8'b11100100;
   2193: result <= 8'b11100100;
   2194: result <= 8'b11100100;
   2195: result <= 8'b11100011;
   2196: result <= 8'b11100011;
   2197: result <= 8'b11100011;
   2198: result <= 8'b11100011;
   2199: result <= 8'b11100011;
   2200: result <= 8'b11100010;
   2201: result <= 8'b11100010;
   2202: result <= 8'b11100010;
   2203: result <= 8'b11100010;
   2204: result <= 8'b11100010;
   2205: result <= 8'b11100001;
   2206: result <= 8'b11100001;
   2207: result <= 8'b11100001;
   2208: result <= 8'b11100001;
   2209: result <= 8'b11100001;
   2210: result <= 8'b11100001;
   2211: result <= 8'b11100000;
   2212: result <= 8'b11100000;
   2213: result <= 8'b11100000;
   2214: result <= 8'b11100000;
   2215: result <= 8'b11100000;
   2216: result <= 8'b11011111;
   2217: result <= 8'b11011111;
   2218: result <= 8'b11011111;
   2219: result <= 8'b11011111;
   2220: result <= 8'b11011111;
   2221: result <= 8'b11011110;
   2222: result <= 8'b11011110;
   2223: result <= 8'b11011110;
   2224: result <= 8'b11011110;
   2225: result <= 8'b11011110;
   2226: result <= 8'b11011101;
   2227: result <= 8'b11011101;
   2228: result <= 8'b11011101;
   2229: result <= 8'b11011101;
   2230: result <= 8'b11011101;
   2231: result <= 8'b11011101;
   2232: result <= 8'b11011100;
   2233: result <= 8'b11011100;
   2234: result <= 8'b11011100;
   2235: result <= 8'b11011100;
   2236: result <= 8'b11011100;
   2237: result <= 8'b11011011;
   2238: result <= 8'b11011011;
   2239: result <= 8'b11011011;
   2240: result <= 8'b11011011;
   2241: result <= 8'b11011011;
   2242: result <= 8'b11011010;
   2243: result <= 8'b11011010;
   2244: result <= 8'b11011010;
   2245: result <= 8'b11011010;
   2246: result <= 8'b11011010;
   2247: result <= 8'b11011010;
   2248: result <= 8'b11011001;
   2249: result <= 8'b11011001;
   2250: result <= 8'b11011001;
   2251: result <= 8'b11011001;
   2252: result <= 8'b11011001;
   2253: result <= 8'b11011000;
   2254: result <= 8'b11011000;
   2255: result <= 8'b11011000;
   2256: result <= 8'b11011000;
   2257: result <= 8'b11011000;
   2258: result <= 8'b11010111;
   2259: result <= 8'b11010111;
   2260: result <= 8'b11010111;
   2261: result <= 8'b11010111;
   2262: result <= 8'b11010111;
   2263: result <= 8'b11010111;
   2264: result <= 8'b11010110;
   2265: result <= 8'b11010110;
   2266: result <= 8'b11010110;
   2267: result <= 8'b11010110;
   2268: result <= 8'b11010110;
   2269: result <= 8'b11010101;
   2270: result <= 8'b11010101;
   2271: result <= 8'b11010101;
   2272: result <= 8'b11010101;
   2273: result <= 8'b11010101;
   2274: result <= 8'b11010101;
   2275: result <= 8'b11010100;
   2276: result <= 8'b11010100;
   2277: result <= 8'b11010100;
   2278: result <= 8'b11010100;
   2279: result <= 8'b11010100;
   2280: result <= 8'b11010011;
   2281: result <= 8'b11010011;
   2282: result <= 8'b11010011;
   2283: result <= 8'b11010011;
   2284: result <= 8'b11010011;
   2285: result <= 8'b11010010;
   2286: result <= 8'b11010010;
   2287: result <= 8'b11010010;
   2288: result <= 8'b11010010;
   2289: result <= 8'b11010010;
   2290: result <= 8'b11010010;
   2291: result <= 8'b11010001;
   2292: result <= 8'b11010001;
   2293: result <= 8'b11010001;
   2294: result <= 8'b11010001;
   2295: result <= 8'b11010001;
   2296: result <= 8'b11010000;
   2297: result <= 8'b11010000;
   2298: result <= 8'b11010000;
   2299: result <= 8'b11010000;
   2300: result <= 8'b11010000;
   2301: result <= 8'b11010000;
   2302: result <= 8'b11001111;
   2303: result <= 8'b11001111;
   2304: result <= 8'b11001111;
   2305: result <= 8'b11001111;
   2306: result <= 8'b11001111;
   2307: result <= 8'b11001110;
   2308: result <= 8'b11001110;
   2309: result <= 8'b11001110;
   2310: result <= 8'b11001110;
   2311: result <= 8'b11001110;
   2312: result <= 8'b11001110;
   2313: result <= 8'b11001101;
   2314: result <= 8'b11001101;
   2315: result <= 8'b11001101;
   2316: result <= 8'b11001101;
   2317: result <= 8'b11001101;
   2318: result <= 8'b11001100;
   2319: result <= 8'b11001100;
   2320: result <= 8'b11001100;
   2321: result <= 8'b11001100;
   2322: result <= 8'b11001100;
   2323: result <= 8'b11001100;
   2324: result <= 8'b11001011;
   2325: result <= 8'b11001011;
   2326: result <= 8'b11001011;
   2327: result <= 8'b11001011;
   2328: result <= 8'b11001011;
   2329: result <= 8'b11001011;
   2330: result <= 8'b11001010;
   2331: result <= 8'b11001010;
   2332: result <= 8'b11001010;
   2333: result <= 8'b11001010;
   2334: result <= 8'b11001010;
   2335: result <= 8'b11001001;
   2336: result <= 8'b11001001;
   2337: result <= 8'b11001001;
   2338: result <= 8'b11001001;
   2339: result <= 8'b11001001;
   2340: result <= 8'b11001001;
   2341: result <= 8'b11001000;
   2342: result <= 8'b11001000;
   2343: result <= 8'b11001000;
   2344: result <= 8'b11001000;
   2345: result <= 8'b11001000;
   2346: result <= 8'b11001000;
   2347: result <= 8'b11000111;
   2348: result <= 8'b11000111;
   2349: result <= 8'b11000111;
   2350: result <= 8'b11000111;
   2351: result <= 8'b11000111;
   2352: result <= 8'b11000110;
   2353: result <= 8'b11000110;
   2354: result <= 8'b11000110;
   2355: result <= 8'b11000110;
   2356: result <= 8'b11000110;
   2357: result <= 8'b11000110;
   2358: result <= 8'b11000101;
   2359: result <= 8'b11000101;
   2360: result <= 8'b11000101;
   2361: result <= 8'b11000101;
   2362: result <= 8'b11000101;
   2363: result <= 8'b11000101;
   2364: result <= 8'b11000100;
   2365: result <= 8'b11000100;
   2366: result <= 8'b11000100;
   2367: result <= 8'b11000100;
   2368: result <= 8'b11000100;
   2369: result <= 8'b11000011;
   2370: result <= 8'b11000011;
   2371: result <= 8'b11000011;
   2372: result <= 8'b11000011;
   2373: result <= 8'b11000011;
   2374: result <= 8'b11000011;
   2375: result <= 8'b11000010;
   2376: result <= 8'b11000010;
   2377: result <= 8'b11000010;
   2378: result <= 8'b11000010;
   2379: result <= 8'b11000010;
   2380: result <= 8'b11000010;
   2381: result <= 8'b11000001;
   2382: result <= 8'b11000001;
   2383: result <= 8'b11000001;
   2384: result <= 8'b11000001;
   2385: result <= 8'b11000001;
   2386: result <= 8'b11000001;
   2387: result <= 8'b11000000;
   2388: result <= 8'b11000000;
   2389: result <= 8'b11000000;
   2390: result <= 8'b11000000;
   2391: result <= 8'b11000000;
   2392: result <= 8'b11000000;
   2393: result <= 8'b10111111;
   2394: result <= 8'b10111111;
   2395: result <= 8'b10111111;
   2396: result <= 8'b10111111;
   2397: result <= 8'b10111111;
   2398: result <= 8'b10111111;
   2399: result <= 8'b10111110;
   2400: result <= 8'b10111110;
   2401: result <= 8'b10111110;
   2402: result <= 8'b10111110;
   2403: result <= 8'b10111110;
   2404: result <= 8'b10111110;
   2405: result <= 8'b10111101;
   2406: result <= 8'b10111101;
   2407: result <= 8'b10111101;
   2408: result <= 8'b10111101;
   2409: result <= 8'b10111101;
   2410: result <= 8'b10111101;
   2411: result <= 8'b10111100;
   2412: result <= 8'b10111100;
   2413: result <= 8'b10111100;
   2414: result <= 8'b10111100;
   2415: result <= 8'b10111100;
   2416: result <= 8'b10111100;
   2417: result <= 8'b10111011;
   2418: result <= 8'b10111011;
   2419: result <= 8'b10111011;
   2420: result <= 8'b10111011;
   2421: result <= 8'b10111011;
   2422: result <= 8'b10111011;
   2423: result <= 8'b10111010;
   2424: result <= 8'b10111010;
   2425: result <= 8'b10111010;
   2426: result <= 8'b10111010;
   2427: result <= 8'b10111010;
   2428: result <= 8'b10111010;
   2429: result <= 8'b10111001;
   2430: result <= 8'b10111001;
   2431: result <= 8'b10111001;
   2432: result <= 8'b10111001;
   2433: result <= 8'b10111001;
   2434: result <= 8'b10111001;
   2435: result <= 8'b10111000;
   2436: result <= 8'b10111000;
   2437: result <= 8'b10111000;
   2438: result <= 8'b10111000;
   2439: result <= 8'b10111000;
   2440: result <= 8'b10111000;
   2441: result <= 8'b10110111;
   2442: result <= 8'b10110111;
   2443: result <= 8'b10110111;
   2444: result <= 8'b10110111;
   2445: result <= 8'b10110111;
   2446: result <= 8'b10110111;
   2447: result <= 8'b10110110;
   2448: result <= 8'b10110110;
   2449: result <= 8'b10110110;
   2450: result <= 8'b10110110;
   2451: result <= 8'b10110110;
   2452: result <= 8'b10110110;
   2453: result <= 8'b10110101;
   2454: result <= 8'b10110101;
   2455: result <= 8'b10110101;
   2456: result <= 8'b10110101;
   2457: result <= 8'b10110101;
   2458: result <= 8'b10110101;
   2459: result <= 8'b10110101;
   2460: result <= 8'b10110100;
   2461: result <= 8'b10110100;
   2462: result <= 8'b10110100;
   2463: result <= 8'b10110100;
   2464: result <= 8'b10110100;
   2465: result <= 8'b10110100;
   2466: result <= 8'b10110011;
   2467: result <= 8'b10110011;
   2468: result <= 8'b10110011;
   2469: result <= 8'b10110011;
   2470: result <= 8'b10110011;
   2471: result <= 8'b10110011;
   2472: result <= 8'b10110010;
   2473: result <= 8'b10110010;
   2474: result <= 8'b10110010;
   2475: result <= 8'b10110010;
   2476: result <= 8'b10110010;
   2477: result <= 8'b10110010;
   2478: result <= 8'b10110010;
   2479: result <= 8'b10110001;
   2480: result <= 8'b10110001;
   2481: result <= 8'b10110001;
   2482: result <= 8'b10110001;
   2483: result <= 8'b10110001;
   2484: result <= 8'b10110001;
   2485: result <= 8'b10110000;
   2486: result <= 8'b10110000;
   2487: result <= 8'b10110000;
   2488: result <= 8'b10110000;
   2489: result <= 8'b10110000;
   2490: result <= 8'b10110000;
   2491: result <= 8'b10110000;
   2492: result <= 8'b10101111;
   2493: result <= 8'b10101111;
   2494: result <= 8'b10101111;
   2495: result <= 8'b10101111;
   2496: result <= 8'b10101111;
   2497: result <= 8'b10101111;
   2498: result <= 8'b10101110;
   2499: result <= 8'b10101110;
   2500: result <= 8'b10101110;
   2501: result <= 8'b10101110;
   2502: result <= 8'b10101110;
   2503: result <= 8'b10101110;
   2504: result <= 8'b10101110;
   2505: result <= 8'b10101101;
   2506: result <= 8'b10101101;
   2507: result <= 8'b10101101;
   2508: result <= 8'b10101101;
   2509: result <= 8'b10101101;
   2510: result <= 8'b10101101;
   2511: result <= 8'b10101101;
   2512: result <= 8'b10101100;
   2513: result <= 8'b10101100;
   2514: result <= 8'b10101100;
   2515: result <= 8'b10101100;
   2516: result <= 8'b10101100;
   2517: result <= 8'b10101100;
   2518: result <= 8'b10101100;
   2519: result <= 8'b10101011;
   2520: result <= 8'b10101011;
   2521: result <= 8'b10101011;
   2522: result <= 8'b10101011;
   2523: result <= 8'b10101011;
   2524: result <= 8'b10101011;
   2525: result <= 8'b10101010;
   2526: result <= 8'b10101010;
   2527: result <= 8'b10101010;
   2528: result <= 8'b10101010;
   2529: result <= 8'b10101010;
   2530: result <= 8'b10101010;
   2531: result <= 8'b10101010;
   2532: result <= 8'b10101001;
   2533: result <= 8'b10101001;
   2534: result <= 8'b10101001;
   2535: result <= 8'b10101001;
   2536: result <= 8'b10101001;
   2537: result <= 8'b10101001;
   2538: result <= 8'b10101001;
   2539: result <= 8'b10101000;
   2540: result <= 8'b10101000;
   2541: result <= 8'b10101000;
   2542: result <= 8'b10101000;
   2543: result <= 8'b10101000;
   2544: result <= 8'b10101000;
   2545: result <= 8'b10101000;
   2546: result <= 8'b10100111;
   2547: result <= 8'b10100111;
   2548: result <= 8'b10100111;
   2549: result <= 8'b10100111;
   2550: result <= 8'b10100111;
   2551: result <= 8'b10100111;
   2552: result <= 8'b10100111;
   2553: result <= 8'b10100110;
   2554: result <= 8'b10100110;
   2555: result <= 8'b10100110;
   2556: result <= 8'b10100110;
   2557: result <= 8'b10100110;
   2558: result <= 8'b10100110;
   2559: result <= 8'b10100110;
   2560: result <= 8'b10100101;
   2561: result <= 8'b10100101;
   2562: result <= 8'b10100101;
   2563: result <= 8'b10100101;
   2564: result <= 8'b10100101;
   2565: result <= 8'b10100101;
   2566: result <= 8'b10100101;
   2567: result <= 8'b10100101;
   2568: result <= 8'b10100100;
   2569: result <= 8'b10100100;
   2570: result <= 8'b10100100;
   2571: result <= 8'b10100100;
   2572: result <= 8'b10100100;
   2573: result <= 8'b10100100;
   2574: result <= 8'b10100100;
   2575: result <= 8'b10100011;
   2576: result <= 8'b10100011;
   2577: result <= 8'b10100011;
   2578: result <= 8'b10100011;
   2579: result <= 8'b10100011;
   2580: result <= 8'b10100011;
   2581: result <= 8'b10100011;
   2582: result <= 8'b10100010;
   2583: result <= 8'b10100010;
   2584: result <= 8'b10100010;
   2585: result <= 8'b10100010;
   2586: result <= 8'b10100010;
   2587: result <= 8'b10100010;
   2588: result <= 8'b10100010;
   2589: result <= 8'b10100010;
   2590: result <= 8'b10100001;
   2591: result <= 8'b10100001;
   2592: result <= 8'b10100001;
   2593: result <= 8'b10100001;
   2594: result <= 8'b10100001;
   2595: result <= 8'b10100001;
   2596: result <= 8'b10100001;
   2597: result <= 8'b10100001;
   2598: result <= 8'b10100000;
   2599: result <= 8'b10100000;
   2600: result <= 8'b10100000;
   2601: result <= 8'b10100000;
   2602: result <= 8'b10100000;
   2603: result <= 8'b10100000;
   2604: result <= 8'b10100000;
   2605: result <= 8'b10011111;
   2606: result <= 8'b10011111;
   2607: result <= 8'b10011111;
   2608: result <= 8'b10011111;
   2609: result <= 8'b10011111;
   2610: result <= 8'b10011111;
   2611: result <= 8'b10011111;
   2612: result <= 8'b10011111;
   2613: result <= 8'b10011110;
   2614: result <= 8'b10011110;
   2615: result <= 8'b10011110;
   2616: result <= 8'b10011110;
   2617: result <= 8'b10011110;
   2618: result <= 8'b10011110;
   2619: result <= 8'b10011110;
   2620: result <= 8'b10011110;
   2621: result <= 8'b10011101;
   2622: result <= 8'b10011101;
   2623: result <= 8'b10011101;
   2624: result <= 8'b10011101;
   2625: result <= 8'b10011101;
   2626: result <= 8'b10011101;
   2627: result <= 8'b10011101;
   2628: result <= 8'b10011101;
   2629: result <= 8'b10011100;
   2630: result <= 8'b10011100;
   2631: result <= 8'b10011100;
   2632: result <= 8'b10011100;
   2633: result <= 8'b10011100;
   2634: result <= 8'b10011100;
   2635: result <= 8'b10011100;
   2636: result <= 8'b10011100;
   2637: result <= 8'b10011011;
   2638: result <= 8'b10011011;
   2639: result <= 8'b10011011;
   2640: result <= 8'b10011011;
   2641: result <= 8'b10011011;
   2642: result <= 8'b10011011;
   2643: result <= 8'b10011011;
   2644: result <= 8'b10011011;
   2645: result <= 8'b10011010;
   2646: result <= 8'b10011010;
   2647: result <= 8'b10011010;
   2648: result <= 8'b10011010;
   2649: result <= 8'b10011010;
   2650: result <= 8'b10011010;
   2651: result <= 8'b10011010;
   2652: result <= 8'b10011010;
   2653: result <= 8'b10011010;
   2654: result <= 8'b10011001;
   2655: result <= 8'b10011001;
   2656: result <= 8'b10011001;
   2657: result <= 8'b10011001;
   2658: result <= 8'b10011001;
   2659: result <= 8'b10011001;
   2660: result <= 8'b10011001;
   2661: result <= 8'b10011001;
   2662: result <= 8'b10011000;
   2663: result <= 8'b10011000;
   2664: result <= 8'b10011000;
   2665: result <= 8'b10011000;
   2666: result <= 8'b10011000;
   2667: result <= 8'b10011000;
   2668: result <= 8'b10011000;
   2669: result <= 8'b10011000;
   2670: result <= 8'b10011000;
   2671: result <= 8'b10010111;
   2672: result <= 8'b10010111;
   2673: result <= 8'b10010111;
   2674: result <= 8'b10010111;
   2675: result <= 8'b10010111;
   2676: result <= 8'b10010111;
   2677: result <= 8'b10010111;
   2678: result <= 8'b10010111;
   2679: result <= 8'b10010111;
   2680: result <= 8'b10010110;
   2681: result <= 8'b10010110;
   2682: result <= 8'b10010110;
   2683: result <= 8'b10010110;
   2684: result <= 8'b10010110;
   2685: result <= 8'b10010110;
   2686: result <= 8'b10010110;
   2687: result <= 8'b10010110;
   2688: result <= 8'b10010110;
   2689: result <= 8'b10010101;
   2690: result <= 8'b10010101;
   2691: result <= 8'b10010101;
   2692: result <= 8'b10010101;
   2693: result <= 8'b10010101;
   2694: result <= 8'b10010101;
   2695: result <= 8'b10010101;
   2696: result <= 8'b10010101;
   2697: result <= 8'b10010101;
   2698: result <= 8'b10010100;
   2699: result <= 8'b10010100;
   2700: result <= 8'b10010100;
   2701: result <= 8'b10010100;
   2702: result <= 8'b10010100;
   2703: result <= 8'b10010100;
   2704: result <= 8'b10010100;
   2705: result <= 8'b10010100;
   2706: result <= 8'b10010100;
   2707: result <= 8'b10010100;
   2708: result <= 8'b10010011;
   2709: result <= 8'b10010011;
   2710: result <= 8'b10010011;
   2711: result <= 8'b10010011;
   2712: result <= 8'b10010011;
   2713: result <= 8'b10010011;
   2714: result <= 8'b10010011;
   2715: result <= 8'b10010011;
   2716: result <= 8'b10010011;
   2717: result <= 8'b10010011;
   2718: result <= 8'b10010010;
   2719: result <= 8'b10010010;
   2720: result <= 8'b10010010;
   2721: result <= 8'b10010010;
   2722: result <= 8'b10010010;
   2723: result <= 8'b10010010;
   2724: result <= 8'b10010010;
   2725: result <= 8'b10010010;
   2726: result <= 8'b10010010;
   2727: result <= 8'b10010010;
   2728: result <= 8'b10010001;
   2729: result <= 8'b10010001;
   2730: result <= 8'b10010001;
   2731: result <= 8'b10010001;
   2732: result <= 8'b10010001;
   2733: result <= 8'b10010001;
   2734: result <= 8'b10010001;
   2735: result <= 8'b10010001;
   2736: result <= 8'b10010001;
   2737: result <= 8'b10010001;
   2738: result <= 8'b10010000;
   2739: result <= 8'b10010000;
   2740: result <= 8'b10010000;
   2741: result <= 8'b10010000;
   2742: result <= 8'b10010000;
   2743: result <= 8'b10010000;
   2744: result <= 8'b10010000;
   2745: result <= 8'b10010000;
   2746: result <= 8'b10010000;
   2747: result <= 8'b10010000;
   2748: result <= 8'b10001111;
   2749: result <= 8'b10001111;
   2750: result <= 8'b10001111;
   2751: result <= 8'b10001111;
   2752: result <= 8'b10001111;
   2753: result <= 8'b10001111;
   2754: result <= 8'b10001111;
   2755: result <= 8'b10001111;
   2756: result <= 8'b10001111;
   2757: result <= 8'b10001111;
   2758: result <= 8'b10001111;
   2759: result <= 8'b10001110;
   2760: result <= 8'b10001110;
   2761: result <= 8'b10001110;
   2762: result <= 8'b10001110;
   2763: result <= 8'b10001110;
   2764: result <= 8'b10001110;
   2765: result <= 8'b10001110;
   2766: result <= 8'b10001110;
   2767: result <= 8'b10001110;
   2768: result <= 8'b10001110;
   2769: result <= 8'b10001110;
   2770: result <= 8'b10001101;
   2771: result <= 8'b10001101;
   2772: result <= 8'b10001101;
   2773: result <= 8'b10001101;
   2774: result <= 8'b10001101;
   2775: result <= 8'b10001101;
   2776: result <= 8'b10001101;
   2777: result <= 8'b10001101;
   2778: result <= 8'b10001101;
   2779: result <= 8'b10001101;
   2780: result <= 8'b10001101;
   2781: result <= 8'b10001101;
   2782: result <= 8'b10001100;
   2783: result <= 8'b10001100;
   2784: result <= 8'b10001100;
   2785: result <= 8'b10001100;
   2786: result <= 8'b10001100;
   2787: result <= 8'b10001100;
   2788: result <= 8'b10001100;
   2789: result <= 8'b10001100;
   2790: result <= 8'b10001100;
   2791: result <= 8'b10001100;
   2792: result <= 8'b10001100;
   2793: result <= 8'b10001100;
   2794: result <= 8'b10001011;
   2795: result <= 8'b10001011;
   2796: result <= 8'b10001011;
   2797: result <= 8'b10001011;
   2798: result <= 8'b10001011;
   2799: result <= 8'b10001011;
   2800: result <= 8'b10001011;
   2801: result <= 8'b10001011;
   2802: result <= 8'b10001011;
   2803: result <= 8'b10001011;
   2804: result <= 8'b10001011;
   2805: result <= 8'b10001011;
   2806: result <= 8'b10001011;
   2807: result <= 8'b10001010;
   2808: result <= 8'b10001010;
   2809: result <= 8'b10001010;
   2810: result <= 8'b10001010;
   2811: result <= 8'b10001010;
   2812: result <= 8'b10001010;
   2813: result <= 8'b10001010;
   2814: result <= 8'b10001010;
   2815: result <= 8'b10001010;
   2816: result <= 8'b10001010;
   2817: result <= 8'b10001010;
   2818: result <= 8'b10001010;
   2819: result <= 8'b10001010;
   2820: result <= 8'b10001001;
   2821: result <= 8'b10001001;
   2822: result <= 8'b10001001;
   2823: result <= 8'b10001001;
   2824: result <= 8'b10001001;
   2825: result <= 8'b10001001;
   2826: result <= 8'b10001001;
   2827: result <= 8'b10001001;
   2828: result <= 8'b10001001;
   2829: result <= 8'b10001001;
   2830: result <= 8'b10001001;
   2831: result <= 8'b10001001;
   2832: result <= 8'b10001001;
   2833: result <= 8'b10001001;
   2834: result <= 8'b10001000;
   2835: result <= 8'b10001000;
   2836: result <= 8'b10001000;
   2837: result <= 8'b10001000;
   2838: result <= 8'b10001000;
   2839: result <= 8'b10001000;
   2840: result <= 8'b10001000;
   2841: result <= 8'b10001000;
   2842: result <= 8'b10001000;
   2843: result <= 8'b10001000;
   2844: result <= 8'b10001000;
   2845: result <= 8'b10001000;
   2846: result <= 8'b10001000;
   2847: result <= 8'b10001000;
   2848: result <= 8'b10000111;
   2849: result <= 8'b10000111;
   2850: result <= 8'b10000111;
   2851: result <= 8'b10000111;
   2852: result <= 8'b10000111;
   2853: result <= 8'b10000111;
   2854: result <= 8'b10000111;
   2855: result <= 8'b10000111;
   2856: result <= 8'b10000111;
   2857: result <= 8'b10000111;
   2858: result <= 8'b10000111;
   2859: result <= 8'b10000111;
   2860: result <= 8'b10000111;
   2861: result <= 8'b10000111;
   2862: result <= 8'b10000111;
   2863: result <= 8'b10000111;
   2864: result <= 8'b10000110;
   2865: result <= 8'b10000110;
   2866: result <= 8'b10000110;
   2867: result <= 8'b10000110;
   2868: result <= 8'b10000110;
   2869: result <= 8'b10000110;
   2870: result <= 8'b10000110;
   2871: result <= 8'b10000110;
   2872: result <= 8'b10000110;
   2873: result <= 8'b10000110;
   2874: result <= 8'b10000110;
   2875: result <= 8'b10000110;
   2876: result <= 8'b10000110;
   2877: result <= 8'b10000110;
   2878: result <= 8'b10000110;
   2879: result <= 8'b10000110;
   2880: result <= 8'b10000110;
   2881: result <= 8'b10000101;
   2882: result <= 8'b10000101;
   2883: result <= 8'b10000101;
   2884: result <= 8'b10000101;
   2885: result <= 8'b10000101;
   2886: result <= 8'b10000101;
   2887: result <= 8'b10000101;
   2888: result <= 8'b10000101;
   2889: result <= 8'b10000101;
   2890: result <= 8'b10000101;
   2891: result <= 8'b10000101;
   2892: result <= 8'b10000101;
   2893: result <= 8'b10000101;
   2894: result <= 8'b10000101;
   2895: result <= 8'b10000101;
   2896: result <= 8'b10000101;
   2897: result <= 8'b10000101;
   2898: result <= 8'b10000101;
   2899: result <= 8'b10000100;
   2900: result <= 8'b10000100;
   2901: result <= 8'b10000100;
   2902: result <= 8'b10000100;
   2903: result <= 8'b10000100;
   2904: result <= 8'b10000100;
   2905: result <= 8'b10000100;
   2906: result <= 8'b10000100;
   2907: result <= 8'b10000100;
   2908: result <= 8'b10000100;
   2909: result <= 8'b10000100;
   2910: result <= 8'b10000100;
   2911: result <= 8'b10000100;
   2912: result <= 8'b10000100;
   2913: result <= 8'b10000100;
   2914: result <= 8'b10000100;
   2915: result <= 8'b10000100;
   2916: result <= 8'b10000100;
   2917: result <= 8'b10000100;
   2918: result <= 8'b10000100;
   2919: result <= 8'b10000100;
   2920: result <= 8'b10000011;
   2921: result <= 8'b10000011;
   2922: result <= 8'b10000011;
   2923: result <= 8'b10000011;
   2924: result <= 8'b10000011;
   2925: result <= 8'b10000011;
   2926: result <= 8'b10000011;
   2927: result <= 8'b10000011;
   2928: result <= 8'b10000011;
   2929: result <= 8'b10000011;
   2930: result <= 8'b10000011;
   2931: result <= 8'b10000011;
   2932: result <= 8'b10000011;
   2933: result <= 8'b10000011;
   2934: result <= 8'b10000011;
   2935: result <= 8'b10000011;
   2936: result <= 8'b10000011;
   2937: result <= 8'b10000011;
   2938: result <= 8'b10000011;
   2939: result <= 8'b10000011;
   2940: result <= 8'b10000011;
   2941: result <= 8'b10000011;
   2942: result <= 8'b10000011;
   2943: result <= 8'b10000010;
   2944: result <= 8'b10000010;
   2945: result <= 8'b10000010;
   2946: result <= 8'b10000010;
   2947: result <= 8'b10000010;
   2948: result <= 8'b10000010;
   2949: result <= 8'b10000010;
   2950: result <= 8'b10000010;
   2951: result <= 8'b10000010;
   2952: result <= 8'b10000010;
   2953: result <= 8'b10000010;
   2954: result <= 8'b10000010;
   2955: result <= 8'b10000010;
   2956: result <= 8'b10000010;
   2957: result <= 8'b10000010;
   2958: result <= 8'b10000010;
   2959: result <= 8'b10000010;
   2960: result <= 8'b10000010;
   2961: result <= 8'b10000010;
   2962: result <= 8'b10000010;
   2963: result <= 8'b10000010;
   2964: result <= 8'b10000010;
   2965: result <= 8'b10000010;
   2966: result <= 8'b10000010;
   2967: result <= 8'b10000010;
   2968: result <= 8'b10000010;
   2969: result <= 8'b10000010;
   2970: result <= 8'b10000010;
   2971: result <= 8'b10000010;
   2972: result <= 8'b10000010;
   2973: result <= 8'b10000001;
   2974: result <= 8'b10000001;
   2975: result <= 8'b10000001;
   2976: result <= 8'b10000001;
   2977: result <= 8'b10000001;
   2978: result <= 8'b10000001;
   2979: result <= 8'b10000001;
   2980: result <= 8'b10000001;
   2981: result <= 8'b10000001;
   2982: result <= 8'b10000001;
   2983: result <= 8'b10000001;
   2984: result <= 8'b10000001;
   2985: result <= 8'b10000001;
   2986: result <= 8'b10000001;
   2987: result <= 8'b10000001;
   2988: result <= 8'b10000001;
   2989: result <= 8'b10000001;
   2990: result <= 8'b10000001;
   2991: result <= 8'b10000001;
   2992: result <= 8'b10000001;
   2993: result <= 8'b10000001;
   2994: result <= 8'b10000001;
   2995: result <= 8'b10000001;
   2996: result <= 8'b10000001;
   2997: result <= 8'b10000001;
   2998: result <= 8'b10000001;
   2999: result <= 8'b10000001;
   3000: result <= 8'b10000001;
   3001: result <= 8'b10000001;
   3002: result <= 8'b10000001;
   3003: result <= 8'b10000001;
   3004: result <= 8'b10000001;
   3005: result <= 8'b10000001;
   3006: result <= 8'b10000001;
   3007: result <= 8'b10000001;
   3008: result <= 8'b10000001;
   3009: result <= 8'b10000001;
   3010: result <= 8'b10000001;
   3011: result <= 8'b10000001;
   3012: result <= 8'b10000001;
   3013: result <= 8'b10000001;
   3014: result <= 8'b10000001;
   3015: result <= 8'b10000000;
   3016: result <= 8'b10000000;
   3017: result <= 8'b10000000;
   3018: result <= 8'b10000000;
   3019: result <= 8'b10000000;
   3020: result <= 8'b10000000;
   3021: result <= 8'b10000000;
   3022: result <= 8'b10000000;
   3023: result <= 8'b10000000;
   3024: result <= 8'b10000000;
   3025: result <= 8'b10000000;
   3026: result <= 8'b10000000;
   3027: result <= 8'b10000000;
   3028: result <= 8'b10000000;
   3029: result <= 8'b10000000;
   3030: result <= 8'b10000000;
   3031: result <= 8'b10000000;
   3032: result <= 8'b10000000;
   3033: result <= 8'b10000000;
   3034: result <= 8'b10000000;
   3035: result <= 8'b10000000;
   3036: result <= 8'b10000000;
   3037: result <= 8'b10000000;
   3038: result <= 8'b10000000;
   3039: result <= 8'b10000000;
   3040: result <= 8'b10000000;
   3041: result <= 8'b10000000;
   3042: result <= 8'b10000000;
   3043: result <= 8'b10000000;
   3044: result <= 8'b10000000;
   3045: result <= 8'b10000000;
   3046: result <= 8'b10000000;
   3047: result <= 8'b10000000;
   3048: result <= 8'b10000000;
   3049: result <= 8'b10000000;
   3050: result <= 8'b10000000;
   3051: result <= 8'b10000000;
   3052: result <= 8'b10000000;
   3053: result <= 8'b10000000;
   3054: result <= 8'b10000000;
   3055: result <= 8'b10000000;
   3056: result <= 8'b10000000;
   3057: result <= 8'b10000000;
   3058: result <= 8'b10000000;
   3059: result <= 8'b10000000;
   3060: result <= 8'b10000000;
   3061: result <= 8'b10000000;
   3062: result <= 8'b10000000;
   3063: result <= 8'b10000000;
   3064: result <= 8'b10000000;
   3065: result <= 8'b10000000;
   3066: result <= 8'b10000000;
   3067: result <= 8'b10000000;
   3068: result <= 8'b10000000;
   3069: result <= 8'b10000000;
   3070: result <= 8'b10000000;
   3071: result <= 8'b10000000;
   3072: result <= 8'b10000000;
   3073: result <= 8'b10000000;
   3074: result <= 8'b10000000;
   3075: result <= 8'b10000000;
   3076: result <= 8'b10000000;
   3077: result <= 8'b10000000;
   3078: result <= 8'b10000000;
   3079: result <= 8'b10000000;
   3080: result <= 8'b10000000;
   3081: result <= 8'b10000000;
   3082: result <= 8'b10000000;
   3083: result <= 8'b10000000;
   3084: result <= 8'b10000000;
   3085: result <= 8'b10000000;
   3086: result <= 8'b10000000;
   3087: result <= 8'b10000000;
   3088: result <= 8'b10000000;
   3089: result <= 8'b10000000;
   3090: result <= 8'b10000000;
   3091: result <= 8'b10000000;
   3092: result <= 8'b10000000;
   3093: result <= 8'b10000000;
   3094: result <= 8'b10000000;
   3095: result <= 8'b10000000;
   3096: result <= 8'b10000000;
   3097: result <= 8'b10000000;
   3098: result <= 8'b10000000;
   3099: result <= 8'b10000000;
   3100: result <= 8'b10000000;
   3101: result <= 8'b10000000;
   3102: result <= 8'b10000000;
   3103: result <= 8'b10000000;
   3104: result <= 8'b10000000;
   3105: result <= 8'b10000000;
   3106: result <= 8'b10000000;
   3107: result <= 8'b10000000;
   3108: result <= 8'b10000000;
   3109: result <= 8'b10000000;
   3110: result <= 8'b10000000;
   3111: result <= 8'b10000000;
   3112: result <= 8'b10000000;
   3113: result <= 8'b10000000;
   3114: result <= 8'b10000000;
   3115: result <= 8'b10000000;
   3116: result <= 8'b10000000;
   3117: result <= 8'b10000000;
   3118: result <= 8'b10000000;
   3119: result <= 8'b10000000;
   3120: result <= 8'b10000000;
   3121: result <= 8'b10000000;
   3122: result <= 8'b10000000;
   3123: result <= 8'b10000000;
   3124: result <= 8'b10000000;
   3125: result <= 8'b10000000;
   3126: result <= 8'b10000000;
   3127: result <= 8'b10000000;
   3128: result <= 8'b10000000;
   3129: result <= 8'b10000000;
   3130: result <= 8'b10000001;
   3131: result <= 8'b10000001;
   3132: result <= 8'b10000001;
   3133: result <= 8'b10000001;
   3134: result <= 8'b10000001;
   3135: result <= 8'b10000001;
   3136: result <= 8'b10000001;
   3137: result <= 8'b10000001;
   3138: result <= 8'b10000001;
   3139: result <= 8'b10000001;
   3140: result <= 8'b10000001;
   3141: result <= 8'b10000001;
   3142: result <= 8'b10000001;
   3143: result <= 8'b10000001;
   3144: result <= 8'b10000001;
   3145: result <= 8'b10000001;
   3146: result <= 8'b10000001;
   3147: result <= 8'b10000001;
   3148: result <= 8'b10000001;
   3149: result <= 8'b10000001;
   3150: result <= 8'b10000001;
   3151: result <= 8'b10000001;
   3152: result <= 8'b10000001;
   3153: result <= 8'b10000001;
   3154: result <= 8'b10000001;
   3155: result <= 8'b10000001;
   3156: result <= 8'b10000001;
   3157: result <= 8'b10000001;
   3158: result <= 8'b10000001;
   3159: result <= 8'b10000001;
   3160: result <= 8'b10000001;
   3161: result <= 8'b10000001;
   3162: result <= 8'b10000001;
   3163: result <= 8'b10000001;
   3164: result <= 8'b10000001;
   3165: result <= 8'b10000001;
   3166: result <= 8'b10000001;
   3167: result <= 8'b10000001;
   3168: result <= 8'b10000001;
   3169: result <= 8'b10000001;
   3170: result <= 8'b10000001;
   3171: result <= 8'b10000001;
   3172: result <= 8'b10000010;
   3173: result <= 8'b10000010;
   3174: result <= 8'b10000010;
   3175: result <= 8'b10000010;
   3176: result <= 8'b10000010;
   3177: result <= 8'b10000010;
   3178: result <= 8'b10000010;
   3179: result <= 8'b10000010;
   3180: result <= 8'b10000010;
   3181: result <= 8'b10000010;
   3182: result <= 8'b10000010;
   3183: result <= 8'b10000010;
   3184: result <= 8'b10000010;
   3185: result <= 8'b10000010;
   3186: result <= 8'b10000010;
   3187: result <= 8'b10000010;
   3188: result <= 8'b10000010;
   3189: result <= 8'b10000010;
   3190: result <= 8'b10000010;
   3191: result <= 8'b10000010;
   3192: result <= 8'b10000010;
   3193: result <= 8'b10000010;
   3194: result <= 8'b10000010;
   3195: result <= 8'b10000010;
   3196: result <= 8'b10000010;
   3197: result <= 8'b10000010;
   3198: result <= 8'b10000010;
   3199: result <= 8'b10000010;
   3200: result <= 8'b10000010;
   3201: result <= 8'b10000010;
   3202: result <= 8'b10000011;
   3203: result <= 8'b10000011;
   3204: result <= 8'b10000011;
   3205: result <= 8'b10000011;
   3206: result <= 8'b10000011;
   3207: result <= 8'b10000011;
   3208: result <= 8'b10000011;
   3209: result <= 8'b10000011;
   3210: result <= 8'b10000011;
   3211: result <= 8'b10000011;
   3212: result <= 8'b10000011;
   3213: result <= 8'b10000011;
   3214: result <= 8'b10000011;
   3215: result <= 8'b10000011;
   3216: result <= 8'b10000011;
   3217: result <= 8'b10000011;
   3218: result <= 8'b10000011;
   3219: result <= 8'b10000011;
   3220: result <= 8'b10000011;
   3221: result <= 8'b10000011;
   3222: result <= 8'b10000011;
   3223: result <= 8'b10000011;
   3224: result <= 8'b10000011;
   3225: result <= 8'b10000100;
   3226: result <= 8'b10000100;
   3227: result <= 8'b10000100;
   3228: result <= 8'b10000100;
   3229: result <= 8'b10000100;
   3230: result <= 8'b10000100;
   3231: result <= 8'b10000100;
   3232: result <= 8'b10000100;
   3233: result <= 8'b10000100;
   3234: result <= 8'b10000100;
   3235: result <= 8'b10000100;
   3236: result <= 8'b10000100;
   3237: result <= 8'b10000100;
   3238: result <= 8'b10000100;
   3239: result <= 8'b10000100;
   3240: result <= 8'b10000100;
   3241: result <= 8'b10000100;
   3242: result <= 8'b10000100;
   3243: result <= 8'b10000100;
   3244: result <= 8'b10000100;
   3245: result <= 8'b10000100;
   3246: result <= 8'b10000101;
   3247: result <= 8'b10000101;
   3248: result <= 8'b10000101;
   3249: result <= 8'b10000101;
   3250: result <= 8'b10000101;
   3251: result <= 8'b10000101;
   3252: result <= 8'b10000101;
   3253: result <= 8'b10000101;
   3254: result <= 8'b10000101;
   3255: result <= 8'b10000101;
   3256: result <= 8'b10000101;
   3257: result <= 8'b10000101;
   3258: result <= 8'b10000101;
   3259: result <= 8'b10000101;
   3260: result <= 8'b10000101;
   3261: result <= 8'b10000101;
   3262: result <= 8'b10000101;
   3263: result <= 8'b10000101;
   3264: result <= 8'b10000110;
   3265: result <= 8'b10000110;
   3266: result <= 8'b10000110;
   3267: result <= 8'b10000110;
   3268: result <= 8'b10000110;
   3269: result <= 8'b10000110;
   3270: result <= 8'b10000110;
   3271: result <= 8'b10000110;
   3272: result <= 8'b10000110;
   3273: result <= 8'b10000110;
   3274: result <= 8'b10000110;
   3275: result <= 8'b10000110;
   3276: result <= 8'b10000110;
   3277: result <= 8'b10000110;
   3278: result <= 8'b10000110;
   3279: result <= 8'b10000110;
   3280: result <= 8'b10000110;
   3281: result <= 8'b10000111;
   3282: result <= 8'b10000111;
   3283: result <= 8'b10000111;
   3284: result <= 8'b10000111;
   3285: result <= 8'b10000111;
   3286: result <= 8'b10000111;
   3287: result <= 8'b10000111;
   3288: result <= 8'b10000111;
   3289: result <= 8'b10000111;
   3290: result <= 8'b10000111;
   3291: result <= 8'b10000111;
   3292: result <= 8'b10000111;
   3293: result <= 8'b10000111;
   3294: result <= 8'b10000111;
   3295: result <= 8'b10000111;
   3296: result <= 8'b10000111;
   3297: result <= 8'b10001000;
   3298: result <= 8'b10001000;
   3299: result <= 8'b10001000;
   3300: result <= 8'b10001000;
   3301: result <= 8'b10001000;
   3302: result <= 8'b10001000;
   3303: result <= 8'b10001000;
   3304: result <= 8'b10001000;
   3305: result <= 8'b10001000;
   3306: result <= 8'b10001000;
   3307: result <= 8'b10001000;
   3308: result <= 8'b10001000;
   3309: result <= 8'b10001000;
   3310: result <= 8'b10001000;
   3311: result <= 8'b10001001;
   3312: result <= 8'b10001001;
   3313: result <= 8'b10001001;
   3314: result <= 8'b10001001;
   3315: result <= 8'b10001001;
   3316: result <= 8'b10001001;
   3317: result <= 8'b10001001;
   3318: result <= 8'b10001001;
   3319: result <= 8'b10001001;
   3320: result <= 8'b10001001;
   3321: result <= 8'b10001001;
   3322: result <= 8'b10001001;
   3323: result <= 8'b10001001;
   3324: result <= 8'b10001001;
   3325: result <= 8'b10001010;
   3326: result <= 8'b10001010;
   3327: result <= 8'b10001010;
   3328: result <= 8'b10001010;
   3329: result <= 8'b10001010;
   3330: result <= 8'b10001010;
   3331: result <= 8'b10001010;
   3332: result <= 8'b10001010;
   3333: result <= 8'b10001010;
   3334: result <= 8'b10001010;
   3335: result <= 8'b10001010;
   3336: result <= 8'b10001010;
   3337: result <= 8'b10001010;
   3338: result <= 8'b10001011;
   3339: result <= 8'b10001011;
   3340: result <= 8'b10001011;
   3341: result <= 8'b10001011;
   3342: result <= 8'b10001011;
   3343: result <= 8'b10001011;
   3344: result <= 8'b10001011;
   3345: result <= 8'b10001011;
   3346: result <= 8'b10001011;
   3347: result <= 8'b10001011;
   3348: result <= 8'b10001011;
   3349: result <= 8'b10001011;
   3350: result <= 8'b10001011;
   3351: result <= 8'b10001100;
   3352: result <= 8'b10001100;
   3353: result <= 8'b10001100;
   3354: result <= 8'b10001100;
   3355: result <= 8'b10001100;
   3356: result <= 8'b10001100;
   3357: result <= 8'b10001100;
   3358: result <= 8'b10001100;
   3359: result <= 8'b10001100;
   3360: result <= 8'b10001100;
   3361: result <= 8'b10001100;
   3362: result <= 8'b10001100;
   3363: result <= 8'b10001101;
   3364: result <= 8'b10001101;
   3365: result <= 8'b10001101;
   3366: result <= 8'b10001101;
   3367: result <= 8'b10001101;
   3368: result <= 8'b10001101;
   3369: result <= 8'b10001101;
   3370: result <= 8'b10001101;
   3371: result <= 8'b10001101;
   3372: result <= 8'b10001101;
   3373: result <= 8'b10001101;
   3374: result <= 8'b10001101;
   3375: result <= 8'b10001110;
   3376: result <= 8'b10001110;
   3377: result <= 8'b10001110;
   3378: result <= 8'b10001110;
   3379: result <= 8'b10001110;
   3380: result <= 8'b10001110;
   3381: result <= 8'b10001110;
   3382: result <= 8'b10001110;
   3383: result <= 8'b10001110;
   3384: result <= 8'b10001110;
   3385: result <= 8'b10001110;
   3386: result <= 8'b10001111;
   3387: result <= 8'b10001111;
   3388: result <= 8'b10001111;
   3389: result <= 8'b10001111;
   3390: result <= 8'b10001111;
   3391: result <= 8'b10001111;
   3392: result <= 8'b10001111;
   3393: result <= 8'b10001111;
   3394: result <= 8'b10001111;
   3395: result <= 8'b10001111;
   3396: result <= 8'b10001111;
   3397: result <= 8'b10010000;
   3398: result <= 8'b10010000;
   3399: result <= 8'b10010000;
   3400: result <= 8'b10010000;
   3401: result <= 8'b10010000;
   3402: result <= 8'b10010000;
   3403: result <= 8'b10010000;
   3404: result <= 8'b10010000;
   3405: result <= 8'b10010000;
   3406: result <= 8'b10010000;
   3407: result <= 8'b10010001;
   3408: result <= 8'b10010001;
   3409: result <= 8'b10010001;
   3410: result <= 8'b10010001;
   3411: result <= 8'b10010001;
   3412: result <= 8'b10010001;
   3413: result <= 8'b10010001;
   3414: result <= 8'b10010001;
   3415: result <= 8'b10010001;
   3416: result <= 8'b10010001;
   3417: result <= 8'b10010010;
   3418: result <= 8'b10010010;
   3419: result <= 8'b10010010;
   3420: result <= 8'b10010010;
   3421: result <= 8'b10010010;
   3422: result <= 8'b10010010;
   3423: result <= 8'b10010010;
   3424: result <= 8'b10010010;
   3425: result <= 8'b10010010;
   3426: result <= 8'b10010010;
   3427: result <= 8'b10010011;
   3428: result <= 8'b10010011;
   3429: result <= 8'b10010011;
   3430: result <= 8'b10010011;
   3431: result <= 8'b10010011;
   3432: result <= 8'b10010011;
   3433: result <= 8'b10010011;
   3434: result <= 8'b10010011;
   3435: result <= 8'b10010011;
   3436: result <= 8'b10010011;
   3437: result <= 8'b10010100;
   3438: result <= 8'b10010100;
   3439: result <= 8'b10010100;
   3440: result <= 8'b10010100;
   3441: result <= 8'b10010100;
   3442: result <= 8'b10010100;
   3443: result <= 8'b10010100;
   3444: result <= 8'b10010100;
   3445: result <= 8'b10010100;
   3446: result <= 8'b10010100;
   3447: result <= 8'b10010101;
   3448: result <= 8'b10010101;
   3449: result <= 8'b10010101;
   3450: result <= 8'b10010101;
   3451: result <= 8'b10010101;
   3452: result <= 8'b10010101;
   3453: result <= 8'b10010101;
   3454: result <= 8'b10010101;
   3455: result <= 8'b10010101;
   3456: result <= 8'b10010110;
   3457: result <= 8'b10010110;
   3458: result <= 8'b10010110;
   3459: result <= 8'b10010110;
   3460: result <= 8'b10010110;
   3461: result <= 8'b10010110;
   3462: result <= 8'b10010110;
   3463: result <= 8'b10010110;
   3464: result <= 8'b10010110;
   3465: result <= 8'b10010111;
   3466: result <= 8'b10010111;
   3467: result <= 8'b10010111;
   3468: result <= 8'b10010111;
   3469: result <= 8'b10010111;
   3470: result <= 8'b10010111;
   3471: result <= 8'b10010111;
   3472: result <= 8'b10010111;
   3473: result <= 8'b10010111;
   3474: result <= 8'b10011000;
   3475: result <= 8'b10011000;
   3476: result <= 8'b10011000;
   3477: result <= 8'b10011000;
   3478: result <= 8'b10011000;
   3479: result <= 8'b10011000;
   3480: result <= 8'b10011000;
   3481: result <= 8'b10011000;
   3482: result <= 8'b10011000;
   3483: result <= 8'b10011001;
   3484: result <= 8'b10011001;
   3485: result <= 8'b10011001;
   3486: result <= 8'b10011001;
   3487: result <= 8'b10011001;
   3488: result <= 8'b10011001;
   3489: result <= 8'b10011001;
   3490: result <= 8'b10011001;
   3491: result <= 8'b10011010;
   3492: result <= 8'b10011010;
   3493: result <= 8'b10011010;
   3494: result <= 8'b10011010;
   3495: result <= 8'b10011010;
   3496: result <= 8'b10011010;
   3497: result <= 8'b10011010;
   3498: result <= 8'b10011010;
   3499: result <= 8'b10011010;
   3500: result <= 8'b10011011;
   3501: result <= 8'b10011011;
   3502: result <= 8'b10011011;
   3503: result <= 8'b10011011;
   3504: result <= 8'b10011011;
   3505: result <= 8'b10011011;
   3506: result <= 8'b10011011;
   3507: result <= 8'b10011011;
   3508: result <= 8'b10011100;
   3509: result <= 8'b10011100;
   3510: result <= 8'b10011100;
   3511: result <= 8'b10011100;
   3512: result <= 8'b10011100;
   3513: result <= 8'b10011100;
   3514: result <= 8'b10011100;
   3515: result <= 8'b10011100;
   3516: result <= 8'b10011101;
   3517: result <= 8'b10011101;
   3518: result <= 8'b10011101;
   3519: result <= 8'b10011101;
   3520: result <= 8'b10011101;
   3521: result <= 8'b10011101;
   3522: result <= 8'b10011101;
   3523: result <= 8'b10011101;
   3524: result <= 8'b10011110;
   3525: result <= 8'b10011110;
   3526: result <= 8'b10011110;
   3527: result <= 8'b10011110;
   3528: result <= 8'b10011110;
   3529: result <= 8'b10011110;
   3530: result <= 8'b10011110;
   3531: result <= 8'b10011110;
   3532: result <= 8'b10011111;
   3533: result <= 8'b10011111;
   3534: result <= 8'b10011111;
   3535: result <= 8'b10011111;
   3536: result <= 8'b10011111;
   3537: result <= 8'b10011111;
   3538: result <= 8'b10011111;
   3539: result <= 8'b10011111;
   3540: result <= 8'b10100000;
   3541: result <= 8'b10100000;
   3542: result <= 8'b10100000;
   3543: result <= 8'b10100000;
   3544: result <= 8'b10100000;
   3545: result <= 8'b10100000;
   3546: result <= 8'b10100000;
   3547: result <= 8'b10100001;
   3548: result <= 8'b10100001;
   3549: result <= 8'b10100001;
   3550: result <= 8'b10100001;
   3551: result <= 8'b10100001;
   3552: result <= 8'b10100001;
   3553: result <= 8'b10100001;
   3554: result <= 8'b10100001;
   3555: result <= 8'b10100010;
   3556: result <= 8'b10100010;
   3557: result <= 8'b10100010;
   3558: result <= 8'b10100010;
   3559: result <= 8'b10100010;
   3560: result <= 8'b10100010;
   3561: result <= 8'b10100010;
   3562: result <= 8'b10100010;
   3563: result <= 8'b10100011;
   3564: result <= 8'b10100011;
   3565: result <= 8'b10100011;
   3566: result <= 8'b10100011;
   3567: result <= 8'b10100011;
   3568: result <= 8'b10100011;
   3569: result <= 8'b10100011;
   3570: result <= 8'b10100100;
   3571: result <= 8'b10100100;
   3572: result <= 8'b10100100;
   3573: result <= 8'b10100100;
   3574: result <= 8'b10100100;
   3575: result <= 8'b10100100;
   3576: result <= 8'b10100100;
   3577: result <= 8'b10100101;
   3578: result <= 8'b10100101;
   3579: result <= 8'b10100101;
   3580: result <= 8'b10100101;
   3581: result <= 8'b10100101;
   3582: result <= 8'b10100101;
   3583: result <= 8'b10100101;
   3584: result <= 8'b10100101;
   3585: result <= 8'b10100110;
   3586: result <= 8'b10100110;
   3587: result <= 8'b10100110;
   3588: result <= 8'b10100110;
   3589: result <= 8'b10100110;
   3590: result <= 8'b10100110;
   3591: result <= 8'b10100110;
   3592: result <= 8'b10100111;
   3593: result <= 8'b10100111;
   3594: result <= 8'b10100111;
   3595: result <= 8'b10100111;
   3596: result <= 8'b10100111;
   3597: result <= 8'b10100111;
   3598: result <= 8'b10100111;
   3599: result <= 8'b10101000;
   3600: result <= 8'b10101000;
   3601: result <= 8'b10101000;
   3602: result <= 8'b10101000;
   3603: result <= 8'b10101000;
   3604: result <= 8'b10101000;
   3605: result <= 8'b10101000;
   3606: result <= 8'b10101001;
   3607: result <= 8'b10101001;
   3608: result <= 8'b10101001;
   3609: result <= 8'b10101001;
   3610: result <= 8'b10101001;
   3611: result <= 8'b10101001;
   3612: result <= 8'b10101001;
   3613: result <= 8'b10101010;
   3614: result <= 8'b10101010;
   3615: result <= 8'b10101010;
   3616: result <= 8'b10101010;
   3617: result <= 8'b10101010;
   3618: result <= 8'b10101010;
   3619: result <= 8'b10101010;
   3620: result <= 8'b10101011;
   3621: result <= 8'b10101011;
   3622: result <= 8'b10101011;
   3623: result <= 8'b10101011;
   3624: result <= 8'b10101011;
   3625: result <= 8'b10101011;
   3626: result <= 8'b10101100;
   3627: result <= 8'b10101100;
   3628: result <= 8'b10101100;
   3629: result <= 8'b10101100;
   3630: result <= 8'b10101100;
   3631: result <= 8'b10101100;
   3632: result <= 8'b10101100;
   3633: result <= 8'b10101101;
   3634: result <= 8'b10101101;
   3635: result <= 8'b10101101;
   3636: result <= 8'b10101101;
   3637: result <= 8'b10101101;
   3638: result <= 8'b10101101;
   3639: result <= 8'b10101101;
   3640: result <= 8'b10101110;
   3641: result <= 8'b10101110;
   3642: result <= 8'b10101110;
   3643: result <= 8'b10101110;
   3644: result <= 8'b10101110;
   3645: result <= 8'b10101110;
   3646: result <= 8'b10101110;
   3647: result <= 8'b10101111;
   3648: result <= 8'b10101111;
   3649: result <= 8'b10101111;
   3650: result <= 8'b10101111;
   3651: result <= 8'b10101111;
   3652: result <= 8'b10101111;
   3653: result <= 8'b10110000;
   3654: result <= 8'b10110000;
   3655: result <= 8'b10110000;
   3656: result <= 8'b10110000;
   3657: result <= 8'b10110000;
   3658: result <= 8'b10110000;
   3659: result <= 8'b10110000;
   3660: result <= 8'b10110001;
   3661: result <= 8'b10110001;
   3662: result <= 8'b10110001;
   3663: result <= 8'b10110001;
   3664: result <= 8'b10110001;
   3665: result <= 8'b10110001;
   3666: result <= 8'b10110010;
   3667: result <= 8'b10110010;
   3668: result <= 8'b10110010;
   3669: result <= 8'b10110010;
   3670: result <= 8'b10110010;
   3671: result <= 8'b10110010;
   3672: result <= 8'b10110010;
   3673: result <= 8'b10110011;
   3674: result <= 8'b10110011;
   3675: result <= 8'b10110011;
   3676: result <= 8'b10110011;
   3677: result <= 8'b10110011;
   3678: result <= 8'b10110011;
   3679: result <= 8'b10110100;
   3680: result <= 8'b10110100;
   3681: result <= 8'b10110100;
   3682: result <= 8'b10110100;
   3683: result <= 8'b10110100;
   3684: result <= 8'b10110100;
   3685: result <= 8'b10110101;
   3686: result <= 8'b10110101;
   3687: result <= 8'b10110101;
   3688: result <= 8'b10110101;
   3689: result <= 8'b10110101;
   3690: result <= 8'b10110101;
   3691: result <= 8'b10110101;
   3692: result <= 8'b10110110;
   3693: result <= 8'b10110110;
   3694: result <= 8'b10110110;
   3695: result <= 8'b10110110;
   3696: result <= 8'b10110110;
   3697: result <= 8'b10110110;
   3698: result <= 8'b10110111;
   3699: result <= 8'b10110111;
   3700: result <= 8'b10110111;
   3701: result <= 8'b10110111;
   3702: result <= 8'b10110111;
   3703: result <= 8'b10110111;
   3704: result <= 8'b10111000;
   3705: result <= 8'b10111000;
   3706: result <= 8'b10111000;
   3707: result <= 8'b10111000;
   3708: result <= 8'b10111000;
   3709: result <= 8'b10111000;
   3710: result <= 8'b10111001;
   3711: result <= 8'b10111001;
   3712: result <= 8'b10111001;
   3713: result <= 8'b10111001;
   3714: result <= 8'b10111001;
   3715: result <= 8'b10111001;
   3716: result <= 8'b10111010;
   3717: result <= 8'b10111010;
   3718: result <= 8'b10111010;
   3719: result <= 8'b10111010;
   3720: result <= 8'b10111010;
   3721: result <= 8'b10111010;
   3722: result <= 8'b10111011;
   3723: result <= 8'b10111011;
   3724: result <= 8'b10111011;
   3725: result <= 8'b10111011;
   3726: result <= 8'b10111011;
   3727: result <= 8'b10111011;
   3728: result <= 8'b10111100;
   3729: result <= 8'b10111100;
   3730: result <= 8'b10111100;
   3731: result <= 8'b10111100;
   3732: result <= 8'b10111100;
   3733: result <= 8'b10111100;
   3734: result <= 8'b10111101;
   3735: result <= 8'b10111101;
   3736: result <= 8'b10111101;
   3737: result <= 8'b10111101;
   3738: result <= 8'b10111101;
   3739: result <= 8'b10111101;
   3740: result <= 8'b10111110;
   3741: result <= 8'b10111110;
   3742: result <= 8'b10111110;
   3743: result <= 8'b10111110;
   3744: result <= 8'b10111110;
   3745: result <= 8'b10111110;
   3746: result <= 8'b10111111;
   3747: result <= 8'b10111111;
   3748: result <= 8'b10111111;
   3749: result <= 8'b10111111;
   3750: result <= 8'b10111111;
   3751: result <= 8'b10111111;
   3752: result <= 8'b11000000;
   3753: result <= 8'b11000000;
   3754: result <= 8'b11000000;
   3755: result <= 8'b11000000;
   3756: result <= 8'b11000000;
   3757: result <= 8'b11000000;
   3758: result <= 8'b11000001;
   3759: result <= 8'b11000001;
   3760: result <= 8'b11000001;
   3761: result <= 8'b11000001;
   3762: result <= 8'b11000001;
   3763: result <= 8'b11000001;
   3764: result <= 8'b11000010;
   3765: result <= 8'b11000010;
   3766: result <= 8'b11000010;
   3767: result <= 8'b11000010;
   3768: result <= 8'b11000010;
   3769: result <= 8'b11000010;
   3770: result <= 8'b11000011;
   3771: result <= 8'b11000011;
   3772: result <= 8'b11000011;
   3773: result <= 8'b11000011;
   3774: result <= 8'b11000011;
   3775: result <= 8'b11000011;
   3776: result <= 8'b11000100;
   3777: result <= 8'b11000100;
   3778: result <= 8'b11000100;
   3779: result <= 8'b11000100;
   3780: result <= 8'b11000100;
   3781: result <= 8'b11000101;
   3782: result <= 8'b11000101;
   3783: result <= 8'b11000101;
   3784: result <= 8'b11000101;
   3785: result <= 8'b11000101;
   3786: result <= 8'b11000101;
   3787: result <= 8'b11000110;
   3788: result <= 8'b11000110;
   3789: result <= 8'b11000110;
   3790: result <= 8'b11000110;
   3791: result <= 8'b11000110;
   3792: result <= 8'b11000110;
   3793: result <= 8'b11000111;
   3794: result <= 8'b11000111;
   3795: result <= 8'b11000111;
   3796: result <= 8'b11000111;
   3797: result <= 8'b11000111;
   3798: result <= 8'b11001000;
   3799: result <= 8'b11001000;
   3800: result <= 8'b11001000;
   3801: result <= 8'b11001000;
   3802: result <= 8'b11001000;
   3803: result <= 8'b11001000;
   3804: result <= 8'b11001001;
   3805: result <= 8'b11001001;
   3806: result <= 8'b11001001;
   3807: result <= 8'b11001001;
   3808: result <= 8'b11001001;
   3809: result <= 8'b11001001;
   3810: result <= 8'b11001010;
   3811: result <= 8'b11001010;
   3812: result <= 8'b11001010;
   3813: result <= 8'b11001010;
   3814: result <= 8'b11001010;
   3815: result <= 8'b11001011;
   3816: result <= 8'b11001011;
   3817: result <= 8'b11001011;
   3818: result <= 8'b11001011;
   3819: result <= 8'b11001011;
   3820: result <= 8'b11001011;
   3821: result <= 8'b11001100;
   3822: result <= 8'b11001100;
   3823: result <= 8'b11001100;
   3824: result <= 8'b11001100;
   3825: result <= 8'b11001100;
   3826: result <= 8'b11001100;
   3827: result <= 8'b11001101;
   3828: result <= 8'b11001101;
   3829: result <= 8'b11001101;
   3830: result <= 8'b11001101;
   3831: result <= 8'b11001101;
   3832: result <= 8'b11001110;
   3833: result <= 8'b11001110;
   3834: result <= 8'b11001110;
   3835: result <= 8'b11001110;
   3836: result <= 8'b11001110;
   3837: result <= 8'b11001110;
   3838: result <= 8'b11001111;
   3839: result <= 8'b11001111;
   3840: result <= 8'b11001111;
   3841: result <= 8'b11001111;
   3842: result <= 8'b11001111;
   3843: result <= 8'b11010000;
   3844: result <= 8'b11010000;
   3845: result <= 8'b11010000;
   3846: result <= 8'b11010000;
   3847: result <= 8'b11010000;
   3848: result <= 8'b11010000;
   3849: result <= 8'b11010001;
   3850: result <= 8'b11010001;
   3851: result <= 8'b11010001;
   3852: result <= 8'b11010001;
   3853: result <= 8'b11010001;
   3854: result <= 8'b11010010;
   3855: result <= 8'b11010010;
   3856: result <= 8'b11010010;
   3857: result <= 8'b11010010;
   3858: result <= 8'b11010010;
   3859: result <= 8'b11010010;
   3860: result <= 8'b11010011;
   3861: result <= 8'b11010011;
   3862: result <= 8'b11010011;
   3863: result <= 8'b11010011;
   3864: result <= 8'b11010011;
   3865: result <= 8'b11010100;
   3866: result <= 8'b11010100;
   3867: result <= 8'b11010100;
   3868: result <= 8'b11010100;
   3869: result <= 8'b11010100;
   3870: result <= 8'b11010101;
   3871: result <= 8'b11010101;
   3872: result <= 8'b11010101;
   3873: result <= 8'b11010101;
   3874: result <= 8'b11010101;
   3875: result <= 8'b11010101;
   3876: result <= 8'b11010110;
   3877: result <= 8'b11010110;
   3878: result <= 8'b11010110;
   3879: result <= 8'b11010110;
   3880: result <= 8'b11010110;
   3881: result <= 8'b11010111;
   3882: result <= 8'b11010111;
   3883: result <= 8'b11010111;
   3884: result <= 8'b11010111;
   3885: result <= 8'b11010111;
   3886: result <= 8'b11010111;
   3887: result <= 8'b11011000;
   3888: result <= 8'b11011000;
   3889: result <= 8'b11011000;
   3890: result <= 8'b11011000;
   3891: result <= 8'b11011000;
   3892: result <= 8'b11011001;
   3893: result <= 8'b11011001;
   3894: result <= 8'b11011001;
   3895: result <= 8'b11011001;
   3896: result <= 8'b11011001;
   3897: result <= 8'b11011010;
   3898: result <= 8'b11011010;
   3899: result <= 8'b11011010;
   3900: result <= 8'b11011010;
   3901: result <= 8'b11011010;
   3902: result <= 8'b11011010;
   3903: result <= 8'b11011011;
   3904: result <= 8'b11011011;
   3905: result <= 8'b11011011;
   3906: result <= 8'b11011011;
   3907: result <= 8'b11011011;
   3908: result <= 8'b11011100;
   3909: result <= 8'b11011100;
   3910: result <= 8'b11011100;
   3911: result <= 8'b11011100;
   3912: result <= 8'b11011100;
   3913: result <= 8'b11011101;
   3914: result <= 8'b11011101;
   3915: result <= 8'b11011101;
   3916: result <= 8'b11011101;
   3917: result <= 8'b11011101;
   3918: result <= 8'b11011101;
   3919: result <= 8'b11011110;
   3920: result <= 8'b11011110;
   3921: result <= 8'b11011110;
   3922: result <= 8'b11011110;
   3923: result <= 8'b11011110;
   3924: result <= 8'b11011111;
   3925: result <= 8'b11011111;
   3926: result <= 8'b11011111;
   3927: result <= 8'b11011111;
   3928: result <= 8'b11011111;
   3929: result <= 8'b11100000;
   3930: result <= 8'b11100000;
   3931: result <= 8'b11100000;
   3932: result <= 8'b11100000;
   3933: result <= 8'b11100000;
   3934: result <= 8'b11100001;
   3935: result <= 8'b11100001;
   3936: result <= 8'b11100001;
   3937: result <= 8'b11100001;
   3938: result <= 8'b11100001;
   3939: result <= 8'b11100001;
   3940: result <= 8'b11100010;
   3941: result <= 8'b11100010;
   3942: result <= 8'b11100010;
   3943: result <= 8'b11100010;
   3944: result <= 8'b11100010;
   3945: result <= 8'b11100011;
   3946: result <= 8'b11100011;
   3947: result <= 8'b11100011;
   3948: result <= 8'b11100011;
   3949: result <= 8'b11100011;
   3950: result <= 8'b11100100;
   3951: result <= 8'b11100100;
   3952: result <= 8'b11100100;
   3953: result <= 8'b11100100;
   3954: result <= 8'b11100100;
   3955: result <= 8'b11100101;
   3956: result <= 8'b11100101;
   3957: result <= 8'b11100101;
   3958: result <= 8'b11100101;
   3959: result <= 8'b11100101;
   3960: result <= 8'b11100101;
   3961: result <= 8'b11100110;
   3962: result <= 8'b11100110;
   3963: result <= 8'b11100110;
   3964: result <= 8'b11100110;
   3965: result <= 8'b11100110;
   3966: result <= 8'b11100111;
   3967: result <= 8'b11100111;
   3968: result <= 8'b11100111;
   3969: result <= 8'b11100111;
   3970: result <= 8'b11100111;
   3971: result <= 8'b11101000;
   3972: result <= 8'b11101000;
   3973: result <= 8'b11101000;
   3974: result <= 8'b11101000;
   3975: result <= 8'b11101000;
   3976: result <= 8'b11101001;
   3977: result <= 8'b11101001;
   3978: result <= 8'b11101001;
   3979: result <= 8'b11101001;
   3980: result <= 8'b11101001;
   3981: result <= 8'b11101010;
   3982: result <= 8'b11101010;
   3983: result <= 8'b11101010;
   3984: result <= 8'b11101010;
   3985: result <= 8'b11101010;
   3986: result <= 8'b11101011;
   3987: result <= 8'b11101011;
   3988: result <= 8'b11101011;
   3989: result <= 8'b11101011;
   3990: result <= 8'b11101011;
   3991: result <= 8'b11101011;
   3992: result <= 8'b11101100;
   3993: result <= 8'b11101100;
   3994: result <= 8'b11101100;
   3995: result <= 8'b11101100;
   3996: result <= 8'b11101100;
   3997: result <= 8'b11101101;
   3998: result <= 8'b11101101;
   3999: result <= 8'b11101101;
   4000: result <= 8'b11101101;
   4001: result <= 8'b11101101;
   4002: result <= 8'b11101110;
   4003: result <= 8'b11101110;
   4004: result <= 8'b11101110;
   4005: result <= 8'b11101110;
   4006: result <= 8'b11101110;
   4007: result <= 8'b11101111;
   4008: result <= 8'b11101111;
   4009: result <= 8'b11101111;
   4010: result <= 8'b11101111;
   4011: result <= 8'b11101111;
   4012: result <= 8'b11110000;
   4013: result <= 8'b11110000;
   4014: result <= 8'b11110000;
   4015: result <= 8'b11110000;
   4016: result <= 8'b11110000;
   4017: result <= 8'b11110001;
   4018: result <= 8'b11110001;
   4019: result <= 8'b11110001;
   4020: result <= 8'b11110001;
   4021: result <= 8'b11110001;
   4022: result <= 8'b11110010;
   4023: result <= 8'b11110010;
   4024: result <= 8'b11110010;
   4025: result <= 8'b11110010;
   4026: result <= 8'b11110010;
   4027: result <= 8'b11110010;
   4028: result <= 8'b11110011;
   4029: result <= 8'b11110011;
   4030: result <= 8'b11110011;
   4031: result <= 8'b11110011;
   4032: result <= 8'b11110011;
   4033: result <= 8'b11110100;
   4034: result <= 8'b11110100;
   4035: result <= 8'b11110100;
   4036: result <= 8'b11110100;
   4037: result <= 8'b11110100;
   4038: result <= 8'b11110101;
   4039: result <= 8'b11110101;
   4040: result <= 8'b11110101;
   4041: result <= 8'b11110101;
   4042: result <= 8'b11110101;
   4043: result <= 8'b11110110;
   4044: result <= 8'b11110110;
   4045: result <= 8'b11110110;
   4046: result <= 8'b11110110;
   4047: result <= 8'b11110110;
   4048: result <= 8'b11110111;
   4049: result <= 8'b11110111;
   4050: result <= 8'b11110111;
   4051: result <= 8'b11110111;
   4052: result <= 8'b11110111;
   4053: result <= 8'b11111000;
   4054: result <= 8'b11111000;
   4055: result <= 8'b11111000;
   4056: result <= 8'b11111000;
   4057: result <= 8'b11111000;
   4058: result <= 8'b11111001;
   4059: result <= 8'b11111001;
   4060: result <= 8'b11111001;
   4061: result <= 8'b11111001;
   4062: result <= 8'b11111001;
   4063: result <= 8'b11111010;
   4064: result <= 8'b11111010;
   4065: result <= 8'b11111010;
   4066: result <= 8'b11111010;
   4067: result <= 8'b11111010;
   4068: result <= 8'b11111011;
   4069: result <= 8'b11111011;
   4070: result <= 8'b11111011;
   4071: result <= 8'b11111011;
   4072: result <= 8'b11111011;
   4073: result <= 8'b11111011;
   4074: result <= 8'b11111100;
   4075: result <= 8'b11111100;
   4076: result <= 8'b11111100;
   4077: result <= 8'b11111100;
   4078: result <= 8'b11111100;
   4079: result <= 8'b11111101;
   4080: result <= 8'b11111101;
   4081: result <= 8'b11111101;
   4082: result <= 8'b11111101;
   4083: result <= 8'b11111101;
   4084: result <= 8'b11111110;
   4085: result <= 8'b11111110;
   4086: result <= 8'b11111110;
   4087: result <= 8'b11111110;
   4088: result <= 8'b11111110;
   4089: result <= 8'b11111111;
   4090: result <= 8'b11111111;
   4091: result <= 8'b11111111;
   4092: result <= 8'b11111111;
   4093: result <= 8'b11111111;
   4094: result <= 8'b00000000;
   4095: result <= 8'b00000000;
   endcase
endmodule
