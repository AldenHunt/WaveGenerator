`timescale 1ns / 1ps
`default_nettype none


//Created by script createsinelookup.py
module sinetable(input wire [15:0] phase, output reg [11:0] result);

always @(*)
  case(phase)
   0: result <= 12'b000000000000;
   1: result <= 12'b000000000000;
   2: result <= 12'b000000000000;
   3: result <= 12'b000000000000;
   4: result <= 12'b000000000000;
   5: result <= 12'b000000000000;
   6: result <= 12'b000000000001;
   7: result <= 12'b000000000001;
   8: result <= 12'b000000000001;
   9: result <= 12'b000000000001;
   10: result <= 12'b000000000001;
   11: result <= 12'b000000000010;
   12: result <= 12'b000000000010;
   13: result <= 12'b000000000010;
   14: result <= 12'b000000000010;
   15: result <= 12'b000000000010;
   16: result <= 12'b000000000011;
   17: result <= 12'b000000000011;
   18: result <= 12'b000000000011;
   19: result <= 12'b000000000011;
   20: result <= 12'b000000000011;
   21: result <= 12'b000000000100;
   22: result <= 12'b000000000100;
   23: result <= 12'b000000000100;
   24: result <= 12'b000000000100;
   25: result <= 12'b000000000100;
   26: result <= 12'b000000000101;
   27: result <= 12'b000000000101;
   28: result <= 12'b000000000101;
   29: result <= 12'b000000000101;
   30: result <= 12'b000000000101;
   31: result <= 12'b000000000110;
   32: result <= 12'b000000000110;
   33: result <= 12'b000000000110;
   34: result <= 12'b000000000110;
   35: result <= 12'b000000000110;
   36: result <= 12'b000000000111;
   37: result <= 12'b000000000111;
   38: result <= 12'b000000000111;
   39: result <= 12'b000000000111;
   40: result <= 12'b000000000111;
   41: result <= 12'b000000001000;
   42: result <= 12'b000000001000;
   43: result <= 12'b000000001000;
   44: result <= 12'b000000001000;
   45: result <= 12'b000000001000;
   46: result <= 12'b000000001001;
   47: result <= 12'b000000001001;
   48: result <= 12'b000000001001;
   49: result <= 12'b000000001001;
   50: result <= 12'b000000001001;
   51: result <= 12'b000000001010;
   52: result <= 12'b000000001010;
   53: result <= 12'b000000001010;
   54: result <= 12'b000000001010;
   55: result <= 12'b000000001010;
   56: result <= 12'b000000001010;
   57: result <= 12'b000000001011;
   58: result <= 12'b000000001011;
   59: result <= 12'b000000001011;
   60: result <= 12'b000000001011;
   61: result <= 12'b000000001011;
   62: result <= 12'b000000001100;
   63: result <= 12'b000000001100;
   64: result <= 12'b000000001100;
   65: result <= 12'b000000001100;
   66: result <= 12'b000000001100;
   67: result <= 12'b000000001101;
   68: result <= 12'b000000001101;
   69: result <= 12'b000000001101;
   70: result <= 12'b000000001101;
   71: result <= 12'b000000001101;
   72: result <= 12'b000000001110;
   73: result <= 12'b000000001110;
   74: result <= 12'b000000001110;
   75: result <= 12'b000000001110;
   76: result <= 12'b000000001110;
   77: result <= 12'b000000001111;
   78: result <= 12'b000000001111;
   79: result <= 12'b000000001111;
   80: result <= 12'b000000001111;
   81: result <= 12'b000000001111;
   82: result <= 12'b000000010000;
   83: result <= 12'b000000010000;
   84: result <= 12'b000000010000;
   85: result <= 12'b000000010000;
   86: result <= 12'b000000010000;
   87: result <= 12'b000000010001;
   88: result <= 12'b000000010001;
   89: result <= 12'b000000010001;
   90: result <= 12'b000000010001;
   91: result <= 12'b000000010001;
   92: result <= 12'b000000010010;
   93: result <= 12'b000000010010;
   94: result <= 12'b000000010010;
   95: result <= 12'b000000010010;
   96: result <= 12'b000000010010;
   97: result <= 12'b000000010011;
   98: result <= 12'b000000010011;
   99: result <= 12'b000000010011;
   100: result <= 12'b000000010011;
   101: result <= 12'b000000010011;
   102: result <= 12'b000000010100;
   103: result <= 12'b000000010100;
   104: result <= 12'b000000010100;
   105: result <= 12'b000000010100;
   106: result <= 12'b000000010100;
   107: result <= 12'b000000010101;
   108: result <= 12'b000000010101;
   109: result <= 12'b000000010101;
   110: result <= 12'b000000010101;
   111: result <= 12'b000000010101;
   112: result <= 12'b000000010101;
   113: result <= 12'b000000010110;
   114: result <= 12'b000000010110;
   115: result <= 12'b000000010110;
   116: result <= 12'b000000010110;
   117: result <= 12'b000000010110;
   118: result <= 12'b000000010111;
   119: result <= 12'b000000010111;
   120: result <= 12'b000000010111;
   121: result <= 12'b000000010111;
   122: result <= 12'b000000010111;
   123: result <= 12'b000000011000;
   124: result <= 12'b000000011000;
   125: result <= 12'b000000011000;
   126: result <= 12'b000000011000;
   127: result <= 12'b000000011000;
   128: result <= 12'b000000011001;
   129: result <= 12'b000000011001;
   130: result <= 12'b000000011001;
   131: result <= 12'b000000011001;
   132: result <= 12'b000000011001;
   133: result <= 12'b000000011010;
   134: result <= 12'b000000011010;
   135: result <= 12'b000000011010;
   136: result <= 12'b000000011010;
   137: result <= 12'b000000011010;
   138: result <= 12'b000000011011;
   139: result <= 12'b000000011011;
   140: result <= 12'b000000011011;
   141: result <= 12'b000000011011;
   142: result <= 12'b000000011011;
   143: result <= 12'b000000011100;
   144: result <= 12'b000000011100;
   145: result <= 12'b000000011100;
   146: result <= 12'b000000011100;
   147: result <= 12'b000000011100;
   148: result <= 12'b000000011101;
   149: result <= 12'b000000011101;
   150: result <= 12'b000000011101;
   151: result <= 12'b000000011101;
   152: result <= 12'b000000011101;
   153: result <= 12'b000000011110;
   154: result <= 12'b000000011110;
   155: result <= 12'b000000011110;
   156: result <= 12'b000000011110;
   157: result <= 12'b000000011110;
   158: result <= 12'b000000011111;
   159: result <= 12'b000000011111;
   160: result <= 12'b000000011111;
   161: result <= 12'b000000011111;
   162: result <= 12'b000000011111;
   163: result <= 12'b000000100000;
   164: result <= 12'b000000100000;
   165: result <= 12'b000000100000;
   166: result <= 12'b000000100000;
   167: result <= 12'b000000100000;
   168: result <= 12'b000000100000;
   169: result <= 12'b000000100001;
   170: result <= 12'b000000100001;
   171: result <= 12'b000000100001;
   172: result <= 12'b000000100001;
   173: result <= 12'b000000100001;
   174: result <= 12'b000000100010;
   175: result <= 12'b000000100010;
   176: result <= 12'b000000100010;
   177: result <= 12'b000000100010;
   178: result <= 12'b000000100010;
   179: result <= 12'b000000100011;
   180: result <= 12'b000000100011;
   181: result <= 12'b000000100011;
   182: result <= 12'b000000100011;
   183: result <= 12'b000000100011;
   184: result <= 12'b000000100100;
   185: result <= 12'b000000100100;
   186: result <= 12'b000000100100;
   187: result <= 12'b000000100100;
   188: result <= 12'b000000100100;
   189: result <= 12'b000000100101;
   190: result <= 12'b000000100101;
   191: result <= 12'b000000100101;
   192: result <= 12'b000000100101;
   193: result <= 12'b000000100101;
   194: result <= 12'b000000100110;
   195: result <= 12'b000000100110;
   196: result <= 12'b000000100110;
   197: result <= 12'b000000100110;
   198: result <= 12'b000000100110;
   199: result <= 12'b000000100111;
   200: result <= 12'b000000100111;
   201: result <= 12'b000000100111;
   202: result <= 12'b000000100111;
   203: result <= 12'b000000100111;
   204: result <= 12'b000000101000;
   205: result <= 12'b000000101000;
   206: result <= 12'b000000101000;
   207: result <= 12'b000000101000;
   208: result <= 12'b000000101000;
   209: result <= 12'b000000101001;
   210: result <= 12'b000000101001;
   211: result <= 12'b000000101001;
   212: result <= 12'b000000101001;
   213: result <= 12'b000000101001;
   214: result <= 12'b000000101010;
   215: result <= 12'b000000101010;
   216: result <= 12'b000000101010;
   217: result <= 12'b000000101010;
   218: result <= 12'b000000101010;
   219: result <= 12'b000000101010;
   220: result <= 12'b000000101011;
   221: result <= 12'b000000101011;
   222: result <= 12'b000000101011;
   223: result <= 12'b000000101011;
   224: result <= 12'b000000101011;
   225: result <= 12'b000000101100;
   226: result <= 12'b000000101100;
   227: result <= 12'b000000101100;
   228: result <= 12'b000000101100;
   229: result <= 12'b000000101100;
   230: result <= 12'b000000101101;
   231: result <= 12'b000000101101;
   232: result <= 12'b000000101101;
   233: result <= 12'b000000101101;
   234: result <= 12'b000000101101;
   235: result <= 12'b000000101110;
   236: result <= 12'b000000101110;
   237: result <= 12'b000000101110;
   238: result <= 12'b000000101110;
   239: result <= 12'b000000101110;
   240: result <= 12'b000000101111;
   241: result <= 12'b000000101111;
   242: result <= 12'b000000101111;
   243: result <= 12'b000000101111;
   244: result <= 12'b000000101111;
   245: result <= 12'b000000110000;
   246: result <= 12'b000000110000;
   247: result <= 12'b000000110000;
   248: result <= 12'b000000110000;
   249: result <= 12'b000000110000;
   250: result <= 12'b000000110001;
   251: result <= 12'b000000110001;
   252: result <= 12'b000000110001;
   253: result <= 12'b000000110001;
   254: result <= 12'b000000110001;
   255: result <= 12'b000000110010;
   256: result <= 12'b000000110010;
   257: result <= 12'b000000110010;
   258: result <= 12'b000000110010;
   259: result <= 12'b000000110010;
   260: result <= 12'b000000110011;
   261: result <= 12'b000000110011;
   262: result <= 12'b000000110011;
   263: result <= 12'b000000110011;
   264: result <= 12'b000000110011;
   265: result <= 12'b000000110100;
   266: result <= 12'b000000110100;
   267: result <= 12'b000000110100;
   268: result <= 12'b000000110100;
   269: result <= 12'b000000110100;
   270: result <= 12'b000000110101;
   271: result <= 12'b000000110101;
   272: result <= 12'b000000110101;
   273: result <= 12'b000000110101;
   274: result <= 12'b000000110101;
   275: result <= 12'b000000110101;
   276: result <= 12'b000000110110;
   277: result <= 12'b000000110110;
   278: result <= 12'b000000110110;
   279: result <= 12'b000000110110;
   280: result <= 12'b000000110110;
   281: result <= 12'b000000110111;
   282: result <= 12'b000000110111;
   283: result <= 12'b000000110111;
   284: result <= 12'b000000110111;
   285: result <= 12'b000000110111;
   286: result <= 12'b000000111000;
   287: result <= 12'b000000111000;
   288: result <= 12'b000000111000;
   289: result <= 12'b000000111000;
   290: result <= 12'b000000111000;
   291: result <= 12'b000000111001;
   292: result <= 12'b000000111001;
   293: result <= 12'b000000111001;
   294: result <= 12'b000000111001;
   295: result <= 12'b000000111001;
   296: result <= 12'b000000111010;
   297: result <= 12'b000000111010;
   298: result <= 12'b000000111010;
   299: result <= 12'b000000111010;
   300: result <= 12'b000000111010;
   301: result <= 12'b000000111011;
   302: result <= 12'b000000111011;
   303: result <= 12'b000000111011;
   304: result <= 12'b000000111011;
   305: result <= 12'b000000111011;
   306: result <= 12'b000000111100;
   307: result <= 12'b000000111100;
   308: result <= 12'b000000111100;
   309: result <= 12'b000000111100;
   310: result <= 12'b000000111100;
   311: result <= 12'b000000111101;
   312: result <= 12'b000000111101;
   313: result <= 12'b000000111101;
   314: result <= 12'b000000111101;
   315: result <= 12'b000000111101;
   316: result <= 12'b000000111110;
   317: result <= 12'b000000111110;
   318: result <= 12'b000000111110;
   319: result <= 12'b000000111110;
   320: result <= 12'b000000111110;
   321: result <= 12'b000000111111;
   322: result <= 12'b000000111111;
   323: result <= 12'b000000111111;
   324: result <= 12'b000000111111;
   325: result <= 12'b000000111111;
   326: result <= 12'b000000111111;
   327: result <= 12'b000001000000;
   328: result <= 12'b000001000000;
   329: result <= 12'b000001000000;
   330: result <= 12'b000001000000;
   331: result <= 12'b000001000000;
   332: result <= 12'b000001000001;
   333: result <= 12'b000001000001;
   334: result <= 12'b000001000001;
   335: result <= 12'b000001000001;
   336: result <= 12'b000001000001;
   337: result <= 12'b000001000010;
   338: result <= 12'b000001000010;
   339: result <= 12'b000001000010;
   340: result <= 12'b000001000010;
   341: result <= 12'b000001000010;
   342: result <= 12'b000001000011;
   343: result <= 12'b000001000011;
   344: result <= 12'b000001000011;
   345: result <= 12'b000001000011;
   346: result <= 12'b000001000011;
   347: result <= 12'b000001000100;
   348: result <= 12'b000001000100;
   349: result <= 12'b000001000100;
   350: result <= 12'b000001000100;
   351: result <= 12'b000001000100;
   352: result <= 12'b000001000101;
   353: result <= 12'b000001000101;
   354: result <= 12'b000001000101;
   355: result <= 12'b000001000101;
   356: result <= 12'b000001000101;
   357: result <= 12'b000001000110;
   358: result <= 12'b000001000110;
   359: result <= 12'b000001000110;
   360: result <= 12'b000001000110;
   361: result <= 12'b000001000110;
   362: result <= 12'b000001000111;
   363: result <= 12'b000001000111;
   364: result <= 12'b000001000111;
   365: result <= 12'b000001000111;
   366: result <= 12'b000001000111;
   367: result <= 12'b000001001000;
   368: result <= 12'b000001001000;
   369: result <= 12'b000001001000;
   370: result <= 12'b000001001000;
   371: result <= 12'b000001001000;
   372: result <= 12'b000001001001;
   373: result <= 12'b000001001001;
   374: result <= 12'b000001001001;
   375: result <= 12'b000001001001;
   376: result <= 12'b000001001001;
   377: result <= 12'b000001001010;
   378: result <= 12'b000001001010;
   379: result <= 12'b000001001010;
   380: result <= 12'b000001001010;
   381: result <= 12'b000001001010;
   382: result <= 12'b000001001010;
   383: result <= 12'b000001001011;
   384: result <= 12'b000001001011;
   385: result <= 12'b000001001011;
   386: result <= 12'b000001001011;
   387: result <= 12'b000001001011;
   388: result <= 12'b000001001100;
   389: result <= 12'b000001001100;
   390: result <= 12'b000001001100;
   391: result <= 12'b000001001100;
   392: result <= 12'b000001001100;
   393: result <= 12'b000001001101;
   394: result <= 12'b000001001101;
   395: result <= 12'b000001001101;
   396: result <= 12'b000001001101;
   397: result <= 12'b000001001101;
   398: result <= 12'b000001001110;
   399: result <= 12'b000001001110;
   400: result <= 12'b000001001110;
   401: result <= 12'b000001001110;
   402: result <= 12'b000001001110;
   403: result <= 12'b000001001111;
   404: result <= 12'b000001001111;
   405: result <= 12'b000001001111;
   406: result <= 12'b000001001111;
   407: result <= 12'b000001001111;
   408: result <= 12'b000001010000;
   409: result <= 12'b000001010000;
   410: result <= 12'b000001010000;
   411: result <= 12'b000001010000;
   412: result <= 12'b000001010000;
   413: result <= 12'b000001010001;
   414: result <= 12'b000001010001;
   415: result <= 12'b000001010001;
   416: result <= 12'b000001010001;
   417: result <= 12'b000001010001;
   418: result <= 12'b000001010010;
   419: result <= 12'b000001010010;
   420: result <= 12'b000001010010;
   421: result <= 12'b000001010010;
   422: result <= 12'b000001010010;
   423: result <= 12'b000001010011;
   424: result <= 12'b000001010011;
   425: result <= 12'b000001010011;
   426: result <= 12'b000001010011;
   427: result <= 12'b000001010011;
   428: result <= 12'b000001010100;
   429: result <= 12'b000001010100;
   430: result <= 12'b000001010100;
   431: result <= 12'b000001010100;
   432: result <= 12'b000001010100;
   433: result <= 12'b000001010100;
   434: result <= 12'b000001010101;
   435: result <= 12'b000001010101;
   436: result <= 12'b000001010101;
   437: result <= 12'b000001010101;
   438: result <= 12'b000001010101;
   439: result <= 12'b000001010110;
   440: result <= 12'b000001010110;
   441: result <= 12'b000001010110;
   442: result <= 12'b000001010110;
   443: result <= 12'b000001010110;
   444: result <= 12'b000001010111;
   445: result <= 12'b000001010111;
   446: result <= 12'b000001010111;
   447: result <= 12'b000001010111;
   448: result <= 12'b000001010111;
   449: result <= 12'b000001011000;
   450: result <= 12'b000001011000;
   451: result <= 12'b000001011000;
   452: result <= 12'b000001011000;
   453: result <= 12'b000001011000;
   454: result <= 12'b000001011001;
   455: result <= 12'b000001011001;
   456: result <= 12'b000001011001;
   457: result <= 12'b000001011001;
   458: result <= 12'b000001011001;
   459: result <= 12'b000001011010;
   460: result <= 12'b000001011010;
   461: result <= 12'b000001011010;
   462: result <= 12'b000001011010;
   463: result <= 12'b000001011010;
   464: result <= 12'b000001011011;
   465: result <= 12'b000001011011;
   466: result <= 12'b000001011011;
   467: result <= 12'b000001011011;
   468: result <= 12'b000001011011;
   469: result <= 12'b000001011100;
   470: result <= 12'b000001011100;
   471: result <= 12'b000001011100;
   472: result <= 12'b000001011100;
   473: result <= 12'b000001011100;
   474: result <= 12'b000001011101;
   475: result <= 12'b000001011101;
   476: result <= 12'b000001011101;
   477: result <= 12'b000001011101;
   478: result <= 12'b000001011101;
   479: result <= 12'b000001011110;
   480: result <= 12'b000001011110;
   481: result <= 12'b000001011110;
   482: result <= 12'b000001011110;
   483: result <= 12'b000001011110;
   484: result <= 12'b000001011110;
   485: result <= 12'b000001011111;
   486: result <= 12'b000001011111;
   487: result <= 12'b000001011111;
   488: result <= 12'b000001011111;
   489: result <= 12'b000001011111;
   490: result <= 12'b000001100000;
   491: result <= 12'b000001100000;
   492: result <= 12'b000001100000;
   493: result <= 12'b000001100000;
   494: result <= 12'b000001100000;
   495: result <= 12'b000001100001;
   496: result <= 12'b000001100001;
   497: result <= 12'b000001100001;
   498: result <= 12'b000001100001;
   499: result <= 12'b000001100001;
   500: result <= 12'b000001100010;
   501: result <= 12'b000001100010;
   502: result <= 12'b000001100010;
   503: result <= 12'b000001100010;
   504: result <= 12'b000001100010;
   505: result <= 12'b000001100011;
   506: result <= 12'b000001100011;
   507: result <= 12'b000001100011;
   508: result <= 12'b000001100011;
   509: result <= 12'b000001100011;
   510: result <= 12'b000001100100;
   511: result <= 12'b000001100100;
   512: result <= 12'b000001100100;
   513: result <= 12'b000001100100;
   514: result <= 12'b000001100100;
   515: result <= 12'b000001100101;
   516: result <= 12'b000001100101;
   517: result <= 12'b000001100101;
   518: result <= 12'b000001100101;
   519: result <= 12'b000001100101;
   520: result <= 12'b000001100110;
   521: result <= 12'b000001100110;
   522: result <= 12'b000001100110;
   523: result <= 12'b000001100110;
   524: result <= 12'b000001100110;
   525: result <= 12'b000001100111;
   526: result <= 12'b000001100111;
   527: result <= 12'b000001100111;
   528: result <= 12'b000001100111;
   529: result <= 12'b000001100111;
   530: result <= 12'b000001101000;
   531: result <= 12'b000001101000;
   532: result <= 12'b000001101000;
   533: result <= 12'b000001101000;
   534: result <= 12'b000001101000;
   535: result <= 12'b000001101001;
   536: result <= 12'b000001101001;
   537: result <= 12'b000001101001;
   538: result <= 12'b000001101001;
   539: result <= 12'b000001101001;
   540: result <= 12'b000001101001;
   541: result <= 12'b000001101010;
   542: result <= 12'b000001101010;
   543: result <= 12'b000001101010;
   544: result <= 12'b000001101010;
   545: result <= 12'b000001101010;
   546: result <= 12'b000001101011;
   547: result <= 12'b000001101011;
   548: result <= 12'b000001101011;
   549: result <= 12'b000001101011;
   550: result <= 12'b000001101011;
   551: result <= 12'b000001101100;
   552: result <= 12'b000001101100;
   553: result <= 12'b000001101100;
   554: result <= 12'b000001101100;
   555: result <= 12'b000001101100;
   556: result <= 12'b000001101101;
   557: result <= 12'b000001101101;
   558: result <= 12'b000001101101;
   559: result <= 12'b000001101101;
   560: result <= 12'b000001101101;
   561: result <= 12'b000001101110;
   562: result <= 12'b000001101110;
   563: result <= 12'b000001101110;
   564: result <= 12'b000001101110;
   565: result <= 12'b000001101110;
   566: result <= 12'b000001101111;
   567: result <= 12'b000001101111;
   568: result <= 12'b000001101111;
   569: result <= 12'b000001101111;
   570: result <= 12'b000001101111;
   571: result <= 12'b000001110000;
   572: result <= 12'b000001110000;
   573: result <= 12'b000001110000;
   574: result <= 12'b000001110000;
   575: result <= 12'b000001110000;
   576: result <= 12'b000001110001;
   577: result <= 12'b000001110001;
   578: result <= 12'b000001110001;
   579: result <= 12'b000001110001;
   580: result <= 12'b000001110001;
   581: result <= 12'b000001110010;
   582: result <= 12'b000001110010;
   583: result <= 12'b000001110010;
   584: result <= 12'b000001110010;
   585: result <= 12'b000001110010;
   586: result <= 12'b000001110011;
   587: result <= 12'b000001110011;
   588: result <= 12'b000001110011;
   589: result <= 12'b000001110011;
   590: result <= 12'b000001110011;
   591: result <= 12'b000001110011;
   592: result <= 12'b000001110100;
   593: result <= 12'b000001110100;
   594: result <= 12'b000001110100;
   595: result <= 12'b000001110100;
   596: result <= 12'b000001110100;
   597: result <= 12'b000001110101;
   598: result <= 12'b000001110101;
   599: result <= 12'b000001110101;
   600: result <= 12'b000001110101;
   601: result <= 12'b000001110101;
   602: result <= 12'b000001110110;
   603: result <= 12'b000001110110;
   604: result <= 12'b000001110110;
   605: result <= 12'b000001110110;
   606: result <= 12'b000001110110;
   607: result <= 12'b000001110111;
   608: result <= 12'b000001110111;
   609: result <= 12'b000001110111;
   610: result <= 12'b000001110111;
   611: result <= 12'b000001110111;
   612: result <= 12'b000001111000;
   613: result <= 12'b000001111000;
   614: result <= 12'b000001111000;
   615: result <= 12'b000001111000;
   616: result <= 12'b000001111000;
   617: result <= 12'b000001111001;
   618: result <= 12'b000001111001;
   619: result <= 12'b000001111001;
   620: result <= 12'b000001111001;
   621: result <= 12'b000001111001;
   622: result <= 12'b000001111010;
   623: result <= 12'b000001111010;
   624: result <= 12'b000001111010;
   625: result <= 12'b000001111010;
   626: result <= 12'b000001111010;
   627: result <= 12'b000001111011;
   628: result <= 12'b000001111011;
   629: result <= 12'b000001111011;
   630: result <= 12'b000001111011;
   631: result <= 12'b000001111011;
   632: result <= 12'b000001111100;
   633: result <= 12'b000001111100;
   634: result <= 12'b000001111100;
   635: result <= 12'b000001111100;
   636: result <= 12'b000001111100;
   637: result <= 12'b000001111100;
   638: result <= 12'b000001111101;
   639: result <= 12'b000001111101;
   640: result <= 12'b000001111101;
   641: result <= 12'b000001111101;
   642: result <= 12'b000001111101;
   643: result <= 12'b000001111110;
   644: result <= 12'b000001111110;
   645: result <= 12'b000001111110;
   646: result <= 12'b000001111110;
   647: result <= 12'b000001111110;
   648: result <= 12'b000001111111;
   649: result <= 12'b000001111111;
   650: result <= 12'b000001111111;
   651: result <= 12'b000001111111;
   652: result <= 12'b000001111111;
   653: result <= 12'b000010000000;
   654: result <= 12'b000010000000;
   655: result <= 12'b000010000000;
   656: result <= 12'b000010000000;
   657: result <= 12'b000010000000;
   658: result <= 12'b000010000001;
   659: result <= 12'b000010000001;
   660: result <= 12'b000010000001;
   661: result <= 12'b000010000001;
   662: result <= 12'b000010000001;
   663: result <= 12'b000010000010;
   664: result <= 12'b000010000010;
   665: result <= 12'b000010000010;
   666: result <= 12'b000010000010;
   667: result <= 12'b000010000010;
   668: result <= 12'b000010000011;
   669: result <= 12'b000010000011;
   670: result <= 12'b000010000011;
   671: result <= 12'b000010000011;
   672: result <= 12'b000010000011;
   673: result <= 12'b000010000100;
   674: result <= 12'b000010000100;
   675: result <= 12'b000010000100;
   676: result <= 12'b000010000100;
   677: result <= 12'b000010000100;
   678: result <= 12'b000010000101;
   679: result <= 12'b000010000101;
   680: result <= 12'b000010000101;
   681: result <= 12'b000010000101;
   682: result <= 12'b000010000101;
   683: result <= 12'b000010000110;
   684: result <= 12'b000010000110;
   685: result <= 12'b000010000110;
   686: result <= 12'b000010000110;
   687: result <= 12'b000010000110;
   688: result <= 12'b000010000110;
   689: result <= 12'b000010000111;
   690: result <= 12'b000010000111;
   691: result <= 12'b000010000111;
   692: result <= 12'b000010000111;
   693: result <= 12'b000010000111;
   694: result <= 12'b000010001000;
   695: result <= 12'b000010001000;
   696: result <= 12'b000010001000;
   697: result <= 12'b000010001000;
   698: result <= 12'b000010001000;
   699: result <= 12'b000010001001;
   700: result <= 12'b000010001001;
   701: result <= 12'b000010001001;
   702: result <= 12'b000010001001;
   703: result <= 12'b000010001001;
   704: result <= 12'b000010001010;
   705: result <= 12'b000010001010;
   706: result <= 12'b000010001010;
   707: result <= 12'b000010001010;
   708: result <= 12'b000010001010;
   709: result <= 12'b000010001011;
   710: result <= 12'b000010001011;
   711: result <= 12'b000010001011;
   712: result <= 12'b000010001011;
   713: result <= 12'b000010001011;
   714: result <= 12'b000010001100;
   715: result <= 12'b000010001100;
   716: result <= 12'b000010001100;
   717: result <= 12'b000010001100;
   718: result <= 12'b000010001100;
   719: result <= 12'b000010001101;
   720: result <= 12'b000010001101;
   721: result <= 12'b000010001101;
   722: result <= 12'b000010001101;
   723: result <= 12'b000010001101;
   724: result <= 12'b000010001110;
   725: result <= 12'b000010001110;
   726: result <= 12'b000010001110;
   727: result <= 12'b000010001110;
   728: result <= 12'b000010001110;
   729: result <= 12'b000010001111;
   730: result <= 12'b000010001111;
   731: result <= 12'b000010001111;
   732: result <= 12'b000010001111;
   733: result <= 12'b000010001111;
   734: result <= 12'b000010010000;
   735: result <= 12'b000010010000;
   736: result <= 12'b000010010000;
   737: result <= 12'b000010010000;
   738: result <= 12'b000010010000;
   739: result <= 12'b000010010000;
   740: result <= 12'b000010010001;
   741: result <= 12'b000010010001;
   742: result <= 12'b000010010001;
   743: result <= 12'b000010010001;
   744: result <= 12'b000010010001;
   745: result <= 12'b000010010010;
   746: result <= 12'b000010010010;
   747: result <= 12'b000010010010;
   748: result <= 12'b000010010010;
   749: result <= 12'b000010010010;
   750: result <= 12'b000010010011;
   751: result <= 12'b000010010011;
   752: result <= 12'b000010010011;
   753: result <= 12'b000010010011;
   754: result <= 12'b000010010011;
   755: result <= 12'b000010010100;
   756: result <= 12'b000010010100;
   757: result <= 12'b000010010100;
   758: result <= 12'b000010010100;
   759: result <= 12'b000010010100;
   760: result <= 12'b000010010101;
   761: result <= 12'b000010010101;
   762: result <= 12'b000010010101;
   763: result <= 12'b000010010101;
   764: result <= 12'b000010010101;
   765: result <= 12'b000010010110;
   766: result <= 12'b000010010110;
   767: result <= 12'b000010010110;
   768: result <= 12'b000010010110;
   769: result <= 12'b000010010110;
   770: result <= 12'b000010010111;
   771: result <= 12'b000010010111;
   772: result <= 12'b000010010111;
   773: result <= 12'b000010010111;
   774: result <= 12'b000010010111;
   775: result <= 12'b000010011000;
   776: result <= 12'b000010011000;
   777: result <= 12'b000010011000;
   778: result <= 12'b000010011000;
   779: result <= 12'b000010011000;
   780: result <= 12'b000010011001;
   781: result <= 12'b000010011001;
   782: result <= 12'b000010011001;
   783: result <= 12'b000010011001;
   784: result <= 12'b000010011001;
   785: result <= 12'b000010011001;
   786: result <= 12'b000010011010;
   787: result <= 12'b000010011010;
   788: result <= 12'b000010011010;
   789: result <= 12'b000010011010;
   790: result <= 12'b000010011010;
   791: result <= 12'b000010011011;
   792: result <= 12'b000010011011;
   793: result <= 12'b000010011011;
   794: result <= 12'b000010011011;
   795: result <= 12'b000010011011;
   796: result <= 12'b000010011100;
   797: result <= 12'b000010011100;
   798: result <= 12'b000010011100;
   799: result <= 12'b000010011100;
   800: result <= 12'b000010011100;
   801: result <= 12'b000010011101;
   802: result <= 12'b000010011101;
   803: result <= 12'b000010011101;
   804: result <= 12'b000010011101;
   805: result <= 12'b000010011101;
   806: result <= 12'b000010011110;
   807: result <= 12'b000010011110;
   808: result <= 12'b000010011110;
   809: result <= 12'b000010011110;
   810: result <= 12'b000010011110;
   811: result <= 12'b000010011111;
   812: result <= 12'b000010011111;
   813: result <= 12'b000010011111;
   814: result <= 12'b000010011111;
   815: result <= 12'b000010011111;
   816: result <= 12'b000010100000;
   817: result <= 12'b000010100000;
   818: result <= 12'b000010100000;
   819: result <= 12'b000010100000;
   820: result <= 12'b000010100000;
   821: result <= 12'b000010100001;
   822: result <= 12'b000010100001;
   823: result <= 12'b000010100001;
   824: result <= 12'b000010100001;
   825: result <= 12'b000010100001;
   826: result <= 12'b000010100010;
   827: result <= 12'b000010100010;
   828: result <= 12'b000010100010;
   829: result <= 12'b000010100010;
   830: result <= 12'b000010100010;
   831: result <= 12'b000010100010;
   832: result <= 12'b000010100011;
   833: result <= 12'b000010100011;
   834: result <= 12'b000010100011;
   835: result <= 12'b000010100011;
   836: result <= 12'b000010100011;
   837: result <= 12'b000010100100;
   838: result <= 12'b000010100100;
   839: result <= 12'b000010100100;
   840: result <= 12'b000010100100;
   841: result <= 12'b000010100100;
   842: result <= 12'b000010100101;
   843: result <= 12'b000010100101;
   844: result <= 12'b000010100101;
   845: result <= 12'b000010100101;
   846: result <= 12'b000010100101;
   847: result <= 12'b000010100110;
   848: result <= 12'b000010100110;
   849: result <= 12'b000010100110;
   850: result <= 12'b000010100110;
   851: result <= 12'b000010100110;
   852: result <= 12'b000010100111;
   853: result <= 12'b000010100111;
   854: result <= 12'b000010100111;
   855: result <= 12'b000010100111;
   856: result <= 12'b000010100111;
   857: result <= 12'b000010101000;
   858: result <= 12'b000010101000;
   859: result <= 12'b000010101000;
   860: result <= 12'b000010101000;
   861: result <= 12'b000010101000;
   862: result <= 12'b000010101001;
   863: result <= 12'b000010101001;
   864: result <= 12'b000010101001;
   865: result <= 12'b000010101001;
   866: result <= 12'b000010101001;
   867: result <= 12'b000010101010;
   868: result <= 12'b000010101010;
   869: result <= 12'b000010101010;
   870: result <= 12'b000010101010;
   871: result <= 12'b000010101010;
   872: result <= 12'b000010101011;
   873: result <= 12'b000010101011;
   874: result <= 12'b000010101011;
   875: result <= 12'b000010101011;
   876: result <= 12'b000010101011;
   877: result <= 12'b000010101011;
   878: result <= 12'b000010101100;
   879: result <= 12'b000010101100;
   880: result <= 12'b000010101100;
   881: result <= 12'b000010101100;
   882: result <= 12'b000010101100;
   883: result <= 12'b000010101101;
   884: result <= 12'b000010101101;
   885: result <= 12'b000010101101;
   886: result <= 12'b000010101101;
   887: result <= 12'b000010101101;
   888: result <= 12'b000010101110;
   889: result <= 12'b000010101110;
   890: result <= 12'b000010101110;
   891: result <= 12'b000010101110;
   892: result <= 12'b000010101110;
   893: result <= 12'b000010101111;
   894: result <= 12'b000010101111;
   895: result <= 12'b000010101111;
   896: result <= 12'b000010101111;
   897: result <= 12'b000010101111;
   898: result <= 12'b000010110000;
   899: result <= 12'b000010110000;
   900: result <= 12'b000010110000;
   901: result <= 12'b000010110000;
   902: result <= 12'b000010110000;
   903: result <= 12'b000010110001;
   904: result <= 12'b000010110001;
   905: result <= 12'b000010110001;
   906: result <= 12'b000010110001;
   907: result <= 12'b000010110001;
   908: result <= 12'b000010110010;
   909: result <= 12'b000010110010;
   910: result <= 12'b000010110010;
   911: result <= 12'b000010110010;
   912: result <= 12'b000010110010;
   913: result <= 12'b000010110011;
   914: result <= 12'b000010110011;
   915: result <= 12'b000010110011;
   916: result <= 12'b000010110011;
   917: result <= 12'b000010110011;
   918: result <= 12'b000010110100;
   919: result <= 12'b000010110100;
   920: result <= 12'b000010110100;
   921: result <= 12'b000010110100;
   922: result <= 12'b000010110100;
   923: result <= 12'b000010110100;
   924: result <= 12'b000010110101;
   925: result <= 12'b000010110101;
   926: result <= 12'b000010110101;
   927: result <= 12'b000010110101;
   928: result <= 12'b000010110101;
   929: result <= 12'b000010110110;
   930: result <= 12'b000010110110;
   931: result <= 12'b000010110110;
   932: result <= 12'b000010110110;
   933: result <= 12'b000010110110;
   934: result <= 12'b000010110111;
   935: result <= 12'b000010110111;
   936: result <= 12'b000010110111;
   937: result <= 12'b000010110111;
   938: result <= 12'b000010110111;
   939: result <= 12'b000010111000;
   940: result <= 12'b000010111000;
   941: result <= 12'b000010111000;
   942: result <= 12'b000010111000;
   943: result <= 12'b000010111000;
   944: result <= 12'b000010111001;
   945: result <= 12'b000010111001;
   946: result <= 12'b000010111001;
   947: result <= 12'b000010111001;
   948: result <= 12'b000010111001;
   949: result <= 12'b000010111010;
   950: result <= 12'b000010111010;
   951: result <= 12'b000010111010;
   952: result <= 12'b000010111010;
   953: result <= 12'b000010111010;
   954: result <= 12'b000010111011;
   955: result <= 12'b000010111011;
   956: result <= 12'b000010111011;
   957: result <= 12'b000010111011;
   958: result <= 12'b000010111011;
   959: result <= 12'b000010111100;
   960: result <= 12'b000010111100;
   961: result <= 12'b000010111100;
   962: result <= 12'b000010111100;
   963: result <= 12'b000010111100;
   964: result <= 12'b000010111101;
   965: result <= 12'b000010111101;
   966: result <= 12'b000010111101;
   967: result <= 12'b000010111101;
   968: result <= 12'b000010111101;
   969: result <= 12'b000010111101;
   970: result <= 12'b000010111110;
   971: result <= 12'b000010111110;
   972: result <= 12'b000010111110;
   973: result <= 12'b000010111110;
   974: result <= 12'b000010111110;
   975: result <= 12'b000010111111;
   976: result <= 12'b000010111111;
   977: result <= 12'b000010111111;
   978: result <= 12'b000010111111;
   979: result <= 12'b000010111111;
   980: result <= 12'b000011000000;
   981: result <= 12'b000011000000;
   982: result <= 12'b000011000000;
   983: result <= 12'b000011000000;
   984: result <= 12'b000011000000;
   985: result <= 12'b000011000001;
   986: result <= 12'b000011000001;
   987: result <= 12'b000011000001;
   988: result <= 12'b000011000001;
   989: result <= 12'b000011000001;
   990: result <= 12'b000011000010;
   991: result <= 12'b000011000010;
   992: result <= 12'b000011000010;
   993: result <= 12'b000011000010;
   994: result <= 12'b000011000010;
   995: result <= 12'b000011000011;
   996: result <= 12'b000011000011;
   997: result <= 12'b000011000011;
   998: result <= 12'b000011000011;
   999: result <= 12'b000011000011;
   1000: result <= 12'b000011000100;
   1001: result <= 12'b000011000100;
   1002: result <= 12'b000011000100;
   1003: result <= 12'b000011000100;
   1004: result <= 12'b000011000100;
   1005: result <= 12'b000011000101;
   1006: result <= 12'b000011000101;
   1007: result <= 12'b000011000101;
   1008: result <= 12'b000011000101;
   1009: result <= 12'b000011000101;
   1010: result <= 12'b000011000110;
   1011: result <= 12'b000011000110;
   1012: result <= 12'b000011000110;
   1013: result <= 12'b000011000110;
   1014: result <= 12'b000011000110;
   1015: result <= 12'b000011000110;
   1016: result <= 12'b000011000111;
   1017: result <= 12'b000011000111;
   1018: result <= 12'b000011000111;
   1019: result <= 12'b000011000111;
   1020: result <= 12'b000011000111;
   1021: result <= 12'b000011001000;
   1022: result <= 12'b000011001000;
   1023: result <= 12'b000011001000;
   1024: result <= 12'b000011001000;
   1025: result <= 12'b000011001000;
   1026: result <= 12'b000011001001;
   1027: result <= 12'b000011001001;
   1028: result <= 12'b000011001001;
   1029: result <= 12'b000011001001;
   1030: result <= 12'b000011001001;
   1031: result <= 12'b000011001010;
   1032: result <= 12'b000011001010;
   1033: result <= 12'b000011001010;
   1034: result <= 12'b000011001010;
   1035: result <= 12'b000011001010;
   1036: result <= 12'b000011001011;
   1037: result <= 12'b000011001011;
   1038: result <= 12'b000011001011;
   1039: result <= 12'b000011001011;
   1040: result <= 12'b000011001011;
   1041: result <= 12'b000011001100;
   1042: result <= 12'b000011001100;
   1043: result <= 12'b000011001100;
   1044: result <= 12'b000011001100;
   1045: result <= 12'b000011001100;
   1046: result <= 12'b000011001101;
   1047: result <= 12'b000011001101;
   1048: result <= 12'b000011001101;
   1049: result <= 12'b000011001101;
   1050: result <= 12'b000011001101;
   1051: result <= 12'b000011001110;
   1052: result <= 12'b000011001110;
   1053: result <= 12'b000011001110;
   1054: result <= 12'b000011001110;
   1055: result <= 12'b000011001110;
   1056: result <= 12'b000011001110;
   1057: result <= 12'b000011001111;
   1058: result <= 12'b000011001111;
   1059: result <= 12'b000011001111;
   1060: result <= 12'b000011001111;
   1061: result <= 12'b000011001111;
   1062: result <= 12'b000011010000;
   1063: result <= 12'b000011010000;
   1064: result <= 12'b000011010000;
   1065: result <= 12'b000011010000;
   1066: result <= 12'b000011010000;
   1067: result <= 12'b000011010001;
   1068: result <= 12'b000011010001;
   1069: result <= 12'b000011010001;
   1070: result <= 12'b000011010001;
   1071: result <= 12'b000011010001;
   1072: result <= 12'b000011010010;
   1073: result <= 12'b000011010010;
   1074: result <= 12'b000011010010;
   1075: result <= 12'b000011010010;
   1076: result <= 12'b000011010010;
   1077: result <= 12'b000011010011;
   1078: result <= 12'b000011010011;
   1079: result <= 12'b000011010011;
   1080: result <= 12'b000011010011;
   1081: result <= 12'b000011010011;
   1082: result <= 12'b000011010100;
   1083: result <= 12'b000011010100;
   1084: result <= 12'b000011010100;
   1085: result <= 12'b000011010100;
   1086: result <= 12'b000011010100;
   1087: result <= 12'b000011010101;
   1088: result <= 12'b000011010101;
   1089: result <= 12'b000011010101;
   1090: result <= 12'b000011010101;
   1091: result <= 12'b000011010101;
   1092: result <= 12'b000011010110;
   1093: result <= 12'b000011010110;
   1094: result <= 12'b000011010110;
   1095: result <= 12'b000011010110;
   1096: result <= 12'b000011010110;
   1097: result <= 12'b000011010110;
   1098: result <= 12'b000011010111;
   1099: result <= 12'b000011010111;
   1100: result <= 12'b000011010111;
   1101: result <= 12'b000011010111;
   1102: result <= 12'b000011010111;
   1103: result <= 12'b000011011000;
   1104: result <= 12'b000011011000;
   1105: result <= 12'b000011011000;
   1106: result <= 12'b000011011000;
   1107: result <= 12'b000011011000;
   1108: result <= 12'b000011011001;
   1109: result <= 12'b000011011001;
   1110: result <= 12'b000011011001;
   1111: result <= 12'b000011011001;
   1112: result <= 12'b000011011001;
   1113: result <= 12'b000011011010;
   1114: result <= 12'b000011011010;
   1115: result <= 12'b000011011010;
   1116: result <= 12'b000011011010;
   1117: result <= 12'b000011011010;
   1118: result <= 12'b000011011011;
   1119: result <= 12'b000011011011;
   1120: result <= 12'b000011011011;
   1121: result <= 12'b000011011011;
   1122: result <= 12'b000011011011;
   1123: result <= 12'b000011011100;
   1124: result <= 12'b000011011100;
   1125: result <= 12'b000011011100;
   1126: result <= 12'b000011011100;
   1127: result <= 12'b000011011100;
   1128: result <= 12'b000011011101;
   1129: result <= 12'b000011011101;
   1130: result <= 12'b000011011101;
   1131: result <= 12'b000011011101;
   1132: result <= 12'b000011011101;
   1133: result <= 12'b000011011110;
   1134: result <= 12'b000011011110;
   1135: result <= 12'b000011011110;
   1136: result <= 12'b000011011110;
   1137: result <= 12'b000011011110;
   1138: result <= 12'b000011011111;
   1139: result <= 12'b000011011111;
   1140: result <= 12'b000011011111;
   1141: result <= 12'b000011011111;
   1142: result <= 12'b000011011111;
   1143: result <= 12'b000011011111;
   1144: result <= 12'b000011100000;
   1145: result <= 12'b000011100000;
   1146: result <= 12'b000011100000;
   1147: result <= 12'b000011100000;
   1148: result <= 12'b000011100000;
   1149: result <= 12'b000011100001;
   1150: result <= 12'b000011100001;
   1151: result <= 12'b000011100001;
   1152: result <= 12'b000011100001;
   1153: result <= 12'b000011100001;
   1154: result <= 12'b000011100010;
   1155: result <= 12'b000011100010;
   1156: result <= 12'b000011100010;
   1157: result <= 12'b000011100010;
   1158: result <= 12'b000011100010;
   1159: result <= 12'b000011100011;
   1160: result <= 12'b000011100011;
   1161: result <= 12'b000011100011;
   1162: result <= 12'b000011100011;
   1163: result <= 12'b000011100011;
   1164: result <= 12'b000011100100;
   1165: result <= 12'b000011100100;
   1166: result <= 12'b000011100100;
   1167: result <= 12'b000011100100;
   1168: result <= 12'b000011100100;
   1169: result <= 12'b000011100101;
   1170: result <= 12'b000011100101;
   1171: result <= 12'b000011100101;
   1172: result <= 12'b000011100101;
   1173: result <= 12'b000011100101;
   1174: result <= 12'b000011100110;
   1175: result <= 12'b000011100110;
   1176: result <= 12'b000011100110;
   1177: result <= 12'b000011100110;
   1178: result <= 12'b000011100110;
   1179: result <= 12'b000011100111;
   1180: result <= 12'b000011100111;
   1181: result <= 12'b000011100111;
   1182: result <= 12'b000011100111;
   1183: result <= 12'b000011100111;
   1184: result <= 12'b000011100111;
   1185: result <= 12'b000011101000;
   1186: result <= 12'b000011101000;
   1187: result <= 12'b000011101000;
   1188: result <= 12'b000011101000;
   1189: result <= 12'b000011101000;
   1190: result <= 12'b000011101001;
   1191: result <= 12'b000011101001;
   1192: result <= 12'b000011101001;
   1193: result <= 12'b000011101001;
   1194: result <= 12'b000011101001;
   1195: result <= 12'b000011101010;
   1196: result <= 12'b000011101010;
   1197: result <= 12'b000011101010;
   1198: result <= 12'b000011101010;
   1199: result <= 12'b000011101010;
   1200: result <= 12'b000011101011;
   1201: result <= 12'b000011101011;
   1202: result <= 12'b000011101011;
   1203: result <= 12'b000011101011;
   1204: result <= 12'b000011101011;
   1205: result <= 12'b000011101100;
   1206: result <= 12'b000011101100;
   1207: result <= 12'b000011101100;
   1208: result <= 12'b000011101100;
   1209: result <= 12'b000011101100;
   1210: result <= 12'b000011101101;
   1211: result <= 12'b000011101101;
   1212: result <= 12'b000011101101;
   1213: result <= 12'b000011101101;
   1214: result <= 12'b000011101101;
   1215: result <= 12'b000011101110;
   1216: result <= 12'b000011101110;
   1217: result <= 12'b000011101110;
   1218: result <= 12'b000011101110;
   1219: result <= 12'b000011101110;
   1220: result <= 12'b000011101111;
   1221: result <= 12'b000011101111;
   1222: result <= 12'b000011101111;
   1223: result <= 12'b000011101111;
   1224: result <= 12'b000011101111;
   1225: result <= 12'b000011101111;
   1226: result <= 12'b000011110000;
   1227: result <= 12'b000011110000;
   1228: result <= 12'b000011110000;
   1229: result <= 12'b000011110000;
   1230: result <= 12'b000011110000;
   1231: result <= 12'b000011110001;
   1232: result <= 12'b000011110001;
   1233: result <= 12'b000011110001;
   1234: result <= 12'b000011110001;
   1235: result <= 12'b000011110001;
   1236: result <= 12'b000011110010;
   1237: result <= 12'b000011110010;
   1238: result <= 12'b000011110010;
   1239: result <= 12'b000011110010;
   1240: result <= 12'b000011110010;
   1241: result <= 12'b000011110011;
   1242: result <= 12'b000011110011;
   1243: result <= 12'b000011110011;
   1244: result <= 12'b000011110011;
   1245: result <= 12'b000011110011;
   1246: result <= 12'b000011110100;
   1247: result <= 12'b000011110100;
   1248: result <= 12'b000011110100;
   1249: result <= 12'b000011110100;
   1250: result <= 12'b000011110100;
   1251: result <= 12'b000011110101;
   1252: result <= 12'b000011110101;
   1253: result <= 12'b000011110101;
   1254: result <= 12'b000011110101;
   1255: result <= 12'b000011110101;
   1256: result <= 12'b000011110110;
   1257: result <= 12'b000011110110;
   1258: result <= 12'b000011110110;
   1259: result <= 12'b000011110110;
   1260: result <= 12'b000011110110;
   1261: result <= 12'b000011110110;
   1262: result <= 12'b000011110111;
   1263: result <= 12'b000011110111;
   1264: result <= 12'b000011110111;
   1265: result <= 12'b000011110111;
   1266: result <= 12'b000011110111;
   1267: result <= 12'b000011111000;
   1268: result <= 12'b000011111000;
   1269: result <= 12'b000011111000;
   1270: result <= 12'b000011111000;
   1271: result <= 12'b000011111000;
   1272: result <= 12'b000011111001;
   1273: result <= 12'b000011111001;
   1274: result <= 12'b000011111001;
   1275: result <= 12'b000011111001;
   1276: result <= 12'b000011111001;
   1277: result <= 12'b000011111010;
   1278: result <= 12'b000011111010;
   1279: result <= 12'b000011111010;
   1280: result <= 12'b000011111010;
   1281: result <= 12'b000011111010;
   1282: result <= 12'b000011111011;
   1283: result <= 12'b000011111011;
   1284: result <= 12'b000011111011;
   1285: result <= 12'b000011111011;
   1286: result <= 12'b000011111011;
   1287: result <= 12'b000011111100;
   1288: result <= 12'b000011111100;
   1289: result <= 12'b000011111100;
   1290: result <= 12'b000011111100;
   1291: result <= 12'b000011111100;
   1292: result <= 12'b000011111101;
   1293: result <= 12'b000011111101;
   1294: result <= 12'b000011111101;
   1295: result <= 12'b000011111101;
   1296: result <= 12'b000011111101;
   1297: result <= 12'b000011111110;
   1298: result <= 12'b000011111110;
   1299: result <= 12'b000011111110;
   1300: result <= 12'b000011111110;
   1301: result <= 12'b000011111110;
   1302: result <= 12'b000011111110;
   1303: result <= 12'b000011111111;
   1304: result <= 12'b000011111111;
   1305: result <= 12'b000011111111;
   1306: result <= 12'b000011111111;
   1307: result <= 12'b000011111111;
   1308: result <= 12'b000100000000;
   1309: result <= 12'b000100000000;
   1310: result <= 12'b000100000000;
   1311: result <= 12'b000100000000;
   1312: result <= 12'b000100000000;
   1313: result <= 12'b000100000001;
   1314: result <= 12'b000100000001;
   1315: result <= 12'b000100000001;
   1316: result <= 12'b000100000001;
   1317: result <= 12'b000100000001;
   1318: result <= 12'b000100000010;
   1319: result <= 12'b000100000010;
   1320: result <= 12'b000100000010;
   1321: result <= 12'b000100000010;
   1322: result <= 12'b000100000010;
   1323: result <= 12'b000100000011;
   1324: result <= 12'b000100000011;
   1325: result <= 12'b000100000011;
   1326: result <= 12'b000100000011;
   1327: result <= 12'b000100000011;
   1328: result <= 12'b000100000100;
   1329: result <= 12'b000100000100;
   1330: result <= 12'b000100000100;
   1331: result <= 12'b000100000100;
   1332: result <= 12'b000100000100;
   1333: result <= 12'b000100000101;
   1334: result <= 12'b000100000101;
   1335: result <= 12'b000100000101;
   1336: result <= 12'b000100000101;
   1337: result <= 12'b000100000101;
   1338: result <= 12'b000100000101;
   1339: result <= 12'b000100000110;
   1340: result <= 12'b000100000110;
   1341: result <= 12'b000100000110;
   1342: result <= 12'b000100000110;
   1343: result <= 12'b000100000110;
   1344: result <= 12'b000100000111;
   1345: result <= 12'b000100000111;
   1346: result <= 12'b000100000111;
   1347: result <= 12'b000100000111;
   1348: result <= 12'b000100000111;
   1349: result <= 12'b000100001000;
   1350: result <= 12'b000100001000;
   1351: result <= 12'b000100001000;
   1352: result <= 12'b000100001000;
   1353: result <= 12'b000100001000;
   1354: result <= 12'b000100001001;
   1355: result <= 12'b000100001001;
   1356: result <= 12'b000100001001;
   1357: result <= 12'b000100001001;
   1358: result <= 12'b000100001001;
   1359: result <= 12'b000100001010;
   1360: result <= 12'b000100001010;
   1361: result <= 12'b000100001010;
   1362: result <= 12'b000100001010;
   1363: result <= 12'b000100001010;
   1364: result <= 12'b000100001011;
   1365: result <= 12'b000100001011;
   1366: result <= 12'b000100001011;
   1367: result <= 12'b000100001011;
   1368: result <= 12'b000100001011;
   1369: result <= 12'b000100001100;
   1370: result <= 12'b000100001100;
   1371: result <= 12'b000100001100;
   1372: result <= 12'b000100001100;
   1373: result <= 12'b000100001100;
   1374: result <= 12'b000100001101;
   1375: result <= 12'b000100001101;
   1376: result <= 12'b000100001101;
   1377: result <= 12'b000100001101;
   1378: result <= 12'b000100001101;
   1379: result <= 12'b000100001101;
   1380: result <= 12'b000100001110;
   1381: result <= 12'b000100001110;
   1382: result <= 12'b000100001110;
   1383: result <= 12'b000100001110;
   1384: result <= 12'b000100001110;
   1385: result <= 12'b000100001111;
   1386: result <= 12'b000100001111;
   1387: result <= 12'b000100001111;
   1388: result <= 12'b000100001111;
   1389: result <= 12'b000100001111;
   1390: result <= 12'b000100010000;
   1391: result <= 12'b000100010000;
   1392: result <= 12'b000100010000;
   1393: result <= 12'b000100010000;
   1394: result <= 12'b000100010000;
   1395: result <= 12'b000100010001;
   1396: result <= 12'b000100010001;
   1397: result <= 12'b000100010001;
   1398: result <= 12'b000100010001;
   1399: result <= 12'b000100010001;
   1400: result <= 12'b000100010010;
   1401: result <= 12'b000100010010;
   1402: result <= 12'b000100010010;
   1403: result <= 12'b000100010010;
   1404: result <= 12'b000100010010;
   1405: result <= 12'b000100010011;
   1406: result <= 12'b000100010011;
   1407: result <= 12'b000100010011;
   1408: result <= 12'b000100010011;
   1409: result <= 12'b000100010011;
   1410: result <= 12'b000100010100;
   1411: result <= 12'b000100010100;
   1412: result <= 12'b000100010100;
   1413: result <= 12'b000100010100;
   1414: result <= 12'b000100010100;
   1415: result <= 12'b000100010100;
   1416: result <= 12'b000100010101;
   1417: result <= 12'b000100010101;
   1418: result <= 12'b000100010101;
   1419: result <= 12'b000100010101;
   1420: result <= 12'b000100010101;
   1421: result <= 12'b000100010110;
   1422: result <= 12'b000100010110;
   1423: result <= 12'b000100010110;
   1424: result <= 12'b000100010110;
   1425: result <= 12'b000100010110;
   1426: result <= 12'b000100010111;
   1427: result <= 12'b000100010111;
   1428: result <= 12'b000100010111;
   1429: result <= 12'b000100010111;
   1430: result <= 12'b000100010111;
   1431: result <= 12'b000100011000;
   1432: result <= 12'b000100011000;
   1433: result <= 12'b000100011000;
   1434: result <= 12'b000100011000;
   1435: result <= 12'b000100011000;
   1436: result <= 12'b000100011001;
   1437: result <= 12'b000100011001;
   1438: result <= 12'b000100011001;
   1439: result <= 12'b000100011001;
   1440: result <= 12'b000100011001;
   1441: result <= 12'b000100011010;
   1442: result <= 12'b000100011010;
   1443: result <= 12'b000100011010;
   1444: result <= 12'b000100011010;
   1445: result <= 12'b000100011010;
   1446: result <= 12'b000100011011;
   1447: result <= 12'b000100011011;
   1448: result <= 12'b000100011011;
   1449: result <= 12'b000100011011;
   1450: result <= 12'b000100011011;
   1451: result <= 12'b000100011011;
   1452: result <= 12'b000100011100;
   1453: result <= 12'b000100011100;
   1454: result <= 12'b000100011100;
   1455: result <= 12'b000100011100;
   1456: result <= 12'b000100011100;
   1457: result <= 12'b000100011101;
   1458: result <= 12'b000100011101;
   1459: result <= 12'b000100011101;
   1460: result <= 12'b000100011101;
   1461: result <= 12'b000100011101;
   1462: result <= 12'b000100011110;
   1463: result <= 12'b000100011110;
   1464: result <= 12'b000100011110;
   1465: result <= 12'b000100011110;
   1466: result <= 12'b000100011110;
   1467: result <= 12'b000100011111;
   1468: result <= 12'b000100011111;
   1469: result <= 12'b000100011111;
   1470: result <= 12'b000100011111;
   1471: result <= 12'b000100011111;
   1472: result <= 12'b000100100000;
   1473: result <= 12'b000100100000;
   1474: result <= 12'b000100100000;
   1475: result <= 12'b000100100000;
   1476: result <= 12'b000100100000;
   1477: result <= 12'b000100100001;
   1478: result <= 12'b000100100001;
   1479: result <= 12'b000100100001;
   1480: result <= 12'b000100100001;
   1481: result <= 12'b000100100001;
   1482: result <= 12'b000100100010;
   1483: result <= 12'b000100100010;
   1484: result <= 12'b000100100010;
   1485: result <= 12'b000100100010;
   1486: result <= 12'b000100100010;
   1487: result <= 12'b000100100010;
   1488: result <= 12'b000100100011;
   1489: result <= 12'b000100100011;
   1490: result <= 12'b000100100011;
   1491: result <= 12'b000100100011;
   1492: result <= 12'b000100100011;
   1493: result <= 12'b000100100100;
   1494: result <= 12'b000100100100;
   1495: result <= 12'b000100100100;
   1496: result <= 12'b000100100100;
   1497: result <= 12'b000100100100;
   1498: result <= 12'b000100100101;
   1499: result <= 12'b000100100101;
   1500: result <= 12'b000100100101;
   1501: result <= 12'b000100100101;
   1502: result <= 12'b000100100101;
   1503: result <= 12'b000100100110;
   1504: result <= 12'b000100100110;
   1505: result <= 12'b000100100110;
   1506: result <= 12'b000100100110;
   1507: result <= 12'b000100100110;
   1508: result <= 12'b000100100111;
   1509: result <= 12'b000100100111;
   1510: result <= 12'b000100100111;
   1511: result <= 12'b000100100111;
   1512: result <= 12'b000100100111;
   1513: result <= 12'b000100101000;
   1514: result <= 12'b000100101000;
   1515: result <= 12'b000100101000;
   1516: result <= 12'b000100101000;
   1517: result <= 12'b000100101000;
   1518: result <= 12'b000100101001;
   1519: result <= 12'b000100101001;
   1520: result <= 12'b000100101001;
   1521: result <= 12'b000100101001;
   1522: result <= 12'b000100101001;
   1523: result <= 12'b000100101001;
   1524: result <= 12'b000100101010;
   1525: result <= 12'b000100101010;
   1526: result <= 12'b000100101010;
   1527: result <= 12'b000100101010;
   1528: result <= 12'b000100101010;
   1529: result <= 12'b000100101011;
   1530: result <= 12'b000100101011;
   1531: result <= 12'b000100101011;
   1532: result <= 12'b000100101011;
   1533: result <= 12'b000100101011;
   1534: result <= 12'b000100101100;
   1535: result <= 12'b000100101100;
   1536: result <= 12'b000100101100;
   1537: result <= 12'b000100101100;
   1538: result <= 12'b000100101100;
   1539: result <= 12'b000100101101;
   1540: result <= 12'b000100101101;
   1541: result <= 12'b000100101101;
   1542: result <= 12'b000100101101;
   1543: result <= 12'b000100101101;
   1544: result <= 12'b000100101110;
   1545: result <= 12'b000100101110;
   1546: result <= 12'b000100101110;
   1547: result <= 12'b000100101110;
   1548: result <= 12'b000100101110;
   1549: result <= 12'b000100101111;
   1550: result <= 12'b000100101111;
   1551: result <= 12'b000100101111;
   1552: result <= 12'b000100101111;
   1553: result <= 12'b000100101111;
   1554: result <= 12'b000100101111;
   1555: result <= 12'b000100110000;
   1556: result <= 12'b000100110000;
   1557: result <= 12'b000100110000;
   1558: result <= 12'b000100110000;
   1559: result <= 12'b000100110000;
   1560: result <= 12'b000100110001;
   1561: result <= 12'b000100110001;
   1562: result <= 12'b000100110001;
   1563: result <= 12'b000100110001;
   1564: result <= 12'b000100110001;
   1565: result <= 12'b000100110010;
   1566: result <= 12'b000100110010;
   1567: result <= 12'b000100110010;
   1568: result <= 12'b000100110010;
   1569: result <= 12'b000100110010;
   1570: result <= 12'b000100110011;
   1571: result <= 12'b000100110011;
   1572: result <= 12'b000100110011;
   1573: result <= 12'b000100110011;
   1574: result <= 12'b000100110011;
   1575: result <= 12'b000100110100;
   1576: result <= 12'b000100110100;
   1577: result <= 12'b000100110100;
   1578: result <= 12'b000100110100;
   1579: result <= 12'b000100110100;
   1580: result <= 12'b000100110101;
   1581: result <= 12'b000100110101;
   1582: result <= 12'b000100110101;
   1583: result <= 12'b000100110101;
   1584: result <= 12'b000100110101;
   1585: result <= 12'b000100110110;
   1586: result <= 12'b000100110110;
   1587: result <= 12'b000100110110;
   1588: result <= 12'b000100110110;
   1589: result <= 12'b000100110110;
   1590: result <= 12'b000100110110;
   1591: result <= 12'b000100110111;
   1592: result <= 12'b000100110111;
   1593: result <= 12'b000100110111;
   1594: result <= 12'b000100110111;
   1595: result <= 12'b000100110111;
   1596: result <= 12'b000100111000;
   1597: result <= 12'b000100111000;
   1598: result <= 12'b000100111000;
   1599: result <= 12'b000100111000;
   1600: result <= 12'b000100111000;
   1601: result <= 12'b000100111001;
   1602: result <= 12'b000100111001;
   1603: result <= 12'b000100111001;
   1604: result <= 12'b000100111001;
   1605: result <= 12'b000100111001;
   1606: result <= 12'b000100111010;
   1607: result <= 12'b000100111010;
   1608: result <= 12'b000100111010;
   1609: result <= 12'b000100111010;
   1610: result <= 12'b000100111010;
   1611: result <= 12'b000100111011;
   1612: result <= 12'b000100111011;
   1613: result <= 12'b000100111011;
   1614: result <= 12'b000100111011;
   1615: result <= 12'b000100111011;
   1616: result <= 12'b000100111100;
   1617: result <= 12'b000100111100;
   1618: result <= 12'b000100111100;
   1619: result <= 12'b000100111100;
   1620: result <= 12'b000100111100;
   1621: result <= 12'b000100111101;
   1622: result <= 12'b000100111101;
   1623: result <= 12'b000100111101;
   1624: result <= 12'b000100111101;
   1625: result <= 12'b000100111101;
   1626: result <= 12'b000100111101;
   1627: result <= 12'b000100111110;
   1628: result <= 12'b000100111110;
   1629: result <= 12'b000100111110;
   1630: result <= 12'b000100111110;
   1631: result <= 12'b000100111110;
   1632: result <= 12'b000100111111;
   1633: result <= 12'b000100111111;
   1634: result <= 12'b000100111111;
   1635: result <= 12'b000100111111;
   1636: result <= 12'b000100111111;
   1637: result <= 12'b000101000000;
   1638: result <= 12'b000101000000;
   1639: result <= 12'b000101000000;
   1640: result <= 12'b000101000000;
   1641: result <= 12'b000101000000;
   1642: result <= 12'b000101000001;
   1643: result <= 12'b000101000001;
   1644: result <= 12'b000101000001;
   1645: result <= 12'b000101000001;
   1646: result <= 12'b000101000001;
   1647: result <= 12'b000101000010;
   1648: result <= 12'b000101000010;
   1649: result <= 12'b000101000010;
   1650: result <= 12'b000101000010;
   1651: result <= 12'b000101000010;
   1652: result <= 12'b000101000011;
   1653: result <= 12'b000101000011;
   1654: result <= 12'b000101000011;
   1655: result <= 12'b000101000011;
   1656: result <= 12'b000101000011;
   1657: result <= 12'b000101000011;
   1658: result <= 12'b000101000100;
   1659: result <= 12'b000101000100;
   1660: result <= 12'b000101000100;
   1661: result <= 12'b000101000100;
   1662: result <= 12'b000101000100;
   1663: result <= 12'b000101000101;
   1664: result <= 12'b000101000101;
   1665: result <= 12'b000101000101;
   1666: result <= 12'b000101000101;
   1667: result <= 12'b000101000101;
   1668: result <= 12'b000101000110;
   1669: result <= 12'b000101000110;
   1670: result <= 12'b000101000110;
   1671: result <= 12'b000101000110;
   1672: result <= 12'b000101000110;
   1673: result <= 12'b000101000111;
   1674: result <= 12'b000101000111;
   1675: result <= 12'b000101000111;
   1676: result <= 12'b000101000111;
   1677: result <= 12'b000101000111;
   1678: result <= 12'b000101001000;
   1679: result <= 12'b000101001000;
   1680: result <= 12'b000101001000;
   1681: result <= 12'b000101001000;
   1682: result <= 12'b000101001000;
   1683: result <= 12'b000101001001;
   1684: result <= 12'b000101001001;
   1685: result <= 12'b000101001001;
   1686: result <= 12'b000101001001;
   1687: result <= 12'b000101001001;
   1688: result <= 12'b000101001001;
   1689: result <= 12'b000101001010;
   1690: result <= 12'b000101001010;
   1691: result <= 12'b000101001010;
   1692: result <= 12'b000101001010;
   1693: result <= 12'b000101001010;
   1694: result <= 12'b000101001011;
   1695: result <= 12'b000101001011;
   1696: result <= 12'b000101001011;
   1697: result <= 12'b000101001011;
   1698: result <= 12'b000101001011;
   1699: result <= 12'b000101001100;
   1700: result <= 12'b000101001100;
   1701: result <= 12'b000101001100;
   1702: result <= 12'b000101001100;
   1703: result <= 12'b000101001100;
   1704: result <= 12'b000101001101;
   1705: result <= 12'b000101001101;
   1706: result <= 12'b000101001101;
   1707: result <= 12'b000101001101;
   1708: result <= 12'b000101001101;
   1709: result <= 12'b000101001110;
   1710: result <= 12'b000101001110;
   1711: result <= 12'b000101001110;
   1712: result <= 12'b000101001110;
   1713: result <= 12'b000101001110;
   1714: result <= 12'b000101001111;
   1715: result <= 12'b000101001111;
   1716: result <= 12'b000101001111;
   1717: result <= 12'b000101001111;
   1718: result <= 12'b000101001111;
   1719: result <= 12'b000101001111;
   1720: result <= 12'b000101010000;
   1721: result <= 12'b000101010000;
   1722: result <= 12'b000101010000;
   1723: result <= 12'b000101010000;
   1724: result <= 12'b000101010000;
   1725: result <= 12'b000101010001;
   1726: result <= 12'b000101010001;
   1727: result <= 12'b000101010001;
   1728: result <= 12'b000101010001;
   1729: result <= 12'b000101010001;
   1730: result <= 12'b000101010010;
   1731: result <= 12'b000101010010;
   1732: result <= 12'b000101010010;
   1733: result <= 12'b000101010010;
   1734: result <= 12'b000101010010;
   1735: result <= 12'b000101010011;
   1736: result <= 12'b000101010011;
   1737: result <= 12'b000101010011;
   1738: result <= 12'b000101010011;
   1739: result <= 12'b000101010011;
   1740: result <= 12'b000101010100;
   1741: result <= 12'b000101010100;
   1742: result <= 12'b000101010100;
   1743: result <= 12'b000101010100;
   1744: result <= 12'b000101010100;
   1745: result <= 12'b000101010101;
   1746: result <= 12'b000101010101;
   1747: result <= 12'b000101010101;
   1748: result <= 12'b000101010101;
   1749: result <= 12'b000101010101;
   1750: result <= 12'b000101010110;
   1751: result <= 12'b000101010110;
   1752: result <= 12'b000101010110;
   1753: result <= 12'b000101010110;
   1754: result <= 12'b000101010110;
   1755: result <= 12'b000101010110;
   1756: result <= 12'b000101010111;
   1757: result <= 12'b000101010111;
   1758: result <= 12'b000101010111;
   1759: result <= 12'b000101010111;
   1760: result <= 12'b000101010111;
   1761: result <= 12'b000101011000;
   1762: result <= 12'b000101011000;
   1763: result <= 12'b000101011000;
   1764: result <= 12'b000101011000;
   1765: result <= 12'b000101011000;
   1766: result <= 12'b000101011001;
   1767: result <= 12'b000101011001;
   1768: result <= 12'b000101011001;
   1769: result <= 12'b000101011001;
   1770: result <= 12'b000101011001;
   1771: result <= 12'b000101011010;
   1772: result <= 12'b000101011010;
   1773: result <= 12'b000101011010;
   1774: result <= 12'b000101011010;
   1775: result <= 12'b000101011010;
   1776: result <= 12'b000101011011;
   1777: result <= 12'b000101011011;
   1778: result <= 12'b000101011011;
   1779: result <= 12'b000101011011;
   1780: result <= 12'b000101011011;
   1781: result <= 12'b000101011100;
   1782: result <= 12'b000101011100;
   1783: result <= 12'b000101011100;
   1784: result <= 12'b000101011100;
   1785: result <= 12'b000101011100;
   1786: result <= 12'b000101011100;
   1787: result <= 12'b000101011101;
   1788: result <= 12'b000101011101;
   1789: result <= 12'b000101011101;
   1790: result <= 12'b000101011101;
   1791: result <= 12'b000101011101;
   1792: result <= 12'b000101011110;
   1793: result <= 12'b000101011110;
   1794: result <= 12'b000101011110;
   1795: result <= 12'b000101011110;
   1796: result <= 12'b000101011110;
   1797: result <= 12'b000101011111;
   1798: result <= 12'b000101011111;
   1799: result <= 12'b000101011111;
   1800: result <= 12'b000101011111;
   1801: result <= 12'b000101011111;
   1802: result <= 12'b000101100000;
   1803: result <= 12'b000101100000;
   1804: result <= 12'b000101100000;
   1805: result <= 12'b000101100000;
   1806: result <= 12'b000101100000;
   1807: result <= 12'b000101100001;
   1808: result <= 12'b000101100001;
   1809: result <= 12'b000101100001;
   1810: result <= 12'b000101100001;
   1811: result <= 12'b000101100001;
   1812: result <= 12'b000101100001;
   1813: result <= 12'b000101100010;
   1814: result <= 12'b000101100010;
   1815: result <= 12'b000101100010;
   1816: result <= 12'b000101100010;
   1817: result <= 12'b000101100010;
   1818: result <= 12'b000101100011;
   1819: result <= 12'b000101100011;
   1820: result <= 12'b000101100011;
   1821: result <= 12'b000101100011;
   1822: result <= 12'b000101100011;
   1823: result <= 12'b000101100100;
   1824: result <= 12'b000101100100;
   1825: result <= 12'b000101100100;
   1826: result <= 12'b000101100100;
   1827: result <= 12'b000101100100;
   1828: result <= 12'b000101100101;
   1829: result <= 12'b000101100101;
   1830: result <= 12'b000101100101;
   1831: result <= 12'b000101100101;
   1832: result <= 12'b000101100101;
   1833: result <= 12'b000101100110;
   1834: result <= 12'b000101100110;
   1835: result <= 12'b000101100110;
   1836: result <= 12'b000101100110;
   1837: result <= 12'b000101100110;
   1838: result <= 12'b000101100111;
   1839: result <= 12'b000101100111;
   1840: result <= 12'b000101100111;
   1841: result <= 12'b000101100111;
   1842: result <= 12'b000101100111;
   1843: result <= 12'b000101100111;
   1844: result <= 12'b000101101000;
   1845: result <= 12'b000101101000;
   1846: result <= 12'b000101101000;
   1847: result <= 12'b000101101000;
   1848: result <= 12'b000101101000;
   1849: result <= 12'b000101101001;
   1850: result <= 12'b000101101001;
   1851: result <= 12'b000101101001;
   1852: result <= 12'b000101101001;
   1853: result <= 12'b000101101001;
   1854: result <= 12'b000101101010;
   1855: result <= 12'b000101101010;
   1856: result <= 12'b000101101010;
   1857: result <= 12'b000101101010;
   1858: result <= 12'b000101101010;
   1859: result <= 12'b000101101011;
   1860: result <= 12'b000101101011;
   1861: result <= 12'b000101101011;
   1862: result <= 12'b000101101011;
   1863: result <= 12'b000101101011;
   1864: result <= 12'b000101101100;
   1865: result <= 12'b000101101100;
   1866: result <= 12'b000101101100;
   1867: result <= 12'b000101101100;
   1868: result <= 12'b000101101100;
   1869: result <= 12'b000101101101;
   1870: result <= 12'b000101101101;
   1871: result <= 12'b000101101101;
   1872: result <= 12'b000101101101;
   1873: result <= 12'b000101101101;
   1874: result <= 12'b000101101101;
   1875: result <= 12'b000101101110;
   1876: result <= 12'b000101101110;
   1877: result <= 12'b000101101110;
   1878: result <= 12'b000101101110;
   1879: result <= 12'b000101101110;
   1880: result <= 12'b000101101111;
   1881: result <= 12'b000101101111;
   1882: result <= 12'b000101101111;
   1883: result <= 12'b000101101111;
   1884: result <= 12'b000101101111;
   1885: result <= 12'b000101110000;
   1886: result <= 12'b000101110000;
   1887: result <= 12'b000101110000;
   1888: result <= 12'b000101110000;
   1889: result <= 12'b000101110000;
   1890: result <= 12'b000101110001;
   1891: result <= 12'b000101110001;
   1892: result <= 12'b000101110001;
   1893: result <= 12'b000101110001;
   1894: result <= 12'b000101110001;
   1895: result <= 12'b000101110010;
   1896: result <= 12'b000101110010;
   1897: result <= 12'b000101110010;
   1898: result <= 12'b000101110010;
   1899: result <= 12'b000101110010;
   1900: result <= 12'b000101110011;
   1901: result <= 12'b000101110011;
   1902: result <= 12'b000101110011;
   1903: result <= 12'b000101110011;
   1904: result <= 12'b000101110011;
   1905: result <= 12'b000101110011;
   1906: result <= 12'b000101110100;
   1907: result <= 12'b000101110100;
   1908: result <= 12'b000101110100;
   1909: result <= 12'b000101110100;
   1910: result <= 12'b000101110100;
   1911: result <= 12'b000101110101;
   1912: result <= 12'b000101110101;
   1913: result <= 12'b000101110101;
   1914: result <= 12'b000101110101;
   1915: result <= 12'b000101110101;
   1916: result <= 12'b000101110110;
   1917: result <= 12'b000101110110;
   1918: result <= 12'b000101110110;
   1919: result <= 12'b000101110110;
   1920: result <= 12'b000101110110;
   1921: result <= 12'b000101110111;
   1922: result <= 12'b000101110111;
   1923: result <= 12'b000101110111;
   1924: result <= 12'b000101110111;
   1925: result <= 12'b000101110111;
   1926: result <= 12'b000101111000;
   1927: result <= 12'b000101111000;
   1928: result <= 12'b000101111000;
   1929: result <= 12'b000101111000;
   1930: result <= 12'b000101111000;
   1931: result <= 12'b000101111000;
   1932: result <= 12'b000101111001;
   1933: result <= 12'b000101111001;
   1934: result <= 12'b000101111001;
   1935: result <= 12'b000101111001;
   1936: result <= 12'b000101111001;
   1937: result <= 12'b000101111010;
   1938: result <= 12'b000101111010;
   1939: result <= 12'b000101111010;
   1940: result <= 12'b000101111010;
   1941: result <= 12'b000101111010;
   1942: result <= 12'b000101111011;
   1943: result <= 12'b000101111011;
   1944: result <= 12'b000101111011;
   1945: result <= 12'b000101111011;
   1946: result <= 12'b000101111011;
   1947: result <= 12'b000101111100;
   1948: result <= 12'b000101111100;
   1949: result <= 12'b000101111100;
   1950: result <= 12'b000101111100;
   1951: result <= 12'b000101111100;
   1952: result <= 12'b000101111101;
   1953: result <= 12'b000101111101;
   1954: result <= 12'b000101111101;
   1955: result <= 12'b000101111101;
   1956: result <= 12'b000101111101;
   1957: result <= 12'b000101111110;
   1958: result <= 12'b000101111110;
   1959: result <= 12'b000101111110;
   1960: result <= 12'b000101111110;
   1961: result <= 12'b000101111110;
   1962: result <= 12'b000101111110;
   1963: result <= 12'b000101111111;
   1964: result <= 12'b000101111111;
   1965: result <= 12'b000101111111;
   1966: result <= 12'b000101111111;
   1967: result <= 12'b000101111111;
   1968: result <= 12'b000110000000;
   1969: result <= 12'b000110000000;
   1970: result <= 12'b000110000000;
   1971: result <= 12'b000110000000;
   1972: result <= 12'b000110000000;
   1973: result <= 12'b000110000001;
   1974: result <= 12'b000110000001;
   1975: result <= 12'b000110000001;
   1976: result <= 12'b000110000001;
   1977: result <= 12'b000110000001;
   1978: result <= 12'b000110000010;
   1979: result <= 12'b000110000010;
   1980: result <= 12'b000110000010;
   1981: result <= 12'b000110000010;
   1982: result <= 12'b000110000010;
   1983: result <= 12'b000110000011;
   1984: result <= 12'b000110000011;
   1985: result <= 12'b000110000011;
   1986: result <= 12'b000110000011;
   1987: result <= 12'b000110000011;
   1988: result <= 12'b000110000011;
   1989: result <= 12'b000110000100;
   1990: result <= 12'b000110000100;
   1991: result <= 12'b000110000100;
   1992: result <= 12'b000110000100;
   1993: result <= 12'b000110000100;
   1994: result <= 12'b000110000101;
   1995: result <= 12'b000110000101;
   1996: result <= 12'b000110000101;
   1997: result <= 12'b000110000101;
   1998: result <= 12'b000110000101;
   1999: result <= 12'b000110000110;
   2000: result <= 12'b000110000110;
   2001: result <= 12'b000110000110;
   2002: result <= 12'b000110000110;
   2003: result <= 12'b000110000110;
   2004: result <= 12'b000110000111;
   2005: result <= 12'b000110000111;
   2006: result <= 12'b000110000111;
   2007: result <= 12'b000110000111;
   2008: result <= 12'b000110000111;
   2009: result <= 12'b000110001000;
   2010: result <= 12'b000110001000;
   2011: result <= 12'b000110001000;
   2012: result <= 12'b000110001000;
   2013: result <= 12'b000110001000;
   2014: result <= 12'b000110001000;
   2015: result <= 12'b000110001001;
   2016: result <= 12'b000110001001;
   2017: result <= 12'b000110001001;
   2018: result <= 12'b000110001001;
   2019: result <= 12'b000110001001;
   2020: result <= 12'b000110001010;
   2021: result <= 12'b000110001010;
   2022: result <= 12'b000110001010;
   2023: result <= 12'b000110001010;
   2024: result <= 12'b000110001010;
   2025: result <= 12'b000110001011;
   2026: result <= 12'b000110001011;
   2027: result <= 12'b000110001011;
   2028: result <= 12'b000110001011;
   2029: result <= 12'b000110001011;
   2030: result <= 12'b000110001100;
   2031: result <= 12'b000110001100;
   2032: result <= 12'b000110001100;
   2033: result <= 12'b000110001100;
   2034: result <= 12'b000110001100;
   2035: result <= 12'b000110001101;
   2036: result <= 12'b000110001101;
   2037: result <= 12'b000110001101;
   2038: result <= 12'b000110001101;
   2039: result <= 12'b000110001101;
   2040: result <= 12'b000110001110;
   2041: result <= 12'b000110001110;
   2042: result <= 12'b000110001110;
   2043: result <= 12'b000110001110;
   2044: result <= 12'b000110001110;
   2045: result <= 12'b000110001110;
   2046: result <= 12'b000110001111;
   2047: result <= 12'b000110001111;
   2048: result <= 12'b000110001111;
   2049: result <= 12'b000110001111;
   2050: result <= 12'b000110001111;
   2051: result <= 12'b000110010000;
   2052: result <= 12'b000110010000;
   2053: result <= 12'b000110010000;
   2054: result <= 12'b000110010000;
   2055: result <= 12'b000110010000;
   2056: result <= 12'b000110010001;
   2057: result <= 12'b000110010001;
   2058: result <= 12'b000110010001;
   2059: result <= 12'b000110010001;
   2060: result <= 12'b000110010001;
   2061: result <= 12'b000110010010;
   2062: result <= 12'b000110010010;
   2063: result <= 12'b000110010010;
   2064: result <= 12'b000110010010;
   2065: result <= 12'b000110010010;
   2066: result <= 12'b000110010011;
   2067: result <= 12'b000110010011;
   2068: result <= 12'b000110010011;
   2069: result <= 12'b000110010011;
   2070: result <= 12'b000110010011;
   2071: result <= 12'b000110010011;
   2072: result <= 12'b000110010100;
   2073: result <= 12'b000110010100;
   2074: result <= 12'b000110010100;
   2075: result <= 12'b000110010100;
   2076: result <= 12'b000110010100;
   2077: result <= 12'b000110010101;
   2078: result <= 12'b000110010101;
   2079: result <= 12'b000110010101;
   2080: result <= 12'b000110010101;
   2081: result <= 12'b000110010101;
   2082: result <= 12'b000110010110;
   2083: result <= 12'b000110010110;
   2084: result <= 12'b000110010110;
   2085: result <= 12'b000110010110;
   2086: result <= 12'b000110010110;
   2087: result <= 12'b000110010111;
   2088: result <= 12'b000110010111;
   2089: result <= 12'b000110010111;
   2090: result <= 12'b000110010111;
   2091: result <= 12'b000110010111;
   2092: result <= 12'b000110011000;
   2093: result <= 12'b000110011000;
   2094: result <= 12'b000110011000;
   2095: result <= 12'b000110011000;
   2096: result <= 12'b000110011000;
   2097: result <= 12'b000110011000;
   2098: result <= 12'b000110011001;
   2099: result <= 12'b000110011001;
   2100: result <= 12'b000110011001;
   2101: result <= 12'b000110011001;
   2102: result <= 12'b000110011001;
   2103: result <= 12'b000110011010;
   2104: result <= 12'b000110011010;
   2105: result <= 12'b000110011010;
   2106: result <= 12'b000110011010;
   2107: result <= 12'b000110011010;
   2108: result <= 12'b000110011011;
   2109: result <= 12'b000110011011;
   2110: result <= 12'b000110011011;
   2111: result <= 12'b000110011011;
   2112: result <= 12'b000110011011;
   2113: result <= 12'b000110011100;
   2114: result <= 12'b000110011100;
   2115: result <= 12'b000110011100;
   2116: result <= 12'b000110011100;
   2117: result <= 12'b000110011100;
   2118: result <= 12'b000110011101;
   2119: result <= 12'b000110011101;
   2120: result <= 12'b000110011101;
   2121: result <= 12'b000110011101;
   2122: result <= 12'b000110011101;
   2123: result <= 12'b000110011101;
   2124: result <= 12'b000110011110;
   2125: result <= 12'b000110011110;
   2126: result <= 12'b000110011110;
   2127: result <= 12'b000110011110;
   2128: result <= 12'b000110011110;
   2129: result <= 12'b000110011111;
   2130: result <= 12'b000110011111;
   2131: result <= 12'b000110011111;
   2132: result <= 12'b000110011111;
   2133: result <= 12'b000110011111;
   2134: result <= 12'b000110100000;
   2135: result <= 12'b000110100000;
   2136: result <= 12'b000110100000;
   2137: result <= 12'b000110100000;
   2138: result <= 12'b000110100000;
   2139: result <= 12'b000110100001;
   2140: result <= 12'b000110100001;
   2141: result <= 12'b000110100001;
   2142: result <= 12'b000110100001;
   2143: result <= 12'b000110100001;
   2144: result <= 12'b000110100010;
   2145: result <= 12'b000110100010;
   2146: result <= 12'b000110100010;
   2147: result <= 12'b000110100010;
   2148: result <= 12'b000110100010;
   2149: result <= 12'b000110100010;
   2150: result <= 12'b000110100011;
   2151: result <= 12'b000110100011;
   2152: result <= 12'b000110100011;
   2153: result <= 12'b000110100011;
   2154: result <= 12'b000110100011;
   2155: result <= 12'b000110100100;
   2156: result <= 12'b000110100100;
   2157: result <= 12'b000110100100;
   2158: result <= 12'b000110100100;
   2159: result <= 12'b000110100100;
   2160: result <= 12'b000110100101;
   2161: result <= 12'b000110100101;
   2162: result <= 12'b000110100101;
   2163: result <= 12'b000110100101;
   2164: result <= 12'b000110100101;
   2165: result <= 12'b000110100110;
   2166: result <= 12'b000110100110;
   2167: result <= 12'b000110100110;
   2168: result <= 12'b000110100110;
   2169: result <= 12'b000110100110;
   2170: result <= 12'b000110100111;
   2171: result <= 12'b000110100111;
   2172: result <= 12'b000110100111;
   2173: result <= 12'b000110100111;
   2174: result <= 12'b000110100111;
   2175: result <= 12'b000110100111;
   2176: result <= 12'b000110101000;
   2177: result <= 12'b000110101000;
   2178: result <= 12'b000110101000;
   2179: result <= 12'b000110101000;
   2180: result <= 12'b000110101000;
   2181: result <= 12'b000110101001;
   2182: result <= 12'b000110101001;
   2183: result <= 12'b000110101001;
   2184: result <= 12'b000110101001;
   2185: result <= 12'b000110101001;
   2186: result <= 12'b000110101010;
   2187: result <= 12'b000110101010;
   2188: result <= 12'b000110101010;
   2189: result <= 12'b000110101010;
   2190: result <= 12'b000110101010;
   2191: result <= 12'b000110101011;
   2192: result <= 12'b000110101011;
   2193: result <= 12'b000110101011;
   2194: result <= 12'b000110101011;
   2195: result <= 12'b000110101011;
   2196: result <= 12'b000110101100;
   2197: result <= 12'b000110101100;
   2198: result <= 12'b000110101100;
   2199: result <= 12'b000110101100;
   2200: result <= 12'b000110101100;
   2201: result <= 12'b000110101100;
   2202: result <= 12'b000110101101;
   2203: result <= 12'b000110101101;
   2204: result <= 12'b000110101101;
   2205: result <= 12'b000110101101;
   2206: result <= 12'b000110101101;
   2207: result <= 12'b000110101110;
   2208: result <= 12'b000110101110;
   2209: result <= 12'b000110101110;
   2210: result <= 12'b000110101110;
   2211: result <= 12'b000110101110;
   2212: result <= 12'b000110101111;
   2213: result <= 12'b000110101111;
   2214: result <= 12'b000110101111;
   2215: result <= 12'b000110101111;
   2216: result <= 12'b000110101111;
   2217: result <= 12'b000110110000;
   2218: result <= 12'b000110110000;
   2219: result <= 12'b000110110000;
   2220: result <= 12'b000110110000;
   2221: result <= 12'b000110110000;
   2222: result <= 12'b000110110000;
   2223: result <= 12'b000110110001;
   2224: result <= 12'b000110110001;
   2225: result <= 12'b000110110001;
   2226: result <= 12'b000110110001;
   2227: result <= 12'b000110110001;
   2228: result <= 12'b000110110010;
   2229: result <= 12'b000110110010;
   2230: result <= 12'b000110110010;
   2231: result <= 12'b000110110010;
   2232: result <= 12'b000110110010;
   2233: result <= 12'b000110110011;
   2234: result <= 12'b000110110011;
   2235: result <= 12'b000110110011;
   2236: result <= 12'b000110110011;
   2237: result <= 12'b000110110011;
   2238: result <= 12'b000110110100;
   2239: result <= 12'b000110110100;
   2240: result <= 12'b000110110100;
   2241: result <= 12'b000110110100;
   2242: result <= 12'b000110110100;
   2243: result <= 12'b000110110101;
   2244: result <= 12'b000110110101;
   2245: result <= 12'b000110110101;
   2246: result <= 12'b000110110101;
   2247: result <= 12'b000110110101;
   2248: result <= 12'b000110110101;
   2249: result <= 12'b000110110110;
   2250: result <= 12'b000110110110;
   2251: result <= 12'b000110110110;
   2252: result <= 12'b000110110110;
   2253: result <= 12'b000110110110;
   2254: result <= 12'b000110110111;
   2255: result <= 12'b000110110111;
   2256: result <= 12'b000110110111;
   2257: result <= 12'b000110110111;
   2258: result <= 12'b000110110111;
   2259: result <= 12'b000110111000;
   2260: result <= 12'b000110111000;
   2261: result <= 12'b000110111000;
   2262: result <= 12'b000110111000;
   2263: result <= 12'b000110111000;
   2264: result <= 12'b000110111001;
   2265: result <= 12'b000110111001;
   2266: result <= 12'b000110111001;
   2267: result <= 12'b000110111001;
   2268: result <= 12'b000110111001;
   2269: result <= 12'b000110111010;
   2270: result <= 12'b000110111010;
   2271: result <= 12'b000110111010;
   2272: result <= 12'b000110111010;
   2273: result <= 12'b000110111010;
   2274: result <= 12'b000110111010;
   2275: result <= 12'b000110111011;
   2276: result <= 12'b000110111011;
   2277: result <= 12'b000110111011;
   2278: result <= 12'b000110111011;
   2279: result <= 12'b000110111011;
   2280: result <= 12'b000110111100;
   2281: result <= 12'b000110111100;
   2282: result <= 12'b000110111100;
   2283: result <= 12'b000110111100;
   2284: result <= 12'b000110111100;
   2285: result <= 12'b000110111101;
   2286: result <= 12'b000110111101;
   2287: result <= 12'b000110111101;
   2288: result <= 12'b000110111101;
   2289: result <= 12'b000110111101;
   2290: result <= 12'b000110111110;
   2291: result <= 12'b000110111110;
   2292: result <= 12'b000110111110;
   2293: result <= 12'b000110111110;
   2294: result <= 12'b000110111110;
   2295: result <= 12'b000110111110;
   2296: result <= 12'b000110111111;
   2297: result <= 12'b000110111111;
   2298: result <= 12'b000110111111;
   2299: result <= 12'b000110111111;
   2300: result <= 12'b000110111111;
   2301: result <= 12'b000111000000;
   2302: result <= 12'b000111000000;
   2303: result <= 12'b000111000000;
   2304: result <= 12'b000111000000;
   2305: result <= 12'b000111000000;
   2306: result <= 12'b000111000001;
   2307: result <= 12'b000111000001;
   2308: result <= 12'b000111000001;
   2309: result <= 12'b000111000001;
   2310: result <= 12'b000111000001;
   2311: result <= 12'b000111000010;
   2312: result <= 12'b000111000010;
   2313: result <= 12'b000111000010;
   2314: result <= 12'b000111000010;
   2315: result <= 12'b000111000010;
   2316: result <= 12'b000111000011;
   2317: result <= 12'b000111000011;
   2318: result <= 12'b000111000011;
   2319: result <= 12'b000111000011;
   2320: result <= 12'b000111000011;
   2321: result <= 12'b000111000011;
   2322: result <= 12'b000111000100;
   2323: result <= 12'b000111000100;
   2324: result <= 12'b000111000100;
   2325: result <= 12'b000111000100;
   2326: result <= 12'b000111000100;
   2327: result <= 12'b000111000101;
   2328: result <= 12'b000111000101;
   2329: result <= 12'b000111000101;
   2330: result <= 12'b000111000101;
   2331: result <= 12'b000111000101;
   2332: result <= 12'b000111000110;
   2333: result <= 12'b000111000110;
   2334: result <= 12'b000111000110;
   2335: result <= 12'b000111000110;
   2336: result <= 12'b000111000110;
   2337: result <= 12'b000111000111;
   2338: result <= 12'b000111000111;
   2339: result <= 12'b000111000111;
   2340: result <= 12'b000111000111;
   2341: result <= 12'b000111000111;
   2342: result <= 12'b000111000111;
   2343: result <= 12'b000111001000;
   2344: result <= 12'b000111001000;
   2345: result <= 12'b000111001000;
   2346: result <= 12'b000111001000;
   2347: result <= 12'b000111001000;
   2348: result <= 12'b000111001001;
   2349: result <= 12'b000111001001;
   2350: result <= 12'b000111001001;
   2351: result <= 12'b000111001001;
   2352: result <= 12'b000111001001;
   2353: result <= 12'b000111001010;
   2354: result <= 12'b000111001010;
   2355: result <= 12'b000111001010;
   2356: result <= 12'b000111001010;
   2357: result <= 12'b000111001010;
   2358: result <= 12'b000111001011;
   2359: result <= 12'b000111001011;
   2360: result <= 12'b000111001011;
   2361: result <= 12'b000111001011;
   2362: result <= 12'b000111001011;
   2363: result <= 12'b000111001100;
   2364: result <= 12'b000111001100;
   2365: result <= 12'b000111001100;
   2366: result <= 12'b000111001100;
   2367: result <= 12'b000111001100;
   2368: result <= 12'b000111001100;
   2369: result <= 12'b000111001101;
   2370: result <= 12'b000111001101;
   2371: result <= 12'b000111001101;
   2372: result <= 12'b000111001101;
   2373: result <= 12'b000111001101;
   2374: result <= 12'b000111001110;
   2375: result <= 12'b000111001110;
   2376: result <= 12'b000111001110;
   2377: result <= 12'b000111001110;
   2378: result <= 12'b000111001110;
   2379: result <= 12'b000111001111;
   2380: result <= 12'b000111001111;
   2381: result <= 12'b000111001111;
   2382: result <= 12'b000111001111;
   2383: result <= 12'b000111001111;
   2384: result <= 12'b000111010000;
   2385: result <= 12'b000111010000;
   2386: result <= 12'b000111010000;
   2387: result <= 12'b000111010000;
   2388: result <= 12'b000111010000;
   2389: result <= 12'b000111010000;
   2390: result <= 12'b000111010001;
   2391: result <= 12'b000111010001;
   2392: result <= 12'b000111010001;
   2393: result <= 12'b000111010001;
   2394: result <= 12'b000111010001;
   2395: result <= 12'b000111010010;
   2396: result <= 12'b000111010010;
   2397: result <= 12'b000111010010;
   2398: result <= 12'b000111010010;
   2399: result <= 12'b000111010010;
   2400: result <= 12'b000111010011;
   2401: result <= 12'b000111010011;
   2402: result <= 12'b000111010011;
   2403: result <= 12'b000111010011;
   2404: result <= 12'b000111010011;
   2405: result <= 12'b000111010100;
   2406: result <= 12'b000111010100;
   2407: result <= 12'b000111010100;
   2408: result <= 12'b000111010100;
   2409: result <= 12'b000111010100;
   2410: result <= 12'b000111010101;
   2411: result <= 12'b000111010101;
   2412: result <= 12'b000111010101;
   2413: result <= 12'b000111010101;
   2414: result <= 12'b000111010101;
   2415: result <= 12'b000111010101;
   2416: result <= 12'b000111010110;
   2417: result <= 12'b000111010110;
   2418: result <= 12'b000111010110;
   2419: result <= 12'b000111010110;
   2420: result <= 12'b000111010110;
   2421: result <= 12'b000111010111;
   2422: result <= 12'b000111010111;
   2423: result <= 12'b000111010111;
   2424: result <= 12'b000111010111;
   2425: result <= 12'b000111010111;
   2426: result <= 12'b000111011000;
   2427: result <= 12'b000111011000;
   2428: result <= 12'b000111011000;
   2429: result <= 12'b000111011000;
   2430: result <= 12'b000111011000;
   2431: result <= 12'b000111011001;
   2432: result <= 12'b000111011001;
   2433: result <= 12'b000111011001;
   2434: result <= 12'b000111011001;
   2435: result <= 12'b000111011001;
   2436: result <= 12'b000111011001;
   2437: result <= 12'b000111011010;
   2438: result <= 12'b000111011010;
   2439: result <= 12'b000111011010;
   2440: result <= 12'b000111011010;
   2441: result <= 12'b000111011010;
   2442: result <= 12'b000111011011;
   2443: result <= 12'b000111011011;
   2444: result <= 12'b000111011011;
   2445: result <= 12'b000111011011;
   2446: result <= 12'b000111011011;
   2447: result <= 12'b000111011100;
   2448: result <= 12'b000111011100;
   2449: result <= 12'b000111011100;
   2450: result <= 12'b000111011100;
   2451: result <= 12'b000111011100;
   2452: result <= 12'b000111011101;
   2453: result <= 12'b000111011101;
   2454: result <= 12'b000111011101;
   2455: result <= 12'b000111011101;
   2456: result <= 12'b000111011101;
   2457: result <= 12'b000111011101;
   2458: result <= 12'b000111011110;
   2459: result <= 12'b000111011110;
   2460: result <= 12'b000111011110;
   2461: result <= 12'b000111011110;
   2462: result <= 12'b000111011110;
   2463: result <= 12'b000111011111;
   2464: result <= 12'b000111011111;
   2465: result <= 12'b000111011111;
   2466: result <= 12'b000111011111;
   2467: result <= 12'b000111011111;
   2468: result <= 12'b000111100000;
   2469: result <= 12'b000111100000;
   2470: result <= 12'b000111100000;
   2471: result <= 12'b000111100000;
   2472: result <= 12'b000111100000;
   2473: result <= 12'b000111100001;
   2474: result <= 12'b000111100001;
   2475: result <= 12'b000111100001;
   2476: result <= 12'b000111100001;
   2477: result <= 12'b000111100001;
   2478: result <= 12'b000111100001;
   2479: result <= 12'b000111100010;
   2480: result <= 12'b000111100010;
   2481: result <= 12'b000111100010;
   2482: result <= 12'b000111100010;
   2483: result <= 12'b000111100010;
   2484: result <= 12'b000111100011;
   2485: result <= 12'b000111100011;
   2486: result <= 12'b000111100011;
   2487: result <= 12'b000111100011;
   2488: result <= 12'b000111100011;
   2489: result <= 12'b000111100100;
   2490: result <= 12'b000111100100;
   2491: result <= 12'b000111100100;
   2492: result <= 12'b000111100100;
   2493: result <= 12'b000111100100;
   2494: result <= 12'b000111100101;
   2495: result <= 12'b000111100101;
   2496: result <= 12'b000111100101;
   2497: result <= 12'b000111100101;
   2498: result <= 12'b000111100101;
   2499: result <= 12'b000111100101;
   2500: result <= 12'b000111100110;
   2501: result <= 12'b000111100110;
   2502: result <= 12'b000111100110;
   2503: result <= 12'b000111100110;
   2504: result <= 12'b000111100110;
   2505: result <= 12'b000111100111;
   2506: result <= 12'b000111100111;
   2507: result <= 12'b000111100111;
   2508: result <= 12'b000111100111;
   2509: result <= 12'b000111100111;
   2510: result <= 12'b000111101000;
   2511: result <= 12'b000111101000;
   2512: result <= 12'b000111101000;
   2513: result <= 12'b000111101000;
   2514: result <= 12'b000111101000;
   2515: result <= 12'b000111101001;
   2516: result <= 12'b000111101001;
   2517: result <= 12'b000111101001;
   2518: result <= 12'b000111101001;
   2519: result <= 12'b000111101001;
   2520: result <= 12'b000111101010;
   2521: result <= 12'b000111101010;
   2522: result <= 12'b000111101010;
   2523: result <= 12'b000111101010;
   2524: result <= 12'b000111101010;
   2525: result <= 12'b000111101010;
   2526: result <= 12'b000111101011;
   2527: result <= 12'b000111101011;
   2528: result <= 12'b000111101011;
   2529: result <= 12'b000111101011;
   2530: result <= 12'b000111101011;
   2531: result <= 12'b000111101100;
   2532: result <= 12'b000111101100;
   2533: result <= 12'b000111101100;
   2534: result <= 12'b000111101100;
   2535: result <= 12'b000111101100;
   2536: result <= 12'b000111101101;
   2537: result <= 12'b000111101101;
   2538: result <= 12'b000111101101;
   2539: result <= 12'b000111101101;
   2540: result <= 12'b000111101101;
   2541: result <= 12'b000111101110;
   2542: result <= 12'b000111101110;
   2543: result <= 12'b000111101110;
   2544: result <= 12'b000111101110;
   2545: result <= 12'b000111101110;
   2546: result <= 12'b000111101110;
   2547: result <= 12'b000111101111;
   2548: result <= 12'b000111101111;
   2549: result <= 12'b000111101111;
   2550: result <= 12'b000111101111;
   2551: result <= 12'b000111101111;
   2552: result <= 12'b000111110000;
   2553: result <= 12'b000111110000;
   2554: result <= 12'b000111110000;
   2555: result <= 12'b000111110000;
   2556: result <= 12'b000111110000;
   2557: result <= 12'b000111110001;
   2558: result <= 12'b000111110001;
   2559: result <= 12'b000111110001;
   2560: result <= 12'b000111110001;
   2561: result <= 12'b000111110001;
   2562: result <= 12'b000111110010;
   2563: result <= 12'b000111110010;
   2564: result <= 12'b000111110010;
   2565: result <= 12'b000111110010;
   2566: result <= 12'b000111110010;
   2567: result <= 12'b000111110010;
   2568: result <= 12'b000111110011;
   2569: result <= 12'b000111110011;
   2570: result <= 12'b000111110011;
   2571: result <= 12'b000111110011;
   2572: result <= 12'b000111110011;
   2573: result <= 12'b000111110100;
   2574: result <= 12'b000111110100;
   2575: result <= 12'b000111110100;
   2576: result <= 12'b000111110100;
   2577: result <= 12'b000111110100;
   2578: result <= 12'b000111110101;
   2579: result <= 12'b000111110101;
   2580: result <= 12'b000111110101;
   2581: result <= 12'b000111110101;
   2582: result <= 12'b000111110101;
   2583: result <= 12'b000111110110;
   2584: result <= 12'b000111110110;
   2585: result <= 12'b000111110110;
   2586: result <= 12'b000111110110;
   2587: result <= 12'b000111110110;
   2588: result <= 12'b000111110110;
   2589: result <= 12'b000111110111;
   2590: result <= 12'b000111110111;
   2591: result <= 12'b000111110111;
   2592: result <= 12'b000111110111;
   2593: result <= 12'b000111110111;
   2594: result <= 12'b000111111000;
   2595: result <= 12'b000111111000;
   2596: result <= 12'b000111111000;
   2597: result <= 12'b000111111000;
   2598: result <= 12'b000111111000;
   2599: result <= 12'b000111111001;
   2600: result <= 12'b000111111001;
   2601: result <= 12'b000111111001;
   2602: result <= 12'b000111111001;
   2603: result <= 12'b000111111001;
   2604: result <= 12'b000111111001;
   2605: result <= 12'b000111111010;
   2606: result <= 12'b000111111010;
   2607: result <= 12'b000111111010;
   2608: result <= 12'b000111111010;
   2609: result <= 12'b000111111010;
   2610: result <= 12'b000111111011;
   2611: result <= 12'b000111111011;
   2612: result <= 12'b000111111011;
   2613: result <= 12'b000111111011;
   2614: result <= 12'b000111111011;
   2615: result <= 12'b000111111100;
   2616: result <= 12'b000111111100;
   2617: result <= 12'b000111111100;
   2618: result <= 12'b000111111100;
   2619: result <= 12'b000111111100;
   2620: result <= 12'b000111111101;
   2621: result <= 12'b000111111101;
   2622: result <= 12'b000111111101;
   2623: result <= 12'b000111111101;
   2624: result <= 12'b000111111101;
   2625: result <= 12'b000111111101;
   2626: result <= 12'b000111111110;
   2627: result <= 12'b000111111110;
   2628: result <= 12'b000111111110;
   2629: result <= 12'b000111111110;
   2630: result <= 12'b000111111110;
   2631: result <= 12'b000111111111;
   2632: result <= 12'b000111111111;
   2633: result <= 12'b000111111111;
   2634: result <= 12'b000111111111;
   2635: result <= 12'b000111111111;
   2636: result <= 12'b001000000000;
   2637: result <= 12'b001000000000;
   2638: result <= 12'b001000000000;
   2639: result <= 12'b001000000000;
   2640: result <= 12'b001000000000;
   2641: result <= 12'b001000000001;
   2642: result <= 12'b001000000001;
   2643: result <= 12'b001000000001;
   2644: result <= 12'b001000000001;
   2645: result <= 12'b001000000001;
   2646: result <= 12'b001000000001;
   2647: result <= 12'b001000000010;
   2648: result <= 12'b001000000010;
   2649: result <= 12'b001000000010;
   2650: result <= 12'b001000000010;
   2651: result <= 12'b001000000010;
   2652: result <= 12'b001000000011;
   2653: result <= 12'b001000000011;
   2654: result <= 12'b001000000011;
   2655: result <= 12'b001000000011;
   2656: result <= 12'b001000000011;
   2657: result <= 12'b001000000100;
   2658: result <= 12'b001000000100;
   2659: result <= 12'b001000000100;
   2660: result <= 12'b001000000100;
   2661: result <= 12'b001000000100;
   2662: result <= 12'b001000000101;
   2663: result <= 12'b001000000101;
   2664: result <= 12'b001000000101;
   2665: result <= 12'b001000000101;
   2666: result <= 12'b001000000101;
   2667: result <= 12'b001000000101;
   2668: result <= 12'b001000000110;
   2669: result <= 12'b001000000110;
   2670: result <= 12'b001000000110;
   2671: result <= 12'b001000000110;
   2672: result <= 12'b001000000110;
   2673: result <= 12'b001000000111;
   2674: result <= 12'b001000000111;
   2675: result <= 12'b001000000111;
   2676: result <= 12'b001000000111;
   2677: result <= 12'b001000000111;
   2678: result <= 12'b001000001000;
   2679: result <= 12'b001000001000;
   2680: result <= 12'b001000001000;
   2681: result <= 12'b001000001000;
   2682: result <= 12'b001000001000;
   2683: result <= 12'b001000001001;
   2684: result <= 12'b001000001001;
   2685: result <= 12'b001000001001;
   2686: result <= 12'b001000001001;
   2687: result <= 12'b001000001001;
   2688: result <= 12'b001000001001;
   2689: result <= 12'b001000001010;
   2690: result <= 12'b001000001010;
   2691: result <= 12'b001000001010;
   2692: result <= 12'b001000001010;
   2693: result <= 12'b001000001010;
   2694: result <= 12'b001000001011;
   2695: result <= 12'b001000001011;
   2696: result <= 12'b001000001011;
   2697: result <= 12'b001000001011;
   2698: result <= 12'b001000001011;
   2699: result <= 12'b001000001100;
   2700: result <= 12'b001000001100;
   2701: result <= 12'b001000001100;
   2702: result <= 12'b001000001100;
   2703: result <= 12'b001000001100;
   2704: result <= 12'b001000001101;
   2705: result <= 12'b001000001101;
   2706: result <= 12'b001000001101;
   2707: result <= 12'b001000001101;
   2708: result <= 12'b001000001101;
   2709: result <= 12'b001000001101;
   2710: result <= 12'b001000001110;
   2711: result <= 12'b001000001110;
   2712: result <= 12'b001000001110;
   2713: result <= 12'b001000001110;
   2714: result <= 12'b001000001110;
   2715: result <= 12'b001000001111;
   2716: result <= 12'b001000001111;
   2717: result <= 12'b001000001111;
   2718: result <= 12'b001000001111;
   2719: result <= 12'b001000001111;
   2720: result <= 12'b001000010000;
   2721: result <= 12'b001000010000;
   2722: result <= 12'b001000010000;
   2723: result <= 12'b001000010000;
   2724: result <= 12'b001000010000;
   2725: result <= 12'b001000010000;
   2726: result <= 12'b001000010001;
   2727: result <= 12'b001000010001;
   2728: result <= 12'b001000010001;
   2729: result <= 12'b001000010001;
   2730: result <= 12'b001000010001;
   2731: result <= 12'b001000010010;
   2732: result <= 12'b001000010010;
   2733: result <= 12'b001000010010;
   2734: result <= 12'b001000010010;
   2735: result <= 12'b001000010010;
   2736: result <= 12'b001000010011;
   2737: result <= 12'b001000010011;
   2738: result <= 12'b001000010011;
   2739: result <= 12'b001000010011;
   2740: result <= 12'b001000010011;
   2741: result <= 12'b001000010100;
   2742: result <= 12'b001000010100;
   2743: result <= 12'b001000010100;
   2744: result <= 12'b001000010100;
   2745: result <= 12'b001000010100;
   2746: result <= 12'b001000010100;
   2747: result <= 12'b001000010101;
   2748: result <= 12'b001000010101;
   2749: result <= 12'b001000010101;
   2750: result <= 12'b001000010101;
   2751: result <= 12'b001000010101;
   2752: result <= 12'b001000010110;
   2753: result <= 12'b001000010110;
   2754: result <= 12'b001000010110;
   2755: result <= 12'b001000010110;
   2756: result <= 12'b001000010110;
   2757: result <= 12'b001000010111;
   2758: result <= 12'b001000010111;
   2759: result <= 12'b001000010111;
   2760: result <= 12'b001000010111;
   2761: result <= 12'b001000010111;
   2762: result <= 12'b001000011000;
   2763: result <= 12'b001000011000;
   2764: result <= 12'b001000011000;
   2765: result <= 12'b001000011000;
   2766: result <= 12'b001000011000;
   2767: result <= 12'b001000011000;
   2768: result <= 12'b001000011001;
   2769: result <= 12'b001000011001;
   2770: result <= 12'b001000011001;
   2771: result <= 12'b001000011001;
   2772: result <= 12'b001000011001;
   2773: result <= 12'b001000011010;
   2774: result <= 12'b001000011010;
   2775: result <= 12'b001000011010;
   2776: result <= 12'b001000011010;
   2777: result <= 12'b001000011010;
   2778: result <= 12'b001000011011;
   2779: result <= 12'b001000011011;
   2780: result <= 12'b001000011011;
   2781: result <= 12'b001000011011;
   2782: result <= 12'b001000011011;
   2783: result <= 12'b001000011011;
   2784: result <= 12'b001000011100;
   2785: result <= 12'b001000011100;
   2786: result <= 12'b001000011100;
   2787: result <= 12'b001000011100;
   2788: result <= 12'b001000011100;
   2789: result <= 12'b001000011101;
   2790: result <= 12'b001000011101;
   2791: result <= 12'b001000011101;
   2792: result <= 12'b001000011101;
   2793: result <= 12'b001000011101;
   2794: result <= 12'b001000011110;
   2795: result <= 12'b001000011110;
   2796: result <= 12'b001000011110;
   2797: result <= 12'b001000011110;
   2798: result <= 12'b001000011110;
   2799: result <= 12'b001000011111;
   2800: result <= 12'b001000011111;
   2801: result <= 12'b001000011111;
   2802: result <= 12'b001000011111;
   2803: result <= 12'b001000011111;
   2804: result <= 12'b001000011111;
   2805: result <= 12'b001000100000;
   2806: result <= 12'b001000100000;
   2807: result <= 12'b001000100000;
   2808: result <= 12'b001000100000;
   2809: result <= 12'b001000100000;
   2810: result <= 12'b001000100001;
   2811: result <= 12'b001000100001;
   2812: result <= 12'b001000100001;
   2813: result <= 12'b001000100001;
   2814: result <= 12'b001000100001;
   2815: result <= 12'b001000100010;
   2816: result <= 12'b001000100010;
   2817: result <= 12'b001000100010;
   2818: result <= 12'b001000100010;
   2819: result <= 12'b001000100010;
   2820: result <= 12'b001000100010;
   2821: result <= 12'b001000100011;
   2822: result <= 12'b001000100011;
   2823: result <= 12'b001000100011;
   2824: result <= 12'b001000100011;
   2825: result <= 12'b001000100011;
   2826: result <= 12'b001000100100;
   2827: result <= 12'b001000100100;
   2828: result <= 12'b001000100100;
   2829: result <= 12'b001000100100;
   2830: result <= 12'b001000100100;
   2831: result <= 12'b001000100101;
   2832: result <= 12'b001000100101;
   2833: result <= 12'b001000100101;
   2834: result <= 12'b001000100101;
   2835: result <= 12'b001000100101;
   2836: result <= 12'b001000100110;
   2837: result <= 12'b001000100110;
   2838: result <= 12'b001000100110;
   2839: result <= 12'b001000100110;
   2840: result <= 12'b001000100110;
   2841: result <= 12'b001000100110;
   2842: result <= 12'b001000100111;
   2843: result <= 12'b001000100111;
   2844: result <= 12'b001000100111;
   2845: result <= 12'b001000100111;
   2846: result <= 12'b001000100111;
   2847: result <= 12'b001000101000;
   2848: result <= 12'b001000101000;
   2849: result <= 12'b001000101000;
   2850: result <= 12'b001000101000;
   2851: result <= 12'b001000101000;
   2852: result <= 12'b001000101001;
   2853: result <= 12'b001000101001;
   2854: result <= 12'b001000101001;
   2855: result <= 12'b001000101001;
   2856: result <= 12'b001000101001;
   2857: result <= 12'b001000101001;
   2858: result <= 12'b001000101010;
   2859: result <= 12'b001000101010;
   2860: result <= 12'b001000101010;
   2861: result <= 12'b001000101010;
   2862: result <= 12'b001000101010;
   2863: result <= 12'b001000101011;
   2864: result <= 12'b001000101011;
   2865: result <= 12'b001000101011;
   2866: result <= 12'b001000101011;
   2867: result <= 12'b001000101011;
   2868: result <= 12'b001000101100;
   2869: result <= 12'b001000101100;
   2870: result <= 12'b001000101100;
   2871: result <= 12'b001000101100;
   2872: result <= 12'b001000101100;
   2873: result <= 12'b001000101101;
   2874: result <= 12'b001000101101;
   2875: result <= 12'b001000101101;
   2876: result <= 12'b001000101101;
   2877: result <= 12'b001000101101;
   2878: result <= 12'b001000101101;
   2879: result <= 12'b001000101110;
   2880: result <= 12'b001000101110;
   2881: result <= 12'b001000101110;
   2882: result <= 12'b001000101110;
   2883: result <= 12'b001000101110;
   2884: result <= 12'b001000101111;
   2885: result <= 12'b001000101111;
   2886: result <= 12'b001000101111;
   2887: result <= 12'b001000101111;
   2888: result <= 12'b001000101111;
   2889: result <= 12'b001000110000;
   2890: result <= 12'b001000110000;
   2891: result <= 12'b001000110000;
   2892: result <= 12'b001000110000;
   2893: result <= 12'b001000110000;
   2894: result <= 12'b001000110000;
   2895: result <= 12'b001000110001;
   2896: result <= 12'b001000110001;
   2897: result <= 12'b001000110001;
   2898: result <= 12'b001000110001;
   2899: result <= 12'b001000110001;
   2900: result <= 12'b001000110010;
   2901: result <= 12'b001000110010;
   2902: result <= 12'b001000110010;
   2903: result <= 12'b001000110010;
   2904: result <= 12'b001000110010;
   2905: result <= 12'b001000110011;
   2906: result <= 12'b001000110011;
   2907: result <= 12'b001000110011;
   2908: result <= 12'b001000110011;
   2909: result <= 12'b001000110011;
   2910: result <= 12'b001000110011;
   2911: result <= 12'b001000110100;
   2912: result <= 12'b001000110100;
   2913: result <= 12'b001000110100;
   2914: result <= 12'b001000110100;
   2915: result <= 12'b001000110100;
   2916: result <= 12'b001000110101;
   2917: result <= 12'b001000110101;
   2918: result <= 12'b001000110101;
   2919: result <= 12'b001000110101;
   2920: result <= 12'b001000110101;
   2921: result <= 12'b001000110110;
   2922: result <= 12'b001000110110;
   2923: result <= 12'b001000110110;
   2924: result <= 12'b001000110110;
   2925: result <= 12'b001000110110;
   2926: result <= 12'b001000110111;
   2927: result <= 12'b001000110111;
   2928: result <= 12'b001000110111;
   2929: result <= 12'b001000110111;
   2930: result <= 12'b001000110111;
   2931: result <= 12'b001000110111;
   2932: result <= 12'b001000111000;
   2933: result <= 12'b001000111000;
   2934: result <= 12'b001000111000;
   2935: result <= 12'b001000111000;
   2936: result <= 12'b001000111000;
   2937: result <= 12'b001000111001;
   2938: result <= 12'b001000111001;
   2939: result <= 12'b001000111001;
   2940: result <= 12'b001000111001;
   2941: result <= 12'b001000111001;
   2942: result <= 12'b001000111010;
   2943: result <= 12'b001000111010;
   2944: result <= 12'b001000111010;
   2945: result <= 12'b001000111010;
   2946: result <= 12'b001000111010;
   2947: result <= 12'b001000111010;
   2948: result <= 12'b001000111011;
   2949: result <= 12'b001000111011;
   2950: result <= 12'b001000111011;
   2951: result <= 12'b001000111011;
   2952: result <= 12'b001000111011;
   2953: result <= 12'b001000111100;
   2954: result <= 12'b001000111100;
   2955: result <= 12'b001000111100;
   2956: result <= 12'b001000111100;
   2957: result <= 12'b001000111100;
   2958: result <= 12'b001000111101;
   2959: result <= 12'b001000111101;
   2960: result <= 12'b001000111101;
   2961: result <= 12'b001000111101;
   2962: result <= 12'b001000111101;
   2963: result <= 12'b001000111101;
   2964: result <= 12'b001000111110;
   2965: result <= 12'b001000111110;
   2966: result <= 12'b001000111110;
   2967: result <= 12'b001000111110;
   2968: result <= 12'b001000111110;
   2969: result <= 12'b001000111111;
   2970: result <= 12'b001000111111;
   2971: result <= 12'b001000111111;
   2972: result <= 12'b001000111111;
   2973: result <= 12'b001000111111;
   2974: result <= 12'b001001000000;
   2975: result <= 12'b001001000000;
   2976: result <= 12'b001001000000;
   2977: result <= 12'b001001000000;
   2978: result <= 12'b001001000000;
   2979: result <= 12'b001001000001;
   2980: result <= 12'b001001000001;
   2981: result <= 12'b001001000001;
   2982: result <= 12'b001001000001;
   2983: result <= 12'b001001000001;
   2984: result <= 12'b001001000001;
   2985: result <= 12'b001001000010;
   2986: result <= 12'b001001000010;
   2987: result <= 12'b001001000010;
   2988: result <= 12'b001001000010;
   2989: result <= 12'b001001000010;
   2990: result <= 12'b001001000011;
   2991: result <= 12'b001001000011;
   2992: result <= 12'b001001000011;
   2993: result <= 12'b001001000011;
   2994: result <= 12'b001001000011;
   2995: result <= 12'b001001000100;
   2996: result <= 12'b001001000100;
   2997: result <= 12'b001001000100;
   2998: result <= 12'b001001000100;
   2999: result <= 12'b001001000100;
   3000: result <= 12'b001001000100;
   3001: result <= 12'b001001000101;
   3002: result <= 12'b001001000101;
   3003: result <= 12'b001001000101;
   3004: result <= 12'b001001000101;
   3005: result <= 12'b001001000101;
   3006: result <= 12'b001001000110;
   3007: result <= 12'b001001000110;
   3008: result <= 12'b001001000110;
   3009: result <= 12'b001001000110;
   3010: result <= 12'b001001000110;
   3011: result <= 12'b001001000111;
   3012: result <= 12'b001001000111;
   3013: result <= 12'b001001000111;
   3014: result <= 12'b001001000111;
   3015: result <= 12'b001001000111;
   3016: result <= 12'b001001000111;
   3017: result <= 12'b001001001000;
   3018: result <= 12'b001001001000;
   3019: result <= 12'b001001001000;
   3020: result <= 12'b001001001000;
   3021: result <= 12'b001001001000;
   3022: result <= 12'b001001001001;
   3023: result <= 12'b001001001001;
   3024: result <= 12'b001001001001;
   3025: result <= 12'b001001001001;
   3026: result <= 12'b001001001001;
   3027: result <= 12'b001001001010;
   3028: result <= 12'b001001001010;
   3029: result <= 12'b001001001010;
   3030: result <= 12'b001001001010;
   3031: result <= 12'b001001001010;
   3032: result <= 12'b001001001010;
   3033: result <= 12'b001001001011;
   3034: result <= 12'b001001001011;
   3035: result <= 12'b001001001011;
   3036: result <= 12'b001001001011;
   3037: result <= 12'b001001001011;
   3038: result <= 12'b001001001100;
   3039: result <= 12'b001001001100;
   3040: result <= 12'b001001001100;
   3041: result <= 12'b001001001100;
   3042: result <= 12'b001001001100;
   3043: result <= 12'b001001001101;
   3044: result <= 12'b001001001101;
   3045: result <= 12'b001001001101;
   3046: result <= 12'b001001001101;
   3047: result <= 12'b001001001101;
   3048: result <= 12'b001001001101;
   3049: result <= 12'b001001001110;
   3050: result <= 12'b001001001110;
   3051: result <= 12'b001001001110;
   3052: result <= 12'b001001001110;
   3053: result <= 12'b001001001110;
   3054: result <= 12'b001001001111;
   3055: result <= 12'b001001001111;
   3056: result <= 12'b001001001111;
   3057: result <= 12'b001001001111;
   3058: result <= 12'b001001001111;
   3059: result <= 12'b001001010000;
   3060: result <= 12'b001001010000;
   3061: result <= 12'b001001010000;
   3062: result <= 12'b001001010000;
   3063: result <= 12'b001001010000;
   3064: result <= 12'b001001010000;
   3065: result <= 12'b001001010001;
   3066: result <= 12'b001001010001;
   3067: result <= 12'b001001010001;
   3068: result <= 12'b001001010001;
   3069: result <= 12'b001001010001;
   3070: result <= 12'b001001010010;
   3071: result <= 12'b001001010010;
   3072: result <= 12'b001001010010;
   3073: result <= 12'b001001010010;
   3074: result <= 12'b001001010010;
   3075: result <= 12'b001001010011;
   3076: result <= 12'b001001010011;
   3077: result <= 12'b001001010011;
   3078: result <= 12'b001001010011;
   3079: result <= 12'b001001010011;
   3080: result <= 12'b001001010100;
   3081: result <= 12'b001001010100;
   3082: result <= 12'b001001010100;
   3083: result <= 12'b001001010100;
   3084: result <= 12'b001001010100;
   3085: result <= 12'b001001010100;
   3086: result <= 12'b001001010101;
   3087: result <= 12'b001001010101;
   3088: result <= 12'b001001010101;
   3089: result <= 12'b001001010101;
   3090: result <= 12'b001001010101;
   3091: result <= 12'b001001010110;
   3092: result <= 12'b001001010110;
   3093: result <= 12'b001001010110;
   3094: result <= 12'b001001010110;
   3095: result <= 12'b001001010110;
   3096: result <= 12'b001001010111;
   3097: result <= 12'b001001010111;
   3098: result <= 12'b001001010111;
   3099: result <= 12'b001001010111;
   3100: result <= 12'b001001010111;
   3101: result <= 12'b001001010111;
   3102: result <= 12'b001001011000;
   3103: result <= 12'b001001011000;
   3104: result <= 12'b001001011000;
   3105: result <= 12'b001001011000;
   3106: result <= 12'b001001011000;
   3107: result <= 12'b001001011001;
   3108: result <= 12'b001001011001;
   3109: result <= 12'b001001011001;
   3110: result <= 12'b001001011001;
   3111: result <= 12'b001001011001;
   3112: result <= 12'b001001011010;
   3113: result <= 12'b001001011010;
   3114: result <= 12'b001001011010;
   3115: result <= 12'b001001011010;
   3116: result <= 12'b001001011010;
   3117: result <= 12'b001001011010;
   3118: result <= 12'b001001011011;
   3119: result <= 12'b001001011011;
   3120: result <= 12'b001001011011;
   3121: result <= 12'b001001011011;
   3122: result <= 12'b001001011011;
   3123: result <= 12'b001001011100;
   3124: result <= 12'b001001011100;
   3125: result <= 12'b001001011100;
   3126: result <= 12'b001001011100;
   3127: result <= 12'b001001011100;
   3128: result <= 12'b001001011101;
   3129: result <= 12'b001001011101;
   3130: result <= 12'b001001011101;
   3131: result <= 12'b001001011101;
   3132: result <= 12'b001001011101;
   3133: result <= 12'b001001011101;
   3134: result <= 12'b001001011110;
   3135: result <= 12'b001001011110;
   3136: result <= 12'b001001011110;
   3137: result <= 12'b001001011110;
   3138: result <= 12'b001001011110;
   3139: result <= 12'b001001011111;
   3140: result <= 12'b001001011111;
   3141: result <= 12'b001001011111;
   3142: result <= 12'b001001011111;
   3143: result <= 12'b001001011111;
   3144: result <= 12'b001001100000;
   3145: result <= 12'b001001100000;
   3146: result <= 12'b001001100000;
   3147: result <= 12'b001001100000;
   3148: result <= 12'b001001100000;
   3149: result <= 12'b001001100000;
   3150: result <= 12'b001001100001;
   3151: result <= 12'b001001100001;
   3152: result <= 12'b001001100001;
   3153: result <= 12'b001001100001;
   3154: result <= 12'b001001100001;
   3155: result <= 12'b001001100010;
   3156: result <= 12'b001001100010;
   3157: result <= 12'b001001100010;
   3158: result <= 12'b001001100010;
   3159: result <= 12'b001001100010;
   3160: result <= 12'b001001100011;
   3161: result <= 12'b001001100011;
   3162: result <= 12'b001001100011;
   3163: result <= 12'b001001100011;
   3164: result <= 12'b001001100011;
   3165: result <= 12'b001001100011;
   3166: result <= 12'b001001100100;
   3167: result <= 12'b001001100100;
   3168: result <= 12'b001001100100;
   3169: result <= 12'b001001100100;
   3170: result <= 12'b001001100100;
   3171: result <= 12'b001001100101;
   3172: result <= 12'b001001100101;
   3173: result <= 12'b001001100101;
   3174: result <= 12'b001001100101;
   3175: result <= 12'b001001100101;
   3176: result <= 12'b001001100110;
   3177: result <= 12'b001001100110;
   3178: result <= 12'b001001100110;
   3179: result <= 12'b001001100110;
   3180: result <= 12'b001001100110;
   3181: result <= 12'b001001100110;
   3182: result <= 12'b001001100111;
   3183: result <= 12'b001001100111;
   3184: result <= 12'b001001100111;
   3185: result <= 12'b001001100111;
   3186: result <= 12'b001001100111;
   3187: result <= 12'b001001101000;
   3188: result <= 12'b001001101000;
   3189: result <= 12'b001001101000;
   3190: result <= 12'b001001101000;
   3191: result <= 12'b001001101000;
   3192: result <= 12'b001001101001;
   3193: result <= 12'b001001101001;
   3194: result <= 12'b001001101001;
   3195: result <= 12'b001001101001;
   3196: result <= 12'b001001101001;
   3197: result <= 12'b001001101001;
   3198: result <= 12'b001001101010;
   3199: result <= 12'b001001101010;
   3200: result <= 12'b001001101010;
   3201: result <= 12'b001001101010;
   3202: result <= 12'b001001101010;
   3203: result <= 12'b001001101011;
   3204: result <= 12'b001001101011;
   3205: result <= 12'b001001101011;
   3206: result <= 12'b001001101011;
   3207: result <= 12'b001001101011;
   3208: result <= 12'b001001101100;
   3209: result <= 12'b001001101100;
   3210: result <= 12'b001001101100;
   3211: result <= 12'b001001101100;
   3212: result <= 12'b001001101100;
   3213: result <= 12'b001001101100;
   3214: result <= 12'b001001101101;
   3215: result <= 12'b001001101101;
   3216: result <= 12'b001001101101;
   3217: result <= 12'b001001101101;
   3218: result <= 12'b001001101101;
   3219: result <= 12'b001001101110;
   3220: result <= 12'b001001101110;
   3221: result <= 12'b001001101110;
   3222: result <= 12'b001001101110;
   3223: result <= 12'b001001101110;
   3224: result <= 12'b001001101110;
   3225: result <= 12'b001001101111;
   3226: result <= 12'b001001101111;
   3227: result <= 12'b001001101111;
   3228: result <= 12'b001001101111;
   3229: result <= 12'b001001101111;
   3230: result <= 12'b001001110000;
   3231: result <= 12'b001001110000;
   3232: result <= 12'b001001110000;
   3233: result <= 12'b001001110000;
   3234: result <= 12'b001001110000;
   3235: result <= 12'b001001110001;
   3236: result <= 12'b001001110001;
   3237: result <= 12'b001001110001;
   3238: result <= 12'b001001110001;
   3239: result <= 12'b001001110001;
   3240: result <= 12'b001001110001;
   3241: result <= 12'b001001110010;
   3242: result <= 12'b001001110010;
   3243: result <= 12'b001001110010;
   3244: result <= 12'b001001110010;
   3245: result <= 12'b001001110010;
   3246: result <= 12'b001001110011;
   3247: result <= 12'b001001110011;
   3248: result <= 12'b001001110011;
   3249: result <= 12'b001001110011;
   3250: result <= 12'b001001110011;
   3251: result <= 12'b001001110100;
   3252: result <= 12'b001001110100;
   3253: result <= 12'b001001110100;
   3254: result <= 12'b001001110100;
   3255: result <= 12'b001001110100;
   3256: result <= 12'b001001110100;
   3257: result <= 12'b001001110101;
   3258: result <= 12'b001001110101;
   3259: result <= 12'b001001110101;
   3260: result <= 12'b001001110101;
   3261: result <= 12'b001001110101;
   3262: result <= 12'b001001110110;
   3263: result <= 12'b001001110110;
   3264: result <= 12'b001001110110;
   3265: result <= 12'b001001110110;
   3266: result <= 12'b001001110110;
   3267: result <= 12'b001001110111;
   3268: result <= 12'b001001110111;
   3269: result <= 12'b001001110111;
   3270: result <= 12'b001001110111;
   3271: result <= 12'b001001110111;
   3272: result <= 12'b001001110111;
   3273: result <= 12'b001001111000;
   3274: result <= 12'b001001111000;
   3275: result <= 12'b001001111000;
   3276: result <= 12'b001001111000;
   3277: result <= 12'b001001111000;
   3278: result <= 12'b001001111001;
   3279: result <= 12'b001001111001;
   3280: result <= 12'b001001111001;
   3281: result <= 12'b001001111001;
   3282: result <= 12'b001001111001;
   3283: result <= 12'b001001111010;
   3284: result <= 12'b001001111010;
   3285: result <= 12'b001001111010;
   3286: result <= 12'b001001111010;
   3287: result <= 12'b001001111010;
   3288: result <= 12'b001001111010;
   3289: result <= 12'b001001111011;
   3290: result <= 12'b001001111011;
   3291: result <= 12'b001001111011;
   3292: result <= 12'b001001111011;
   3293: result <= 12'b001001111011;
   3294: result <= 12'b001001111100;
   3295: result <= 12'b001001111100;
   3296: result <= 12'b001001111100;
   3297: result <= 12'b001001111100;
   3298: result <= 12'b001001111100;
   3299: result <= 12'b001001111101;
   3300: result <= 12'b001001111101;
   3301: result <= 12'b001001111101;
   3302: result <= 12'b001001111101;
   3303: result <= 12'b001001111101;
   3304: result <= 12'b001001111101;
   3305: result <= 12'b001001111110;
   3306: result <= 12'b001001111110;
   3307: result <= 12'b001001111110;
   3308: result <= 12'b001001111110;
   3309: result <= 12'b001001111110;
   3310: result <= 12'b001001111111;
   3311: result <= 12'b001001111111;
   3312: result <= 12'b001001111111;
   3313: result <= 12'b001001111111;
   3314: result <= 12'b001001111111;
   3315: result <= 12'b001001111111;
   3316: result <= 12'b001010000000;
   3317: result <= 12'b001010000000;
   3318: result <= 12'b001010000000;
   3319: result <= 12'b001010000000;
   3320: result <= 12'b001010000000;
   3321: result <= 12'b001010000001;
   3322: result <= 12'b001010000001;
   3323: result <= 12'b001010000001;
   3324: result <= 12'b001010000001;
   3325: result <= 12'b001010000001;
   3326: result <= 12'b001010000010;
   3327: result <= 12'b001010000010;
   3328: result <= 12'b001010000010;
   3329: result <= 12'b001010000010;
   3330: result <= 12'b001010000010;
   3331: result <= 12'b001010000010;
   3332: result <= 12'b001010000011;
   3333: result <= 12'b001010000011;
   3334: result <= 12'b001010000011;
   3335: result <= 12'b001010000011;
   3336: result <= 12'b001010000011;
   3337: result <= 12'b001010000100;
   3338: result <= 12'b001010000100;
   3339: result <= 12'b001010000100;
   3340: result <= 12'b001010000100;
   3341: result <= 12'b001010000100;
   3342: result <= 12'b001010000101;
   3343: result <= 12'b001010000101;
   3344: result <= 12'b001010000101;
   3345: result <= 12'b001010000101;
   3346: result <= 12'b001010000101;
   3347: result <= 12'b001010000101;
   3348: result <= 12'b001010000110;
   3349: result <= 12'b001010000110;
   3350: result <= 12'b001010000110;
   3351: result <= 12'b001010000110;
   3352: result <= 12'b001010000110;
   3353: result <= 12'b001010000111;
   3354: result <= 12'b001010000111;
   3355: result <= 12'b001010000111;
   3356: result <= 12'b001010000111;
   3357: result <= 12'b001010000111;
   3358: result <= 12'b001010001000;
   3359: result <= 12'b001010001000;
   3360: result <= 12'b001010001000;
   3361: result <= 12'b001010001000;
   3362: result <= 12'b001010001000;
   3363: result <= 12'b001010001000;
   3364: result <= 12'b001010001001;
   3365: result <= 12'b001010001001;
   3366: result <= 12'b001010001001;
   3367: result <= 12'b001010001001;
   3368: result <= 12'b001010001001;
   3369: result <= 12'b001010001010;
   3370: result <= 12'b001010001010;
   3371: result <= 12'b001010001010;
   3372: result <= 12'b001010001010;
   3373: result <= 12'b001010001010;
   3374: result <= 12'b001010001010;
   3375: result <= 12'b001010001011;
   3376: result <= 12'b001010001011;
   3377: result <= 12'b001010001011;
   3378: result <= 12'b001010001011;
   3379: result <= 12'b001010001011;
   3380: result <= 12'b001010001100;
   3381: result <= 12'b001010001100;
   3382: result <= 12'b001010001100;
   3383: result <= 12'b001010001100;
   3384: result <= 12'b001010001100;
   3385: result <= 12'b001010001101;
   3386: result <= 12'b001010001101;
   3387: result <= 12'b001010001101;
   3388: result <= 12'b001010001101;
   3389: result <= 12'b001010001101;
   3390: result <= 12'b001010001101;
   3391: result <= 12'b001010001110;
   3392: result <= 12'b001010001110;
   3393: result <= 12'b001010001110;
   3394: result <= 12'b001010001110;
   3395: result <= 12'b001010001110;
   3396: result <= 12'b001010001111;
   3397: result <= 12'b001010001111;
   3398: result <= 12'b001010001111;
   3399: result <= 12'b001010001111;
   3400: result <= 12'b001010001111;
   3401: result <= 12'b001010010000;
   3402: result <= 12'b001010010000;
   3403: result <= 12'b001010010000;
   3404: result <= 12'b001010010000;
   3405: result <= 12'b001010010000;
   3406: result <= 12'b001010010000;
   3407: result <= 12'b001010010001;
   3408: result <= 12'b001010010001;
   3409: result <= 12'b001010010001;
   3410: result <= 12'b001010010001;
   3411: result <= 12'b001010010001;
   3412: result <= 12'b001010010010;
   3413: result <= 12'b001010010010;
   3414: result <= 12'b001010010010;
   3415: result <= 12'b001010010010;
   3416: result <= 12'b001010010010;
   3417: result <= 12'b001010010010;
   3418: result <= 12'b001010010011;
   3419: result <= 12'b001010010011;
   3420: result <= 12'b001010010011;
   3421: result <= 12'b001010010011;
   3422: result <= 12'b001010010011;
   3423: result <= 12'b001010010100;
   3424: result <= 12'b001010010100;
   3425: result <= 12'b001010010100;
   3426: result <= 12'b001010010100;
   3427: result <= 12'b001010010100;
   3428: result <= 12'b001010010101;
   3429: result <= 12'b001010010101;
   3430: result <= 12'b001010010101;
   3431: result <= 12'b001010010101;
   3432: result <= 12'b001010010101;
   3433: result <= 12'b001010010101;
   3434: result <= 12'b001010010110;
   3435: result <= 12'b001010010110;
   3436: result <= 12'b001010010110;
   3437: result <= 12'b001010010110;
   3438: result <= 12'b001010010110;
   3439: result <= 12'b001010010111;
   3440: result <= 12'b001010010111;
   3441: result <= 12'b001010010111;
   3442: result <= 12'b001010010111;
   3443: result <= 12'b001010010111;
   3444: result <= 12'b001010011000;
   3445: result <= 12'b001010011000;
   3446: result <= 12'b001010011000;
   3447: result <= 12'b001010011000;
   3448: result <= 12'b001010011000;
   3449: result <= 12'b001010011000;
   3450: result <= 12'b001010011001;
   3451: result <= 12'b001010011001;
   3452: result <= 12'b001010011001;
   3453: result <= 12'b001010011001;
   3454: result <= 12'b001010011001;
   3455: result <= 12'b001010011010;
   3456: result <= 12'b001010011010;
   3457: result <= 12'b001010011010;
   3458: result <= 12'b001010011010;
   3459: result <= 12'b001010011010;
   3460: result <= 12'b001010011010;
   3461: result <= 12'b001010011011;
   3462: result <= 12'b001010011011;
   3463: result <= 12'b001010011011;
   3464: result <= 12'b001010011011;
   3465: result <= 12'b001010011011;
   3466: result <= 12'b001010011100;
   3467: result <= 12'b001010011100;
   3468: result <= 12'b001010011100;
   3469: result <= 12'b001010011100;
   3470: result <= 12'b001010011100;
   3471: result <= 12'b001010011101;
   3472: result <= 12'b001010011101;
   3473: result <= 12'b001010011101;
   3474: result <= 12'b001010011101;
   3475: result <= 12'b001010011101;
   3476: result <= 12'b001010011101;
   3477: result <= 12'b001010011110;
   3478: result <= 12'b001010011110;
   3479: result <= 12'b001010011110;
   3480: result <= 12'b001010011110;
   3481: result <= 12'b001010011110;
   3482: result <= 12'b001010011111;
   3483: result <= 12'b001010011111;
   3484: result <= 12'b001010011111;
   3485: result <= 12'b001010011111;
   3486: result <= 12'b001010011111;
   3487: result <= 12'b001010011111;
   3488: result <= 12'b001010100000;
   3489: result <= 12'b001010100000;
   3490: result <= 12'b001010100000;
   3491: result <= 12'b001010100000;
   3492: result <= 12'b001010100000;
   3493: result <= 12'b001010100001;
   3494: result <= 12'b001010100001;
   3495: result <= 12'b001010100001;
   3496: result <= 12'b001010100001;
   3497: result <= 12'b001010100001;
   3498: result <= 12'b001010100010;
   3499: result <= 12'b001010100010;
   3500: result <= 12'b001010100010;
   3501: result <= 12'b001010100010;
   3502: result <= 12'b001010100010;
   3503: result <= 12'b001010100010;
   3504: result <= 12'b001010100011;
   3505: result <= 12'b001010100011;
   3506: result <= 12'b001010100011;
   3507: result <= 12'b001010100011;
   3508: result <= 12'b001010100011;
   3509: result <= 12'b001010100100;
   3510: result <= 12'b001010100100;
   3511: result <= 12'b001010100100;
   3512: result <= 12'b001010100100;
   3513: result <= 12'b001010100100;
   3514: result <= 12'b001010100100;
   3515: result <= 12'b001010100101;
   3516: result <= 12'b001010100101;
   3517: result <= 12'b001010100101;
   3518: result <= 12'b001010100101;
   3519: result <= 12'b001010100101;
   3520: result <= 12'b001010100110;
   3521: result <= 12'b001010100110;
   3522: result <= 12'b001010100110;
   3523: result <= 12'b001010100110;
   3524: result <= 12'b001010100110;
   3525: result <= 12'b001010100111;
   3526: result <= 12'b001010100111;
   3527: result <= 12'b001010100111;
   3528: result <= 12'b001010100111;
   3529: result <= 12'b001010100111;
   3530: result <= 12'b001010100111;
   3531: result <= 12'b001010101000;
   3532: result <= 12'b001010101000;
   3533: result <= 12'b001010101000;
   3534: result <= 12'b001010101000;
   3535: result <= 12'b001010101000;
   3536: result <= 12'b001010101001;
   3537: result <= 12'b001010101001;
   3538: result <= 12'b001010101001;
   3539: result <= 12'b001010101001;
   3540: result <= 12'b001010101001;
   3541: result <= 12'b001010101001;
   3542: result <= 12'b001010101010;
   3543: result <= 12'b001010101010;
   3544: result <= 12'b001010101010;
   3545: result <= 12'b001010101010;
   3546: result <= 12'b001010101010;
   3547: result <= 12'b001010101011;
   3548: result <= 12'b001010101011;
   3549: result <= 12'b001010101011;
   3550: result <= 12'b001010101011;
   3551: result <= 12'b001010101011;
   3552: result <= 12'b001010101100;
   3553: result <= 12'b001010101100;
   3554: result <= 12'b001010101100;
   3555: result <= 12'b001010101100;
   3556: result <= 12'b001010101100;
   3557: result <= 12'b001010101100;
   3558: result <= 12'b001010101101;
   3559: result <= 12'b001010101101;
   3560: result <= 12'b001010101101;
   3561: result <= 12'b001010101101;
   3562: result <= 12'b001010101101;
   3563: result <= 12'b001010101110;
   3564: result <= 12'b001010101110;
   3565: result <= 12'b001010101110;
   3566: result <= 12'b001010101110;
   3567: result <= 12'b001010101110;
   3568: result <= 12'b001010101110;
   3569: result <= 12'b001010101111;
   3570: result <= 12'b001010101111;
   3571: result <= 12'b001010101111;
   3572: result <= 12'b001010101111;
   3573: result <= 12'b001010101111;
   3574: result <= 12'b001010110000;
   3575: result <= 12'b001010110000;
   3576: result <= 12'b001010110000;
   3577: result <= 12'b001010110000;
   3578: result <= 12'b001010110000;
   3579: result <= 12'b001010110001;
   3580: result <= 12'b001010110001;
   3581: result <= 12'b001010110001;
   3582: result <= 12'b001010110001;
   3583: result <= 12'b001010110001;
   3584: result <= 12'b001010110001;
   3585: result <= 12'b001010110010;
   3586: result <= 12'b001010110010;
   3587: result <= 12'b001010110010;
   3588: result <= 12'b001010110010;
   3589: result <= 12'b001010110010;
   3590: result <= 12'b001010110011;
   3591: result <= 12'b001010110011;
   3592: result <= 12'b001010110011;
   3593: result <= 12'b001010110011;
   3594: result <= 12'b001010110011;
   3595: result <= 12'b001010110011;
   3596: result <= 12'b001010110100;
   3597: result <= 12'b001010110100;
   3598: result <= 12'b001010110100;
   3599: result <= 12'b001010110100;
   3600: result <= 12'b001010110100;
   3601: result <= 12'b001010110101;
   3602: result <= 12'b001010110101;
   3603: result <= 12'b001010110101;
   3604: result <= 12'b001010110101;
   3605: result <= 12'b001010110101;
   3606: result <= 12'b001010110110;
   3607: result <= 12'b001010110110;
   3608: result <= 12'b001010110110;
   3609: result <= 12'b001010110110;
   3610: result <= 12'b001010110110;
   3611: result <= 12'b001010110110;
   3612: result <= 12'b001010110111;
   3613: result <= 12'b001010110111;
   3614: result <= 12'b001010110111;
   3615: result <= 12'b001010110111;
   3616: result <= 12'b001010110111;
   3617: result <= 12'b001010111000;
   3618: result <= 12'b001010111000;
   3619: result <= 12'b001010111000;
   3620: result <= 12'b001010111000;
   3621: result <= 12'b001010111000;
   3622: result <= 12'b001010111000;
   3623: result <= 12'b001010111001;
   3624: result <= 12'b001010111001;
   3625: result <= 12'b001010111001;
   3626: result <= 12'b001010111001;
   3627: result <= 12'b001010111001;
   3628: result <= 12'b001010111010;
   3629: result <= 12'b001010111010;
   3630: result <= 12'b001010111010;
   3631: result <= 12'b001010111010;
   3632: result <= 12'b001010111010;
   3633: result <= 12'b001010111011;
   3634: result <= 12'b001010111011;
   3635: result <= 12'b001010111011;
   3636: result <= 12'b001010111011;
   3637: result <= 12'b001010111011;
   3638: result <= 12'b001010111011;
   3639: result <= 12'b001010111100;
   3640: result <= 12'b001010111100;
   3641: result <= 12'b001010111100;
   3642: result <= 12'b001010111100;
   3643: result <= 12'b001010111100;
   3644: result <= 12'b001010111101;
   3645: result <= 12'b001010111101;
   3646: result <= 12'b001010111101;
   3647: result <= 12'b001010111101;
   3648: result <= 12'b001010111101;
   3649: result <= 12'b001010111101;
   3650: result <= 12'b001010111110;
   3651: result <= 12'b001010111110;
   3652: result <= 12'b001010111110;
   3653: result <= 12'b001010111110;
   3654: result <= 12'b001010111110;
   3655: result <= 12'b001010111111;
   3656: result <= 12'b001010111111;
   3657: result <= 12'b001010111111;
   3658: result <= 12'b001010111111;
   3659: result <= 12'b001010111111;
   3660: result <= 12'b001010111111;
   3661: result <= 12'b001011000000;
   3662: result <= 12'b001011000000;
   3663: result <= 12'b001011000000;
   3664: result <= 12'b001011000000;
   3665: result <= 12'b001011000000;
   3666: result <= 12'b001011000001;
   3667: result <= 12'b001011000001;
   3668: result <= 12'b001011000001;
   3669: result <= 12'b001011000001;
   3670: result <= 12'b001011000001;
   3671: result <= 12'b001011000010;
   3672: result <= 12'b001011000010;
   3673: result <= 12'b001011000010;
   3674: result <= 12'b001011000010;
   3675: result <= 12'b001011000010;
   3676: result <= 12'b001011000010;
   3677: result <= 12'b001011000011;
   3678: result <= 12'b001011000011;
   3679: result <= 12'b001011000011;
   3680: result <= 12'b001011000011;
   3681: result <= 12'b001011000011;
   3682: result <= 12'b001011000100;
   3683: result <= 12'b001011000100;
   3684: result <= 12'b001011000100;
   3685: result <= 12'b001011000100;
   3686: result <= 12'b001011000100;
   3687: result <= 12'b001011000100;
   3688: result <= 12'b001011000101;
   3689: result <= 12'b001011000101;
   3690: result <= 12'b001011000101;
   3691: result <= 12'b001011000101;
   3692: result <= 12'b001011000101;
   3693: result <= 12'b001011000110;
   3694: result <= 12'b001011000110;
   3695: result <= 12'b001011000110;
   3696: result <= 12'b001011000110;
   3697: result <= 12'b001011000110;
   3698: result <= 12'b001011000110;
   3699: result <= 12'b001011000111;
   3700: result <= 12'b001011000111;
   3701: result <= 12'b001011000111;
   3702: result <= 12'b001011000111;
   3703: result <= 12'b001011000111;
   3704: result <= 12'b001011001000;
   3705: result <= 12'b001011001000;
   3706: result <= 12'b001011001000;
   3707: result <= 12'b001011001000;
   3708: result <= 12'b001011001000;
   3709: result <= 12'b001011001001;
   3710: result <= 12'b001011001001;
   3711: result <= 12'b001011001001;
   3712: result <= 12'b001011001001;
   3713: result <= 12'b001011001001;
   3714: result <= 12'b001011001001;
   3715: result <= 12'b001011001010;
   3716: result <= 12'b001011001010;
   3717: result <= 12'b001011001010;
   3718: result <= 12'b001011001010;
   3719: result <= 12'b001011001010;
   3720: result <= 12'b001011001011;
   3721: result <= 12'b001011001011;
   3722: result <= 12'b001011001011;
   3723: result <= 12'b001011001011;
   3724: result <= 12'b001011001011;
   3725: result <= 12'b001011001011;
   3726: result <= 12'b001011001100;
   3727: result <= 12'b001011001100;
   3728: result <= 12'b001011001100;
   3729: result <= 12'b001011001100;
   3730: result <= 12'b001011001100;
   3731: result <= 12'b001011001101;
   3732: result <= 12'b001011001101;
   3733: result <= 12'b001011001101;
   3734: result <= 12'b001011001101;
   3735: result <= 12'b001011001101;
   3736: result <= 12'b001011001101;
   3737: result <= 12'b001011001110;
   3738: result <= 12'b001011001110;
   3739: result <= 12'b001011001110;
   3740: result <= 12'b001011001110;
   3741: result <= 12'b001011001110;
   3742: result <= 12'b001011001111;
   3743: result <= 12'b001011001111;
   3744: result <= 12'b001011001111;
   3745: result <= 12'b001011001111;
   3746: result <= 12'b001011001111;
   3747: result <= 12'b001011001111;
   3748: result <= 12'b001011010000;
   3749: result <= 12'b001011010000;
   3750: result <= 12'b001011010000;
   3751: result <= 12'b001011010000;
   3752: result <= 12'b001011010000;
   3753: result <= 12'b001011010001;
   3754: result <= 12'b001011010001;
   3755: result <= 12'b001011010001;
   3756: result <= 12'b001011010001;
   3757: result <= 12'b001011010001;
   3758: result <= 12'b001011010010;
   3759: result <= 12'b001011010010;
   3760: result <= 12'b001011010010;
   3761: result <= 12'b001011010010;
   3762: result <= 12'b001011010010;
   3763: result <= 12'b001011010010;
   3764: result <= 12'b001011010011;
   3765: result <= 12'b001011010011;
   3766: result <= 12'b001011010011;
   3767: result <= 12'b001011010011;
   3768: result <= 12'b001011010011;
   3769: result <= 12'b001011010100;
   3770: result <= 12'b001011010100;
   3771: result <= 12'b001011010100;
   3772: result <= 12'b001011010100;
   3773: result <= 12'b001011010100;
   3774: result <= 12'b001011010100;
   3775: result <= 12'b001011010101;
   3776: result <= 12'b001011010101;
   3777: result <= 12'b001011010101;
   3778: result <= 12'b001011010101;
   3779: result <= 12'b001011010101;
   3780: result <= 12'b001011010110;
   3781: result <= 12'b001011010110;
   3782: result <= 12'b001011010110;
   3783: result <= 12'b001011010110;
   3784: result <= 12'b001011010110;
   3785: result <= 12'b001011010110;
   3786: result <= 12'b001011010111;
   3787: result <= 12'b001011010111;
   3788: result <= 12'b001011010111;
   3789: result <= 12'b001011010111;
   3790: result <= 12'b001011010111;
   3791: result <= 12'b001011011000;
   3792: result <= 12'b001011011000;
   3793: result <= 12'b001011011000;
   3794: result <= 12'b001011011000;
   3795: result <= 12'b001011011000;
   3796: result <= 12'b001011011000;
   3797: result <= 12'b001011011001;
   3798: result <= 12'b001011011001;
   3799: result <= 12'b001011011001;
   3800: result <= 12'b001011011001;
   3801: result <= 12'b001011011001;
   3802: result <= 12'b001011011010;
   3803: result <= 12'b001011011010;
   3804: result <= 12'b001011011010;
   3805: result <= 12'b001011011010;
   3806: result <= 12'b001011011010;
   3807: result <= 12'b001011011011;
   3808: result <= 12'b001011011011;
   3809: result <= 12'b001011011011;
   3810: result <= 12'b001011011011;
   3811: result <= 12'b001011011011;
   3812: result <= 12'b001011011011;
   3813: result <= 12'b001011011100;
   3814: result <= 12'b001011011100;
   3815: result <= 12'b001011011100;
   3816: result <= 12'b001011011100;
   3817: result <= 12'b001011011100;
   3818: result <= 12'b001011011101;
   3819: result <= 12'b001011011101;
   3820: result <= 12'b001011011101;
   3821: result <= 12'b001011011101;
   3822: result <= 12'b001011011101;
   3823: result <= 12'b001011011101;
   3824: result <= 12'b001011011110;
   3825: result <= 12'b001011011110;
   3826: result <= 12'b001011011110;
   3827: result <= 12'b001011011110;
   3828: result <= 12'b001011011110;
   3829: result <= 12'b001011011111;
   3830: result <= 12'b001011011111;
   3831: result <= 12'b001011011111;
   3832: result <= 12'b001011011111;
   3833: result <= 12'b001011011111;
   3834: result <= 12'b001011011111;
   3835: result <= 12'b001011100000;
   3836: result <= 12'b001011100000;
   3837: result <= 12'b001011100000;
   3838: result <= 12'b001011100000;
   3839: result <= 12'b001011100000;
   3840: result <= 12'b001011100001;
   3841: result <= 12'b001011100001;
   3842: result <= 12'b001011100001;
   3843: result <= 12'b001011100001;
   3844: result <= 12'b001011100001;
   3845: result <= 12'b001011100001;
   3846: result <= 12'b001011100010;
   3847: result <= 12'b001011100010;
   3848: result <= 12'b001011100010;
   3849: result <= 12'b001011100010;
   3850: result <= 12'b001011100010;
   3851: result <= 12'b001011100011;
   3852: result <= 12'b001011100011;
   3853: result <= 12'b001011100011;
   3854: result <= 12'b001011100011;
   3855: result <= 12'b001011100011;
   3856: result <= 12'b001011100011;
   3857: result <= 12'b001011100100;
   3858: result <= 12'b001011100100;
   3859: result <= 12'b001011100100;
   3860: result <= 12'b001011100100;
   3861: result <= 12'b001011100100;
   3862: result <= 12'b001011100101;
   3863: result <= 12'b001011100101;
   3864: result <= 12'b001011100101;
   3865: result <= 12'b001011100101;
   3866: result <= 12'b001011100101;
   3867: result <= 12'b001011100110;
   3868: result <= 12'b001011100110;
   3869: result <= 12'b001011100110;
   3870: result <= 12'b001011100110;
   3871: result <= 12'b001011100110;
   3872: result <= 12'b001011100110;
   3873: result <= 12'b001011100111;
   3874: result <= 12'b001011100111;
   3875: result <= 12'b001011100111;
   3876: result <= 12'b001011100111;
   3877: result <= 12'b001011100111;
   3878: result <= 12'b001011101000;
   3879: result <= 12'b001011101000;
   3880: result <= 12'b001011101000;
   3881: result <= 12'b001011101000;
   3882: result <= 12'b001011101000;
   3883: result <= 12'b001011101000;
   3884: result <= 12'b001011101001;
   3885: result <= 12'b001011101001;
   3886: result <= 12'b001011101001;
   3887: result <= 12'b001011101001;
   3888: result <= 12'b001011101001;
   3889: result <= 12'b001011101010;
   3890: result <= 12'b001011101010;
   3891: result <= 12'b001011101010;
   3892: result <= 12'b001011101010;
   3893: result <= 12'b001011101010;
   3894: result <= 12'b001011101010;
   3895: result <= 12'b001011101011;
   3896: result <= 12'b001011101011;
   3897: result <= 12'b001011101011;
   3898: result <= 12'b001011101011;
   3899: result <= 12'b001011101011;
   3900: result <= 12'b001011101100;
   3901: result <= 12'b001011101100;
   3902: result <= 12'b001011101100;
   3903: result <= 12'b001011101100;
   3904: result <= 12'b001011101100;
   3905: result <= 12'b001011101100;
   3906: result <= 12'b001011101101;
   3907: result <= 12'b001011101101;
   3908: result <= 12'b001011101101;
   3909: result <= 12'b001011101101;
   3910: result <= 12'b001011101101;
   3911: result <= 12'b001011101110;
   3912: result <= 12'b001011101110;
   3913: result <= 12'b001011101110;
   3914: result <= 12'b001011101110;
   3915: result <= 12'b001011101110;
   3916: result <= 12'b001011101110;
   3917: result <= 12'b001011101111;
   3918: result <= 12'b001011101111;
   3919: result <= 12'b001011101111;
   3920: result <= 12'b001011101111;
   3921: result <= 12'b001011101111;
   3922: result <= 12'b001011110000;
   3923: result <= 12'b001011110000;
   3924: result <= 12'b001011110000;
   3925: result <= 12'b001011110000;
   3926: result <= 12'b001011110000;
   3927: result <= 12'b001011110000;
   3928: result <= 12'b001011110001;
   3929: result <= 12'b001011110001;
   3930: result <= 12'b001011110001;
   3931: result <= 12'b001011110001;
   3932: result <= 12'b001011110001;
   3933: result <= 12'b001011110010;
   3934: result <= 12'b001011110010;
   3935: result <= 12'b001011110010;
   3936: result <= 12'b001011110010;
   3937: result <= 12'b001011110010;
   3938: result <= 12'b001011110010;
   3939: result <= 12'b001011110011;
   3940: result <= 12'b001011110011;
   3941: result <= 12'b001011110011;
   3942: result <= 12'b001011110011;
   3943: result <= 12'b001011110011;
   3944: result <= 12'b001011110100;
   3945: result <= 12'b001011110100;
   3946: result <= 12'b001011110100;
   3947: result <= 12'b001011110100;
   3948: result <= 12'b001011110100;
   3949: result <= 12'b001011110100;
   3950: result <= 12'b001011110101;
   3951: result <= 12'b001011110101;
   3952: result <= 12'b001011110101;
   3953: result <= 12'b001011110101;
   3954: result <= 12'b001011110101;
   3955: result <= 12'b001011110110;
   3956: result <= 12'b001011110110;
   3957: result <= 12'b001011110110;
   3958: result <= 12'b001011110110;
   3959: result <= 12'b001011110110;
   3960: result <= 12'b001011110110;
   3961: result <= 12'b001011110111;
   3962: result <= 12'b001011110111;
   3963: result <= 12'b001011110111;
   3964: result <= 12'b001011110111;
   3965: result <= 12'b001011110111;
   3966: result <= 12'b001011111000;
   3967: result <= 12'b001011111000;
   3968: result <= 12'b001011111000;
   3969: result <= 12'b001011111000;
   3970: result <= 12'b001011111000;
   3971: result <= 12'b001011111001;
   3972: result <= 12'b001011111001;
   3973: result <= 12'b001011111001;
   3974: result <= 12'b001011111001;
   3975: result <= 12'b001011111001;
   3976: result <= 12'b001011111001;
   3977: result <= 12'b001011111010;
   3978: result <= 12'b001011111010;
   3979: result <= 12'b001011111010;
   3980: result <= 12'b001011111010;
   3981: result <= 12'b001011111010;
   3982: result <= 12'b001011111011;
   3983: result <= 12'b001011111011;
   3984: result <= 12'b001011111011;
   3985: result <= 12'b001011111011;
   3986: result <= 12'b001011111011;
   3987: result <= 12'b001011111011;
   3988: result <= 12'b001011111100;
   3989: result <= 12'b001011111100;
   3990: result <= 12'b001011111100;
   3991: result <= 12'b001011111100;
   3992: result <= 12'b001011111100;
   3993: result <= 12'b001011111101;
   3994: result <= 12'b001011111101;
   3995: result <= 12'b001011111101;
   3996: result <= 12'b001011111101;
   3997: result <= 12'b001011111101;
   3998: result <= 12'b001011111101;
   3999: result <= 12'b001011111110;
   4000: result <= 12'b001011111110;
   4001: result <= 12'b001011111110;
   4002: result <= 12'b001011111110;
   4003: result <= 12'b001011111110;
   4004: result <= 12'b001011111111;
   4005: result <= 12'b001011111111;
   4006: result <= 12'b001011111111;
   4007: result <= 12'b001011111111;
   4008: result <= 12'b001011111111;
   4009: result <= 12'b001011111111;
   4010: result <= 12'b001100000000;
   4011: result <= 12'b001100000000;
   4012: result <= 12'b001100000000;
   4013: result <= 12'b001100000000;
   4014: result <= 12'b001100000000;
   4015: result <= 12'b001100000001;
   4016: result <= 12'b001100000001;
   4017: result <= 12'b001100000001;
   4018: result <= 12'b001100000001;
   4019: result <= 12'b001100000001;
   4020: result <= 12'b001100000001;
   4021: result <= 12'b001100000010;
   4022: result <= 12'b001100000010;
   4023: result <= 12'b001100000010;
   4024: result <= 12'b001100000010;
   4025: result <= 12'b001100000010;
   4026: result <= 12'b001100000011;
   4027: result <= 12'b001100000011;
   4028: result <= 12'b001100000011;
   4029: result <= 12'b001100000011;
   4030: result <= 12'b001100000011;
   4031: result <= 12'b001100000011;
   4032: result <= 12'b001100000100;
   4033: result <= 12'b001100000100;
   4034: result <= 12'b001100000100;
   4035: result <= 12'b001100000100;
   4036: result <= 12'b001100000100;
   4037: result <= 12'b001100000101;
   4038: result <= 12'b001100000101;
   4039: result <= 12'b001100000101;
   4040: result <= 12'b001100000101;
   4041: result <= 12'b001100000101;
   4042: result <= 12'b001100000101;
   4043: result <= 12'b001100000110;
   4044: result <= 12'b001100000110;
   4045: result <= 12'b001100000110;
   4046: result <= 12'b001100000110;
   4047: result <= 12'b001100000110;
   4048: result <= 12'b001100000111;
   4049: result <= 12'b001100000111;
   4050: result <= 12'b001100000111;
   4051: result <= 12'b001100000111;
   4052: result <= 12'b001100000111;
   4053: result <= 12'b001100000111;
   4054: result <= 12'b001100001000;
   4055: result <= 12'b001100001000;
   4056: result <= 12'b001100001000;
   4057: result <= 12'b001100001000;
   4058: result <= 12'b001100001000;
   4059: result <= 12'b001100001001;
   4060: result <= 12'b001100001001;
   4061: result <= 12'b001100001001;
   4062: result <= 12'b001100001001;
   4063: result <= 12'b001100001001;
   4064: result <= 12'b001100001001;
   4065: result <= 12'b001100001010;
   4066: result <= 12'b001100001010;
   4067: result <= 12'b001100001010;
   4068: result <= 12'b001100001010;
   4069: result <= 12'b001100001010;
   4070: result <= 12'b001100001011;
   4071: result <= 12'b001100001011;
   4072: result <= 12'b001100001011;
   4073: result <= 12'b001100001011;
   4074: result <= 12'b001100001011;
   4075: result <= 12'b001100001011;
   4076: result <= 12'b001100001100;
   4077: result <= 12'b001100001100;
   4078: result <= 12'b001100001100;
   4079: result <= 12'b001100001100;
   4080: result <= 12'b001100001100;
   4081: result <= 12'b001100001101;
   4082: result <= 12'b001100001101;
   4083: result <= 12'b001100001101;
   4084: result <= 12'b001100001101;
   4085: result <= 12'b001100001101;
   4086: result <= 12'b001100001101;
   4087: result <= 12'b001100001110;
   4088: result <= 12'b001100001110;
   4089: result <= 12'b001100001110;
   4090: result <= 12'b001100001110;
   4091: result <= 12'b001100001110;
   4092: result <= 12'b001100001111;
   4093: result <= 12'b001100001111;
   4094: result <= 12'b001100001111;
   4095: result <= 12'b001100001111;
   4096: result <= 12'b001100001111;
   4097: result <= 12'b001100001111;
   4098: result <= 12'b001100010000;
   4099: result <= 12'b001100010000;
   4100: result <= 12'b001100010000;
   4101: result <= 12'b001100010000;
   4102: result <= 12'b001100010000;
   4103: result <= 12'b001100010001;
   4104: result <= 12'b001100010001;
   4105: result <= 12'b001100010001;
   4106: result <= 12'b001100010001;
   4107: result <= 12'b001100010001;
   4108: result <= 12'b001100010001;
   4109: result <= 12'b001100010010;
   4110: result <= 12'b001100010010;
   4111: result <= 12'b001100010010;
   4112: result <= 12'b001100010010;
   4113: result <= 12'b001100010010;
   4114: result <= 12'b001100010010;
   4115: result <= 12'b001100010011;
   4116: result <= 12'b001100010011;
   4117: result <= 12'b001100010011;
   4118: result <= 12'b001100010011;
   4119: result <= 12'b001100010011;
   4120: result <= 12'b001100010100;
   4121: result <= 12'b001100010100;
   4122: result <= 12'b001100010100;
   4123: result <= 12'b001100010100;
   4124: result <= 12'b001100010100;
   4125: result <= 12'b001100010100;
   4126: result <= 12'b001100010101;
   4127: result <= 12'b001100010101;
   4128: result <= 12'b001100010101;
   4129: result <= 12'b001100010101;
   4130: result <= 12'b001100010101;
   4131: result <= 12'b001100010110;
   4132: result <= 12'b001100010110;
   4133: result <= 12'b001100010110;
   4134: result <= 12'b001100010110;
   4135: result <= 12'b001100010110;
   4136: result <= 12'b001100010110;
   4137: result <= 12'b001100010111;
   4138: result <= 12'b001100010111;
   4139: result <= 12'b001100010111;
   4140: result <= 12'b001100010111;
   4141: result <= 12'b001100010111;
   4142: result <= 12'b001100011000;
   4143: result <= 12'b001100011000;
   4144: result <= 12'b001100011000;
   4145: result <= 12'b001100011000;
   4146: result <= 12'b001100011000;
   4147: result <= 12'b001100011000;
   4148: result <= 12'b001100011001;
   4149: result <= 12'b001100011001;
   4150: result <= 12'b001100011001;
   4151: result <= 12'b001100011001;
   4152: result <= 12'b001100011001;
   4153: result <= 12'b001100011010;
   4154: result <= 12'b001100011010;
   4155: result <= 12'b001100011010;
   4156: result <= 12'b001100011010;
   4157: result <= 12'b001100011010;
   4158: result <= 12'b001100011010;
   4159: result <= 12'b001100011011;
   4160: result <= 12'b001100011011;
   4161: result <= 12'b001100011011;
   4162: result <= 12'b001100011011;
   4163: result <= 12'b001100011011;
   4164: result <= 12'b001100011100;
   4165: result <= 12'b001100011100;
   4166: result <= 12'b001100011100;
   4167: result <= 12'b001100011100;
   4168: result <= 12'b001100011100;
   4169: result <= 12'b001100011100;
   4170: result <= 12'b001100011101;
   4171: result <= 12'b001100011101;
   4172: result <= 12'b001100011101;
   4173: result <= 12'b001100011101;
   4174: result <= 12'b001100011101;
   4175: result <= 12'b001100011110;
   4176: result <= 12'b001100011110;
   4177: result <= 12'b001100011110;
   4178: result <= 12'b001100011110;
   4179: result <= 12'b001100011110;
   4180: result <= 12'b001100011110;
   4181: result <= 12'b001100011111;
   4182: result <= 12'b001100011111;
   4183: result <= 12'b001100011111;
   4184: result <= 12'b001100011111;
   4185: result <= 12'b001100011111;
   4186: result <= 12'b001100100000;
   4187: result <= 12'b001100100000;
   4188: result <= 12'b001100100000;
   4189: result <= 12'b001100100000;
   4190: result <= 12'b001100100000;
   4191: result <= 12'b001100100000;
   4192: result <= 12'b001100100001;
   4193: result <= 12'b001100100001;
   4194: result <= 12'b001100100001;
   4195: result <= 12'b001100100001;
   4196: result <= 12'b001100100001;
   4197: result <= 12'b001100100010;
   4198: result <= 12'b001100100010;
   4199: result <= 12'b001100100010;
   4200: result <= 12'b001100100010;
   4201: result <= 12'b001100100010;
   4202: result <= 12'b001100100010;
   4203: result <= 12'b001100100011;
   4204: result <= 12'b001100100011;
   4205: result <= 12'b001100100011;
   4206: result <= 12'b001100100011;
   4207: result <= 12'b001100100011;
   4208: result <= 12'b001100100100;
   4209: result <= 12'b001100100100;
   4210: result <= 12'b001100100100;
   4211: result <= 12'b001100100100;
   4212: result <= 12'b001100100100;
   4213: result <= 12'b001100100100;
   4214: result <= 12'b001100100101;
   4215: result <= 12'b001100100101;
   4216: result <= 12'b001100100101;
   4217: result <= 12'b001100100101;
   4218: result <= 12'b001100100101;
   4219: result <= 12'b001100100101;
   4220: result <= 12'b001100100110;
   4221: result <= 12'b001100100110;
   4222: result <= 12'b001100100110;
   4223: result <= 12'b001100100110;
   4224: result <= 12'b001100100110;
   4225: result <= 12'b001100100111;
   4226: result <= 12'b001100100111;
   4227: result <= 12'b001100100111;
   4228: result <= 12'b001100100111;
   4229: result <= 12'b001100100111;
   4230: result <= 12'b001100100111;
   4231: result <= 12'b001100101000;
   4232: result <= 12'b001100101000;
   4233: result <= 12'b001100101000;
   4234: result <= 12'b001100101000;
   4235: result <= 12'b001100101000;
   4236: result <= 12'b001100101001;
   4237: result <= 12'b001100101001;
   4238: result <= 12'b001100101001;
   4239: result <= 12'b001100101001;
   4240: result <= 12'b001100101001;
   4241: result <= 12'b001100101001;
   4242: result <= 12'b001100101010;
   4243: result <= 12'b001100101010;
   4244: result <= 12'b001100101010;
   4245: result <= 12'b001100101010;
   4246: result <= 12'b001100101010;
   4247: result <= 12'b001100101011;
   4248: result <= 12'b001100101011;
   4249: result <= 12'b001100101011;
   4250: result <= 12'b001100101011;
   4251: result <= 12'b001100101011;
   4252: result <= 12'b001100101011;
   4253: result <= 12'b001100101100;
   4254: result <= 12'b001100101100;
   4255: result <= 12'b001100101100;
   4256: result <= 12'b001100101100;
   4257: result <= 12'b001100101100;
   4258: result <= 12'b001100101101;
   4259: result <= 12'b001100101101;
   4260: result <= 12'b001100101101;
   4261: result <= 12'b001100101101;
   4262: result <= 12'b001100101101;
   4263: result <= 12'b001100101101;
   4264: result <= 12'b001100101110;
   4265: result <= 12'b001100101110;
   4266: result <= 12'b001100101110;
   4267: result <= 12'b001100101110;
   4268: result <= 12'b001100101110;
   4269: result <= 12'b001100101111;
   4270: result <= 12'b001100101111;
   4271: result <= 12'b001100101111;
   4272: result <= 12'b001100101111;
   4273: result <= 12'b001100101111;
   4274: result <= 12'b001100101111;
   4275: result <= 12'b001100110000;
   4276: result <= 12'b001100110000;
   4277: result <= 12'b001100110000;
   4278: result <= 12'b001100110000;
   4279: result <= 12'b001100110000;
   4280: result <= 12'b001100110000;
   4281: result <= 12'b001100110001;
   4282: result <= 12'b001100110001;
   4283: result <= 12'b001100110001;
   4284: result <= 12'b001100110001;
   4285: result <= 12'b001100110001;
   4286: result <= 12'b001100110010;
   4287: result <= 12'b001100110010;
   4288: result <= 12'b001100110010;
   4289: result <= 12'b001100110010;
   4290: result <= 12'b001100110010;
   4291: result <= 12'b001100110010;
   4292: result <= 12'b001100110011;
   4293: result <= 12'b001100110011;
   4294: result <= 12'b001100110011;
   4295: result <= 12'b001100110011;
   4296: result <= 12'b001100110011;
   4297: result <= 12'b001100110100;
   4298: result <= 12'b001100110100;
   4299: result <= 12'b001100110100;
   4300: result <= 12'b001100110100;
   4301: result <= 12'b001100110100;
   4302: result <= 12'b001100110100;
   4303: result <= 12'b001100110101;
   4304: result <= 12'b001100110101;
   4305: result <= 12'b001100110101;
   4306: result <= 12'b001100110101;
   4307: result <= 12'b001100110101;
   4308: result <= 12'b001100110110;
   4309: result <= 12'b001100110110;
   4310: result <= 12'b001100110110;
   4311: result <= 12'b001100110110;
   4312: result <= 12'b001100110110;
   4313: result <= 12'b001100110110;
   4314: result <= 12'b001100110111;
   4315: result <= 12'b001100110111;
   4316: result <= 12'b001100110111;
   4317: result <= 12'b001100110111;
   4318: result <= 12'b001100110111;
   4319: result <= 12'b001100111000;
   4320: result <= 12'b001100111000;
   4321: result <= 12'b001100111000;
   4322: result <= 12'b001100111000;
   4323: result <= 12'b001100111000;
   4324: result <= 12'b001100111000;
   4325: result <= 12'b001100111001;
   4326: result <= 12'b001100111001;
   4327: result <= 12'b001100111001;
   4328: result <= 12'b001100111001;
   4329: result <= 12'b001100111001;
   4330: result <= 12'b001100111001;
   4331: result <= 12'b001100111010;
   4332: result <= 12'b001100111010;
   4333: result <= 12'b001100111010;
   4334: result <= 12'b001100111010;
   4335: result <= 12'b001100111010;
   4336: result <= 12'b001100111011;
   4337: result <= 12'b001100111011;
   4338: result <= 12'b001100111011;
   4339: result <= 12'b001100111011;
   4340: result <= 12'b001100111011;
   4341: result <= 12'b001100111011;
   4342: result <= 12'b001100111100;
   4343: result <= 12'b001100111100;
   4344: result <= 12'b001100111100;
   4345: result <= 12'b001100111100;
   4346: result <= 12'b001100111100;
   4347: result <= 12'b001100111101;
   4348: result <= 12'b001100111101;
   4349: result <= 12'b001100111101;
   4350: result <= 12'b001100111101;
   4351: result <= 12'b001100111101;
   4352: result <= 12'b001100111101;
   4353: result <= 12'b001100111110;
   4354: result <= 12'b001100111110;
   4355: result <= 12'b001100111110;
   4356: result <= 12'b001100111110;
   4357: result <= 12'b001100111110;
   4358: result <= 12'b001100111111;
   4359: result <= 12'b001100111111;
   4360: result <= 12'b001100111111;
   4361: result <= 12'b001100111111;
   4362: result <= 12'b001100111111;
   4363: result <= 12'b001100111111;
   4364: result <= 12'b001101000000;
   4365: result <= 12'b001101000000;
   4366: result <= 12'b001101000000;
   4367: result <= 12'b001101000000;
   4368: result <= 12'b001101000000;
   4369: result <= 12'b001101000000;
   4370: result <= 12'b001101000001;
   4371: result <= 12'b001101000001;
   4372: result <= 12'b001101000001;
   4373: result <= 12'b001101000001;
   4374: result <= 12'b001101000001;
   4375: result <= 12'b001101000010;
   4376: result <= 12'b001101000010;
   4377: result <= 12'b001101000010;
   4378: result <= 12'b001101000010;
   4379: result <= 12'b001101000010;
   4380: result <= 12'b001101000010;
   4381: result <= 12'b001101000011;
   4382: result <= 12'b001101000011;
   4383: result <= 12'b001101000011;
   4384: result <= 12'b001101000011;
   4385: result <= 12'b001101000011;
   4386: result <= 12'b001101000100;
   4387: result <= 12'b001101000100;
   4388: result <= 12'b001101000100;
   4389: result <= 12'b001101000100;
   4390: result <= 12'b001101000100;
   4391: result <= 12'b001101000100;
   4392: result <= 12'b001101000101;
   4393: result <= 12'b001101000101;
   4394: result <= 12'b001101000101;
   4395: result <= 12'b001101000101;
   4396: result <= 12'b001101000101;
   4397: result <= 12'b001101000110;
   4398: result <= 12'b001101000110;
   4399: result <= 12'b001101000110;
   4400: result <= 12'b001101000110;
   4401: result <= 12'b001101000110;
   4402: result <= 12'b001101000110;
   4403: result <= 12'b001101000111;
   4404: result <= 12'b001101000111;
   4405: result <= 12'b001101000111;
   4406: result <= 12'b001101000111;
   4407: result <= 12'b001101000111;
   4408: result <= 12'b001101000111;
   4409: result <= 12'b001101001000;
   4410: result <= 12'b001101001000;
   4411: result <= 12'b001101001000;
   4412: result <= 12'b001101001000;
   4413: result <= 12'b001101001000;
   4414: result <= 12'b001101001001;
   4415: result <= 12'b001101001001;
   4416: result <= 12'b001101001001;
   4417: result <= 12'b001101001001;
   4418: result <= 12'b001101001001;
   4419: result <= 12'b001101001001;
   4420: result <= 12'b001101001010;
   4421: result <= 12'b001101001010;
   4422: result <= 12'b001101001010;
   4423: result <= 12'b001101001010;
   4424: result <= 12'b001101001010;
   4425: result <= 12'b001101001011;
   4426: result <= 12'b001101001011;
   4427: result <= 12'b001101001011;
   4428: result <= 12'b001101001011;
   4429: result <= 12'b001101001011;
   4430: result <= 12'b001101001011;
   4431: result <= 12'b001101001100;
   4432: result <= 12'b001101001100;
   4433: result <= 12'b001101001100;
   4434: result <= 12'b001101001100;
   4435: result <= 12'b001101001100;
   4436: result <= 12'b001101001100;
   4437: result <= 12'b001101001101;
   4438: result <= 12'b001101001101;
   4439: result <= 12'b001101001101;
   4440: result <= 12'b001101001101;
   4441: result <= 12'b001101001101;
   4442: result <= 12'b001101001110;
   4443: result <= 12'b001101001110;
   4444: result <= 12'b001101001110;
   4445: result <= 12'b001101001110;
   4446: result <= 12'b001101001110;
   4447: result <= 12'b001101001110;
   4448: result <= 12'b001101001111;
   4449: result <= 12'b001101001111;
   4450: result <= 12'b001101001111;
   4451: result <= 12'b001101001111;
   4452: result <= 12'b001101001111;
   4453: result <= 12'b001101010000;
   4454: result <= 12'b001101010000;
   4455: result <= 12'b001101010000;
   4456: result <= 12'b001101010000;
   4457: result <= 12'b001101010000;
   4458: result <= 12'b001101010000;
   4459: result <= 12'b001101010001;
   4460: result <= 12'b001101010001;
   4461: result <= 12'b001101010001;
   4462: result <= 12'b001101010001;
   4463: result <= 12'b001101010001;
   4464: result <= 12'b001101010001;
   4465: result <= 12'b001101010010;
   4466: result <= 12'b001101010010;
   4467: result <= 12'b001101010010;
   4468: result <= 12'b001101010010;
   4469: result <= 12'b001101010010;
   4470: result <= 12'b001101010011;
   4471: result <= 12'b001101010011;
   4472: result <= 12'b001101010011;
   4473: result <= 12'b001101010011;
   4474: result <= 12'b001101010011;
   4475: result <= 12'b001101010011;
   4476: result <= 12'b001101010100;
   4477: result <= 12'b001101010100;
   4478: result <= 12'b001101010100;
   4479: result <= 12'b001101010100;
   4480: result <= 12'b001101010100;
   4481: result <= 12'b001101010101;
   4482: result <= 12'b001101010101;
   4483: result <= 12'b001101010101;
   4484: result <= 12'b001101010101;
   4485: result <= 12'b001101010101;
   4486: result <= 12'b001101010101;
   4487: result <= 12'b001101010110;
   4488: result <= 12'b001101010110;
   4489: result <= 12'b001101010110;
   4490: result <= 12'b001101010110;
   4491: result <= 12'b001101010110;
   4492: result <= 12'b001101010110;
   4493: result <= 12'b001101010111;
   4494: result <= 12'b001101010111;
   4495: result <= 12'b001101010111;
   4496: result <= 12'b001101010111;
   4497: result <= 12'b001101010111;
   4498: result <= 12'b001101011000;
   4499: result <= 12'b001101011000;
   4500: result <= 12'b001101011000;
   4501: result <= 12'b001101011000;
   4502: result <= 12'b001101011000;
   4503: result <= 12'b001101011000;
   4504: result <= 12'b001101011001;
   4505: result <= 12'b001101011001;
   4506: result <= 12'b001101011001;
   4507: result <= 12'b001101011001;
   4508: result <= 12'b001101011001;
   4509: result <= 12'b001101011010;
   4510: result <= 12'b001101011010;
   4511: result <= 12'b001101011010;
   4512: result <= 12'b001101011010;
   4513: result <= 12'b001101011010;
   4514: result <= 12'b001101011010;
   4515: result <= 12'b001101011011;
   4516: result <= 12'b001101011011;
   4517: result <= 12'b001101011011;
   4518: result <= 12'b001101011011;
   4519: result <= 12'b001101011011;
   4520: result <= 12'b001101011011;
   4521: result <= 12'b001101011100;
   4522: result <= 12'b001101011100;
   4523: result <= 12'b001101011100;
   4524: result <= 12'b001101011100;
   4525: result <= 12'b001101011100;
   4526: result <= 12'b001101011101;
   4527: result <= 12'b001101011101;
   4528: result <= 12'b001101011101;
   4529: result <= 12'b001101011101;
   4530: result <= 12'b001101011101;
   4531: result <= 12'b001101011101;
   4532: result <= 12'b001101011110;
   4533: result <= 12'b001101011110;
   4534: result <= 12'b001101011110;
   4535: result <= 12'b001101011110;
   4536: result <= 12'b001101011110;
   4537: result <= 12'b001101011111;
   4538: result <= 12'b001101011111;
   4539: result <= 12'b001101011111;
   4540: result <= 12'b001101011111;
   4541: result <= 12'b001101011111;
   4542: result <= 12'b001101011111;
   4543: result <= 12'b001101100000;
   4544: result <= 12'b001101100000;
   4545: result <= 12'b001101100000;
   4546: result <= 12'b001101100000;
   4547: result <= 12'b001101100000;
   4548: result <= 12'b001101100000;
   4549: result <= 12'b001101100001;
   4550: result <= 12'b001101100001;
   4551: result <= 12'b001101100001;
   4552: result <= 12'b001101100001;
   4553: result <= 12'b001101100001;
   4554: result <= 12'b001101100010;
   4555: result <= 12'b001101100010;
   4556: result <= 12'b001101100010;
   4557: result <= 12'b001101100010;
   4558: result <= 12'b001101100010;
   4559: result <= 12'b001101100010;
   4560: result <= 12'b001101100011;
   4561: result <= 12'b001101100011;
   4562: result <= 12'b001101100011;
   4563: result <= 12'b001101100011;
   4564: result <= 12'b001101100011;
   4565: result <= 12'b001101100011;
   4566: result <= 12'b001101100100;
   4567: result <= 12'b001101100100;
   4568: result <= 12'b001101100100;
   4569: result <= 12'b001101100100;
   4570: result <= 12'b001101100100;
   4571: result <= 12'b001101100101;
   4572: result <= 12'b001101100101;
   4573: result <= 12'b001101100101;
   4574: result <= 12'b001101100101;
   4575: result <= 12'b001101100101;
   4576: result <= 12'b001101100101;
   4577: result <= 12'b001101100110;
   4578: result <= 12'b001101100110;
   4579: result <= 12'b001101100110;
   4580: result <= 12'b001101100110;
   4581: result <= 12'b001101100110;
   4582: result <= 12'b001101100111;
   4583: result <= 12'b001101100111;
   4584: result <= 12'b001101100111;
   4585: result <= 12'b001101100111;
   4586: result <= 12'b001101100111;
   4587: result <= 12'b001101100111;
   4588: result <= 12'b001101101000;
   4589: result <= 12'b001101101000;
   4590: result <= 12'b001101101000;
   4591: result <= 12'b001101101000;
   4592: result <= 12'b001101101000;
   4593: result <= 12'b001101101000;
   4594: result <= 12'b001101101001;
   4595: result <= 12'b001101101001;
   4596: result <= 12'b001101101001;
   4597: result <= 12'b001101101001;
   4598: result <= 12'b001101101001;
   4599: result <= 12'b001101101010;
   4600: result <= 12'b001101101010;
   4601: result <= 12'b001101101010;
   4602: result <= 12'b001101101010;
   4603: result <= 12'b001101101010;
   4604: result <= 12'b001101101010;
   4605: result <= 12'b001101101011;
   4606: result <= 12'b001101101011;
   4607: result <= 12'b001101101011;
   4608: result <= 12'b001101101011;
   4609: result <= 12'b001101101011;
   4610: result <= 12'b001101101011;
   4611: result <= 12'b001101101100;
   4612: result <= 12'b001101101100;
   4613: result <= 12'b001101101100;
   4614: result <= 12'b001101101100;
   4615: result <= 12'b001101101100;
   4616: result <= 12'b001101101101;
   4617: result <= 12'b001101101101;
   4618: result <= 12'b001101101101;
   4619: result <= 12'b001101101101;
   4620: result <= 12'b001101101101;
   4621: result <= 12'b001101101101;
   4622: result <= 12'b001101101110;
   4623: result <= 12'b001101101110;
   4624: result <= 12'b001101101110;
   4625: result <= 12'b001101101110;
   4626: result <= 12'b001101101110;
   4627: result <= 12'b001101101111;
   4628: result <= 12'b001101101111;
   4629: result <= 12'b001101101111;
   4630: result <= 12'b001101101111;
   4631: result <= 12'b001101101111;
   4632: result <= 12'b001101101111;
   4633: result <= 12'b001101110000;
   4634: result <= 12'b001101110000;
   4635: result <= 12'b001101110000;
   4636: result <= 12'b001101110000;
   4637: result <= 12'b001101110000;
   4638: result <= 12'b001101110000;
   4639: result <= 12'b001101110001;
   4640: result <= 12'b001101110001;
   4641: result <= 12'b001101110001;
   4642: result <= 12'b001101110001;
   4643: result <= 12'b001101110001;
   4644: result <= 12'b001101110010;
   4645: result <= 12'b001101110010;
   4646: result <= 12'b001101110010;
   4647: result <= 12'b001101110010;
   4648: result <= 12'b001101110010;
   4649: result <= 12'b001101110010;
   4650: result <= 12'b001101110011;
   4651: result <= 12'b001101110011;
   4652: result <= 12'b001101110011;
   4653: result <= 12'b001101110011;
   4654: result <= 12'b001101110011;
   4655: result <= 12'b001101110011;
   4656: result <= 12'b001101110100;
   4657: result <= 12'b001101110100;
   4658: result <= 12'b001101110100;
   4659: result <= 12'b001101110100;
   4660: result <= 12'b001101110100;
   4661: result <= 12'b001101110101;
   4662: result <= 12'b001101110101;
   4663: result <= 12'b001101110101;
   4664: result <= 12'b001101110101;
   4665: result <= 12'b001101110101;
   4666: result <= 12'b001101110101;
   4667: result <= 12'b001101110110;
   4668: result <= 12'b001101110110;
   4669: result <= 12'b001101110110;
   4670: result <= 12'b001101110110;
   4671: result <= 12'b001101110110;
   4672: result <= 12'b001101110110;
   4673: result <= 12'b001101110111;
   4674: result <= 12'b001101110111;
   4675: result <= 12'b001101110111;
   4676: result <= 12'b001101110111;
   4677: result <= 12'b001101110111;
   4678: result <= 12'b001101111000;
   4679: result <= 12'b001101111000;
   4680: result <= 12'b001101111000;
   4681: result <= 12'b001101111000;
   4682: result <= 12'b001101111000;
   4683: result <= 12'b001101111000;
   4684: result <= 12'b001101111001;
   4685: result <= 12'b001101111001;
   4686: result <= 12'b001101111001;
   4687: result <= 12'b001101111001;
   4688: result <= 12'b001101111001;
   4689: result <= 12'b001101111001;
   4690: result <= 12'b001101111010;
   4691: result <= 12'b001101111010;
   4692: result <= 12'b001101111010;
   4693: result <= 12'b001101111010;
   4694: result <= 12'b001101111010;
   4695: result <= 12'b001101111011;
   4696: result <= 12'b001101111011;
   4697: result <= 12'b001101111011;
   4698: result <= 12'b001101111011;
   4699: result <= 12'b001101111011;
   4700: result <= 12'b001101111011;
   4701: result <= 12'b001101111100;
   4702: result <= 12'b001101111100;
   4703: result <= 12'b001101111100;
   4704: result <= 12'b001101111100;
   4705: result <= 12'b001101111100;
   4706: result <= 12'b001101111100;
   4707: result <= 12'b001101111101;
   4708: result <= 12'b001101111101;
   4709: result <= 12'b001101111101;
   4710: result <= 12'b001101111101;
   4711: result <= 12'b001101111101;
   4712: result <= 12'b001101111110;
   4713: result <= 12'b001101111110;
   4714: result <= 12'b001101111110;
   4715: result <= 12'b001101111110;
   4716: result <= 12'b001101111110;
   4717: result <= 12'b001101111110;
   4718: result <= 12'b001101111111;
   4719: result <= 12'b001101111111;
   4720: result <= 12'b001101111111;
   4721: result <= 12'b001101111111;
   4722: result <= 12'b001101111111;
   4723: result <= 12'b001101111111;
   4724: result <= 12'b001110000000;
   4725: result <= 12'b001110000000;
   4726: result <= 12'b001110000000;
   4727: result <= 12'b001110000000;
   4728: result <= 12'b001110000000;
   4729: result <= 12'b001110000001;
   4730: result <= 12'b001110000001;
   4731: result <= 12'b001110000001;
   4732: result <= 12'b001110000001;
   4733: result <= 12'b001110000001;
   4734: result <= 12'b001110000001;
   4735: result <= 12'b001110000010;
   4736: result <= 12'b001110000010;
   4737: result <= 12'b001110000010;
   4738: result <= 12'b001110000010;
   4739: result <= 12'b001110000010;
   4740: result <= 12'b001110000010;
   4741: result <= 12'b001110000011;
   4742: result <= 12'b001110000011;
   4743: result <= 12'b001110000011;
   4744: result <= 12'b001110000011;
   4745: result <= 12'b001110000011;
   4746: result <= 12'b001110000100;
   4747: result <= 12'b001110000100;
   4748: result <= 12'b001110000100;
   4749: result <= 12'b001110000100;
   4750: result <= 12'b001110000100;
   4751: result <= 12'b001110000100;
   4752: result <= 12'b001110000101;
   4753: result <= 12'b001110000101;
   4754: result <= 12'b001110000101;
   4755: result <= 12'b001110000101;
   4756: result <= 12'b001110000101;
   4757: result <= 12'b001110000101;
   4758: result <= 12'b001110000110;
   4759: result <= 12'b001110000110;
   4760: result <= 12'b001110000110;
   4761: result <= 12'b001110000110;
   4762: result <= 12'b001110000110;
   4763: result <= 12'b001110000111;
   4764: result <= 12'b001110000111;
   4765: result <= 12'b001110000111;
   4766: result <= 12'b001110000111;
   4767: result <= 12'b001110000111;
   4768: result <= 12'b001110000111;
   4769: result <= 12'b001110001000;
   4770: result <= 12'b001110001000;
   4771: result <= 12'b001110001000;
   4772: result <= 12'b001110001000;
   4773: result <= 12'b001110001000;
   4774: result <= 12'b001110001000;
   4775: result <= 12'b001110001001;
   4776: result <= 12'b001110001001;
   4777: result <= 12'b001110001001;
   4778: result <= 12'b001110001001;
   4779: result <= 12'b001110001001;
   4780: result <= 12'b001110001010;
   4781: result <= 12'b001110001010;
   4782: result <= 12'b001110001010;
   4783: result <= 12'b001110001010;
   4784: result <= 12'b001110001010;
   4785: result <= 12'b001110001010;
   4786: result <= 12'b001110001011;
   4787: result <= 12'b001110001011;
   4788: result <= 12'b001110001011;
   4789: result <= 12'b001110001011;
   4790: result <= 12'b001110001011;
   4791: result <= 12'b001110001011;
   4792: result <= 12'b001110001100;
   4793: result <= 12'b001110001100;
   4794: result <= 12'b001110001100;
   4795: result <= 12'b001110001100;
   4796: result <= 12'b001110001100;
   4797: result <= 12'b001110001101;
   4798: result <= 12'b001110001101;
   4799: result <= 12'b001110001101;
   4800: result <= 12'b001110001101;
   4801: result <= 12'b001110001101;
   4802: result <= 12'b001110001101;
   4803: result <= 12'b001110001110;
   4804: result <= 12'b001110001110;
   4805: result <= 12'b001110001110;
   4806: result <= 12'b001110001110;
   4807: result <= 12'b001110001110;
   4808: result <= 12'b001110001110;
   4809: result <= 12'b001110001111;
   4810: result <= 12'b001110001111;
   4811: result <= 12'b001110001111;
   4812: result <= 12'b001110001111;
   4813: result <= 12'b001110001111;
   4814: result <= 12'b001110010000;
   4815: result <= 12'b001110010000;
   4816: result <= 12'b001110010000;
   4817: result <= 12'b001110010000;
   4818: result <= 12'b001110010000;
   4819: result <= 12'b001110010000;
   4820: result <= 12'b001110010001;
   4821: result <= 12'b001110010001;
   4822: result <= 12'b001110010001;
   4823: result <= 12'b001110010001;
   4824: result <= 12'b001110010001;
   4825: result <= 12'b001110010001;
   4826: result <= 12'b001110010010;
   4827: result <= 12'b001110010010;
   4828: result <= 12'b001110010010;
   4829: result <= 12'b001110010010;
   4830: result <= 12'b001110010010;
   4831: result <= 12'b001110010011;
   4832: result <= 12'b001110010011;
   4833: result <= 12'b001110010011;
   4834: result <= 12'b001110010011;
   4835: result <= 12'b001110010011;
   4836: result <= 12'b001110010011;
   4837: result <= 12'b001110010100;
   4838: result <= 12'b001110010100;
   4839: result <= 12'b001110010100;
   4840: result <= 12'b001110010100;
   4841: result <= 12'b001110010100;
   4842: result <= 12'b001110010100;
   4843: result <= 12'b001110010101;
   4844: result <= 12'b001110010101;
   4845: result <= 12'b001110010101;
   4846: result <= 12'b001110010101;
   4847: result <= 12'b001110010101;
   4848: result <= 12'b001110010101;
   4849: result <= 12'b001110010110;
   4850: result <= 12'b001110010110;
   4851: result <= 12'b001110010110;
   4852: result <= 12'b001110010110;
   4853: result <= 12'b001110010110;
   4854: result <= 12'b001110010111;
   4855: result <= 12'b001110010111;
   4856: result <= 12'b001110010111;
   4857: result <= 12'b001110010111;
   4858: result <= 12'b001110010111;
   4859: result <= 12'b001110010111;
   4860: result <= 12'b001110011000;
   4861: result <= 12'b001110011000;
   4862: result <= 12'b001110011000;
   4863: result <= 12'b001110011000;
   4864: result <= 12'b001110011000;
   4865: result <= 12'b001110011000;
   4866: result <= 12'b001110011001;
   4867: result <= 12'b001110011001;
   4868: result <= 12'b001110011001;
   4869: result <= 12'b001110011001;
   4870: result <= 12'b001110011001;
   4871: result <= 12'b001110011010;
   4872: result <= 12'b001110011010;
   4873: result <= 12'b001110011010;
   4874: result <= 12'b001110011010;
   4875: result <= 12'b001110011010;
   4876: result <= 12'b001110011010;
   4877: result <= 12'b001110011011;
   4878: result <= 12'b001110011011;
   4879: result <= 12'b001110011011;
   4880: result <= 12'b001110011011;
   4881: result <= 12'b001110011011;
   4882: result <= 12'b001110011011;
   4883: result <= 12'b001110011100;
   4884: result <= 12'b001110011100;
   4885: result <= 12'b001110011100;
   4886: result <= 12'b001110011100;
   4887: result <= 12'b001110011100;
   4888: result <= 12'b001110011101;
   4889: result <= 12'b001110011101;
   4890: result <= 12'b001110011101;
   4891: result <= 12'b001110011101;
   4892: result <= 12'b001110011101;
   4893: result <= 12'b001110011101;
   4894: result <= 12'b001110011110;
   4895: result <= 12'b001110011110;
   4896: result <= 12'b001110011110;
   4897: result <= 12'b001110011110;
   4898: result <= 12'b001110011110;
   4899: result <= 12'b001110011110;
   4900: result <= 12'b001110011111;
   4901: result <= 12'b001110011111;
   4902: result <= 12'b001110011111;
   4903: result <= 12'b001110011111;
   4904: result <= 12'b001110011111;
   4905: result <= 12'b001110011111;
   4906: result <= 12'b001110100000;
   4907: result <= 12'b001110100000;
   4908: result <= 12'b001110100000;
   4909: result <= 12'b001110100000;
   4910: result <= 12'b001110100000;
   4911: result <= 12'b001110100001;
   4912: result <= 12'b001110100001;
   4913: result <= 12'b001110100001;
   4914: result <= 12'b001110100001;
   4915: result <= 12'b001110100001;
   4916: result <= 12'b001110100001;
   4917: result <= 12'b001110100010;
   4918: result <= 12'b001110100010;
   4919: result <= 12'b001110100010;
   4920: result <= 12'b001110100010;
   4921: result <= 12'b001110100010;
   4922: result <= 12'b001110100010;
   4923: result <= 12'b001110100011;
   4924: result <= 12'b001110100011;
   4925: result <= 12'b001110100011;
   4926: result <= 12'b001110100011;
   4927: result <= 12'b001110100011;
   4928: result <= 12'b001110100100;
   4929: result <= 12'b001110100100;
   4930: result <= 12'b001110100100;
   4931: result <= 12'b001110100100;
   4932: result <= 12'b001110100100;
   4933: result <= 12'b001110100100;
   4934: result <= 12'b001110100101;
   4935: result <= 12'b001110100101;
   4936: result <= 12'b001110100101;
   4937: result <= 12'b001110100101;
   4938: result <= 12'b001110100101;
   4939: result <= 12'b001110100101;
   4940: result <= 12'b001110100110;
   4941: result <= 12'b001110100110;
   4942: result <= 12'b001110100110;
   4943: result <= 12'b001110100110;
   4944: result <= 12'b001110100110;
   4945: result <= 12'b001110100110;
   4946: result <= 12'b001110100111;
   4947: result <= 12'b001110100111;
   4948: result <= 12'b001110100111;
   4949: result <= 12'b001110100111;
   4950: result <= 12'b001110100111;
   4951: result <= 12'b001110101000;
   4952: result <= 12'b001110101000;
   4953: result <= 12'b001110101000;
   4954: result <= 12'b001110101000;
   4955: result <= 12'b001110101000;
   4956: result <= 12'b001110101000;
   4957: result <= 12'b001110101001;
   4958: result <= 12'b001110101001;
   4959: result <= 12'b001110101001;
   4960: result <= 12'b001110101001;
   4961: result <= 12'b001110101001;
   4962: result <= 12'b001110101001;
   4963: result <= 12'b001110101010;
   4964: result <= 12'b001110101010;
   4965: result <= 12'b001110101010;
   4966: result <= 12'b001110101010;
   4967: result <= 12'b001110101010;
   4968: result <= 12'b001110101010;
   4969: result <= 12'b001110101011;
   4970: result <= 12'b001110101011;
   4971: result <= 12'b001110101011;
   4972: result <= 12'b001110101011;
   4973: result <= 12'b001110101011;
   4974: result <= 12'b001110101100;
   4975: result <= 12'b001110101100;
   4976: result <= 12'b001110101100;
   4977: result <= 12'b001110101100;
   4978: result <= 12'b001110101100;
   4979: result <= 12'b001110101100;
   4980: result <= 12'b001110101101;
   4981: result <= 12'b001110101101;
   4982: result <= 12'b001110101101;
   4983: result <= 12'b001110101101;
   4984: result <= 12'b001110101101;
   4985: result <= 12'b001110101101;
   4986: result <= 12'b001110101110;
   4987: result <= 12'b001110101110;
   4988: result <= 12'b001110101110;
   4989: result <= 12'b001110101110;
   4990: result <= 12'b001110101110;
   4991: result <= 12'b001110101111;
   4992: result <= 12'b001110101111;
   4993: result <= 12'b001110101111;
   4994: result <= 12'b001110101111;
   4995: result <= 12'b001110101111;
   4996: result <= 12'b001110101111;
   4997: result <= 12'b001110110000;
   4998: result <= 12'b001110110000;
   4999: result <= 12'b001110110000;
   5000: result <= 12'b001110110000;
   5001: result <= 12'b001110110000;
   5002: result <= 12'b001110110000;
   5003: result <= 12'b001110110001;
   5004: result <= 12'b001110110001;
   5005: result <= 12'b001110110001;
   5006: result <= 12'b001110110001;
   5007: result <= 12'b001110110001;
   5008: result <= 12'b001110110001;
   5009: result <= 12'b001110110010;
   5010: result <= 12'b001110110010;
   5011: result <= 12'b001110110010;
   5012: result <= 12'b001110110010;
   5013: result <= 12'b001110110010;
   5014: result <= 12'b001110110011;
   5015: result <= 12'b001110110011;
   5016: result <= 12'b001110110011;
   5017: result <= 12'b001110110011;
   5018: result <= 12'b001110110011;
   5019: result <= 12'b001110110011;
   5020: result <= 12'b001110110100;
   5021: result <= 12'b001110110100;
   5022: result <= 12'b001110110100;
   5023: result <= 12'b001110110100;
   5024: result <= 12'b001110110100;
   5025: result <= 12'b001110110100;
   5026: result <= 12'b001110110101;
   5027: result <= 12'b001110110101;
   5028: result <= 12'b001110110101;
   5029: result <= 12'b001110110101;
   5030: result <= 12'b001110110101;
   5031: result <= 12'b001110110101;
   5032: result <= 12'b001110110110;
   5033: result <= 12'b001110110110;
   5034: result <= 12'b001110110110;
   5035: result <= 12'b001110110110;
   5036: result <= 12'b001110110110;
   5037: result <= 12'b001110110111;
   5038: result <= 12'b001110110111;
   5039: result <= 12'b001110110111;
   5040: result <= 12'b001110110111;
   5041: result <= 12'b001110110111;
   5042: result <= 12'b001110110111;
   5043: result <= 12'b001110111000;
   5044: result <= 12'b001110111000;
   5045: result <= 12'b001110111000;
   5046: result <= 12'b001110111000;
   5047: result <= 12'b001110111000;
   5048: result <= 12'b001110111000;
   5049: result <= 12'b001110111001;
   5050: result <= 12'b001110111001;
   5051: result <= 12'b001110111001;
   5052: result <= 12'b001110111001;
   5053: result <= 12'b001110111001;
   5054: result <= 12'b001110111001;
   5055: result <= 12'b001110111010;
   5056: result <= 12'b001110111010;
   5057: result <= 12'b001110111010;
   5058: result <= 12'b001110111010;
   5059: result <= 12'b001110111010;
   5060: result <= 12'b001110111011;
   5061: result <= 12'b001110111011;
   5062: result <= 12'b001110111011;
   5063: result <= 12'b001110111011;
   5064: result <= 12'b001110111011;
   5065: result <= 12'b001110111011;
   5066: result <= 12'b001110111100;
   5067: result <= 12'b001110111100;
   5068: result <= 12'b001110111100;
   5069: result <= 12'b001110111100;
   5070: result <= 12'b001110111100;
   5071: result <= 12'b001110111100;
   5072: result <= 12'b001110111101;
   5073: result <= 12'b001110111101;
   5074: result <= 12'b001110111101;
   5075: result <= 12'b001110111101;
   5076: result <= 12'b001110111101;
   5077: result <= 12'b001110111101;
   5078: result <= 12'b001110111110;
   5079: result <= 12'b001110111110;
   5080: result <= 12'b001110111110;
   5081: result <= 12'b001110111110;
   5082: result <= 12'b001110111110;
   5083: result <= 12'b001110111111;
   5084: result <= 12'b001110111111;
   5085: result <= 12'b001110111111;
   5086: result <= 12'b001110111111;
   5087: result <= 12'b001110111111;
   5088: result <= 12'b001110111111;
   5089: result <= 12'b001111000000;
   5090: result <= 12'b001111000000;
   5091: result <= 12'b001111000000;
   5092: result <= 12'b001111000000;
   5093: result <= 12'b001111000000;
   5094: result <= 12'b001111000000;
   5095: result <= 12'b001111000001;
   5096: result <= 12'b001111000001;
   5097: result <= 12'b001111000001;
   5098: result <= 12'b001111000001;
   5099: result <= 12'b001111000001;
   5100: result <= 12'b001111000001;
   5101: result <= 12'b001111000010;
   5102: result <= 12'b001111000010;
   5103: result <= 12'b001111000010;
   5104: result <= 12'b001111000010;
   5105: result <= 12'b001111000010;
   5106: result <= 12'b001111000010;
   5107: result <= 12'b001111000011;
   5108: result <= 12'b001111000011;
   5109: result <= 12'b001111000011;
   5110: result <= 12'b001111000011;
   5111: result <= 12'b001111000011;
   5112: result <= 12'b001111000100;
   5113: result <= 12'b001111000100;
   5114: result <= 12'b001111000100;
   5115: result <= 12'b001111000100;
   5116: result <= 12'b001111000100;
   5117: result <= 12'b001111000100;
   5118: result <= 12'b001111000101;
   5119: result <= 12'b001111000101;
   5120: result <= 12'b001111000101;
   5121: result <= 12'b001111000101;
   5122: result <= 12'b001111000101;
   5123: result <= 12'b001111000101;
   5124: result <= 12'b001111000110;
   5125: result <= 12'b001111000110;
   5126: result <= 12'b001111000110;
   5127: result <= 12'b001111000110;
   5128: result <= 12'b001111000110;
   5129: result <= 12'b001111000110;
   5130: result <= 12'b001111000111;
   5131: result <= 12'b001111000111;
   5132: result <= 12'b001111000111;
   5133: result <= 12'b001111000111;
   5134: result <= 12'b001111000111;
   5135: result <= 12'b001111001000;
   5136: result <= 12'b001111001000;
   5137: result <= 12'b001111001000;
   5138: result <= 12'b001111001000;
   5139: result <= 12'b001111001000;
   5140: result <= 12'b001111001000;
   5141: result <= 12'b001111001001;
   5142: result <= 12'b001111001001;
   5143: result <= 12'b001111001001;
   5144: result <= 12'b001111001001;
   5145: result <= 12'b001111001001;
   5146: result <= 12'b001111001001;
   5147: result <= 12'b001111001010;
   5148: result <= 12'b001111001010;
   5149: result <= 12'b001111001010;
   5150: result <= 12'b001111001010;
   5151: result <= 12'b001111001010;
   5152: result <= 12'b001111001010;
   5153: result <= 12'b001111001011;
   5154: result <= 12'b001111001011;
   5155: result <= 12'b001111001011;
   5156: result <= 12'b001111001011;
   5157: result <= 12'b001111001011;
   5158: result <= 12'b001111001011;
   5159: result <= 12'b001111001100;
   5160: result <= 12'b001111001100;
   5161: result <= 12'b001111001100;
   5162: result <= 12'b001111001100;
   5163: result <= 12'b001111001100;
   5164: result <= 12'b001111001101;
   5165: result <= 12'b001111001101;
   5166: result <= 12'b001111001101;
   5167: result <= 12'b001111001101;
   5168: result <= 12'b001111001101;
   5169: result <= 12'b001111001101;
   5170: result <= 12'b001111001110;
   5171: result <= 12'b001111001110;
   5172: result <= 12'b001111001110;
   5173: result <= 12'b001111001110;
   5174: result <= 12'b001111001110;
   5175: result <= 12'b001111001110;
   5176: result <= 12'b001111001111;
   5177: result <= 12'b001111001111;
   5178: result <= 12'b001111001111;
   5179: result <= 12'b001111001111;
   5180: result <= 12'b001111001111;
   5181: result <= 12'b001111001111;
   5182: result <= 12'b001111010000;
   5183: result <= 12'b001111010000;
   5184: result <= 12'b001111010000;
   5185: result <= 12'b001111010000;
   5186: result <= 12'b001111010000;
   5187: result <= 12'b001111010001;
   5188: result <= 12'b001111010001;
   5189: result <= 12'b001111010001;
   5190: result <= 12'b001111010001;
   5191: result <= 12'b001111010001;
   5192: result <= 12'b001111010001;
   5193: result <= 12'b001111010010;
   5194: result <= 12'b001111010010;
   5195: result <= 12'b001111010010;
   5196: result <= 12'b001111010010;
   5197: result <= 12'b001111010010;
   5198: result <= 12'b001111010010;
   5199: result <= 12'b001111010011;
   5200: result <= 12'b001111010011;
   5201: result <= 12'b001111010011;
   5202: result <= 12'b001111010011;
   5203: result <= 12'b001111010011;
   5204: result <= 12'b001111010011;
   5205: result <= 12'b001111010100;
   5206: result <= 12'b001111010100;
   5207: result <= 12'b001111010100;
   5208: result <= 12'b001111010100;
   5209: result <= 12'b001111010100;
   5210: result <= 12'b001111010100;
   5211: result <= 12'b001111010101;
   5212: result <= 12'b001111010101;
   5213: result <= 12'b001111010101;
   5214: result <= 12'b001111010101;
   5215: result <= 12'b001111010101;
   5216: result <= 12'b001111010110;
   5217: result <= 12'b001111010110;
   5218: result <= 12'b001111010110;
   5219: result <= 12'b001111010110;
   5220: result <= 12'b001111010110;
   5221: result <= 12'b001111010110;
   5222: result <= 12'b001111010111;
   5223: result <= 12'b001111010111;
   5224: result <= 12'b001111010111;
   5225: result <= 12'b001111010111;
   5226: result <= 12'b001111010111;
   5227: result <= 12'b001111010111;
   5228: result <= 12'b001111011000;
   5229: result <= 12'b001111011000;
   5230: result <= 12'b001111011000;
   5231: result <= 12'b001111011000;
   5232: result <= 12'b001111011000;
   5233: result <= 12'b001111011000;
   5234: result <= 12'b001111011001;
   5235: result <= 12'b001111011001;
   5236: result <= 12'b001111011001;
   5237: result <= 12'b001111011001;
   5238: result <= 12'b001111011001;
   5239: result <= 12'b001111011001;
   5240: result <= 12'b001111011010;
   5241: result <= 12'b001111011010;
   5242: result <= 12'b001111011010;
   5243: result <= 12'b001111011010;
   5244: result <= 12'b001111011010;
   5245: result <= 12'b001111011010;
   5246: result <= 12'b001111011011;
   5247: result <= 12'b001111011011;
   5248: result <= 12'b001111011011;
   5249: result <= 12'b001111011011;
   5250: result <= 12'b001111011011;
   5251: result <= 12'b001111011100;
   5252: result <= 12'b001111011100;
   5253: result <= 12'b001111011100;
   5254: result <= 12'b001111011100;
   5255: result <= 12'b001111011100;
   5256: result <= 12'b001111011100;
   5257: result <= 12'b001111011101;
   5258: result <= 12'b001111011101;
   5259: result <= 12'b001111011101;
   5260: result <= 12'b001111011101;
   5261: result <= 12'b001111011101;
   5262: result <= 12'b001111011101;
   5263: result <= 12'b001111011110;
   5264: result <= 12'b001111011110;
   5265: result <= 12'b001111011110;
   5266: result <= 12'b001111011110;
   5267: result <= 12'b001111011110;
   5268: result <= 12'b001111011110;
   5269: result <= 12'b001111011111;
   5270: result <= 12'b001111011111;
   5271: result <= 12'b001111011111;
   5272: result <= 12'b001111011111;
   5273: result <= 12'b001111011111;
   5274: result <= 12'b001111011111;
   5275: result <= 12'b001111100000;
   5276: result <= 12'b001111100000;
   5277: result <= 12'b001111100000;
   5278: result <= 12'b001111100000;
   5279: result <= 12'b001111100000;
   5280: result <= 12'b001111100001;
   5281: result <= 12'b001111100001;
   5282: result <= 12'b001111100001;
   5283: result <= 12'b001111100001;
   5284: result <= 12'b001111100001;
   5285: result <= 12'b001111100001;
   5286: result <= 12'b001111100010;
   5287: result <= 12'b001111100010;
   5288: result <= 12'b001111100010;
   5289: result <= 12'b001111100010;
   5290: result <= 12'b001111100010;
   5291: result <= 12'b001111100010;
   5292: result <= 12'b001111100011;
   5293: result <= 12'b001111100011;
   5294: result <= 12'b001111100011;
   5295: result <= 12'b001111100011;
   5296: result <= 12'b001111100011;
   5297: result <= 12'b001111100011;
   5298: result <= 12'b001111100100;
   5299: result <= 12'b001111100100;
   5300: result <= 12'b001111100100;
   5301: result <= 12'b001111100100;
   5302: result <= 12'b001111100100;
   5303: result <= 12'b001111100100;
   5304: result <= 12'b001111100101;
   5305: result <= 12'b001111100101;
   5306: result <= 12'b001111100101;
   5307: result <= 12'b001111100101;
   5308: result <= 12'b001111100101;
   5309: result <= 12'b001111100101;
   5310: result <= 12'b001111100110;
   5311: result <= 12'b001111100110;
   5312: result <= 12'b001111100110;
   5313: result <= 12'b001111100110;
   5314: result <= 12'b001111100110;
   5315: result <= 12'b001111100111;
   5316: result <= 12'b001111100111;
   5317: result <= 12'b001111100111;
   5318: result <= 12'b001111100111;
   5319: result <= 12'b001111100111;
   5320: result <= 12'b001111100111;
   5321: result <= 12'b001111101000;
   5322: result <= 12'b001111101000;
   5323: result <= 12'b001111101000;
   5324: result <= 12'b001111101000;
   5325: result <= 12'b001111101000;
   5326: result <= 12'b001111101000;
   5327: result <= 12'b001111101001;
   5328: result <= 12'b001111101001;
   5329: result <= 12'b001111101001;
   5330: result <= 12'b001111101001;
   5331: result <= 12'b001111101001;
   5332: result <= 12'b001111101001;
   5333: result <= 12'b001111101010;
   5334: result <= 12'b001111101010;
   5335: result <= 12'b001111101010;
   5336: result <= 12'b001111101010;
   5337: result <= 12'b001111101010;
   5338: result <= 12'b001111101010;
   5339: result <= 12'b001111101011;
   5340: result <= 12'b001111101011;
   5341: result <= 12'b001111101011;
   5342: result <= 12'b001111101011;
   5343: result <= 12'b001111101011;
   5344: result <= 12'b001111101011;
   5345: result <= 12'b001111101100;
   5346: result <= 12'b001111101100;
   5347: result <= 12'b001111101100;
   5348: result <= 12'b001111101100;
   5349: result <= 12'b001111101100;
   5350: result <= 12'b001111101101;
   5351: result <= 12'b001111101101;
   5352: result <= 12'b001111101101;
   5353: result <= 12'b001111101101;
   5354: result <= 12'b001111101101;
   5355: result <= 12'b001111101101;
   5356: result <= 12'b001111101110;
   5357: result <= 12'b001111101110;
   5358: result <= 12'b001111101110;
   5359: result <= 12'b001111101110;
   5360: result <= 12'b001111101110;
   5361: result <= 12'b001111101110;
   5362: result <= 12'b001111101111;
   5363: result <= 12'b001111101111;
   5364: result <= 12'b001111101111;
   5365: result <= 12'b001111101111;
   5366: result <= 12'b001111101111;
   5367: result <= 12'b001111101111;
   5368: result <= 12'b001111110000;
   5369: result <= 12'b001111110000;
   5370: result <= 12'b001111110000;
   5371: result <= 12'b001111110000;
   5372: result <= 12'b001111110000;
   5373: result <= 12'b001111110000;
   5374: result <= 12'b001111110001;
   5375: result <= 12'b001111110001;
   5376: result <= 12'b001111110001;
   5377: result <= 12'b001111110001;
   5378: result <= 12'b001111110001;
   5379: result <= 12'b001111110001;
   5380: result <= 12'b001111110010;
   5381: result <= 12'b001111110010;
   5382: result <= 12'b001111110010;
   5383: result <= 12'b001111110010;
   5384: result <= 12'b001111110010;
   5385: result <= 12'b001111110010;
   5386: result <= 12'b001111110011;
   5387: result <= 12'b001111110011;
   5388: result <= 12'b001111110011;
   5389: result <= 12'b001111110011;
   5390: result <= 12'b001111110011;
   5391: result <= 12'b001111110100;
   5392: result <= 12'b001111110100;
   5393: result <= 12'b001111110100;
   5394: result <= 12'b001111110100;
   5395: result <= 12'b001111110100;
   5396: result <= 12'b001111110100;
   5397: result <= 12'b001111110101;
   5398: result <= 12'b001111110101;
   5399: result <= 12'b001111110101;
   5400: result <= 12'b001111110101;
   5401: result <= 12'b001111110101;
   5402: result <= 12'b001111110101;
   5403: result <= 12'b001111110110;
   5404: result <= 12'b001111110110;
   5405: result <= 12'b001111110110;
   5406: result <= 12'b001111110110;
   5407: result <= 12'b001111110110;
   5408: result <= 12'b001111110110;
   5409: result <= 12'b001111110111;
   5410: result <= 12'b001111110111;
   5411: result <= 12'b001111110111;
   5412: result <= 12'b001111110111;
   5413: result <= 12'b001111110111;
   5414: result <= 12'b001111110111;
   5415: result <= 12'b001111111000;
   5416: result <= 12'b001111111000;
   5417: result <= 12'b001111111000;
   5418: result <= 12'b001111111000;
   5419: result <= 12'b001111111000;
   5420: result <= 12'b001111111000;
   5421: result <= 12'b001111111001;
   5422: result <= 12'b001111111001;
   5423: result <= 12'b001111111001;
   5424: result <= 12'b001111111001;
   5425: result <= 12'b001111111001;
   5426: result <= 12'b001111111001;
   5427: result <= 12'b001111111010;
   5428: result <= 12'b001111111010;
   5429: result <= 12'b001111111010;
   5430: result <= 12'b001111111010;
   5431: result <= 12'b001111111010;
   5432: result <= 12'b001111111011;
   5433: result <= 12'b001111111011;
   5434: result <= 12'b001111111011;
   5435: result <= 12'b001111111011;
   5436: result <= 12'b001111111011;
   5437: result <= 12'b001111111011;
   5438: result <= 12'b001111111100;
   5439: result <= 12'b001111111100;
   5440: result <= 12'b001111111100;
   5441: result <= 12'b001111111100;
   5442: result <= 12'b001111111100;
   5443: result <= 12'b001111111100;
   5444: result <= 12'b001111111101;
   5445: result <= 12'b001111111101;
   5446: result <= 12'b001111111101;
   5447: result <= 12'b001111111101;
   5448: result <= 12'b001111111101;
   5449: result <= 12'b001111111101;
   5450: result <= 12'b001111111110;
   5451: result <= 12'b001111111110;
   5452: result <= 12'b001111111110;
   5453: result <= 12'b001111111110;
   5454: result <= 12'b001111111110;
   5455: result <= 12'b001111111110;
   5456: result <= 12'b001111111111;
   5457: result <= 12'b001111111111;
   5458: result <= 12'b001111111111;
   5459: result <= 12'b001111111111;
   5460: result <= 12'b001111111111;
   5461: result <= 12'b001111111111;
   5462: result <= 12'b010000000000;
   5463: result <= 12'b010000000000;
   5464: result <= 12'b010000000000;
   5465: result <= 12'b010000000000;
   5466: result <= 12'b010000000000;
   5467: result <= 12'b010000000000;
   5468: result <= 12'b010000000001;
   5469: result <= 12'b010000000001;
   5470: result <= 12'b010000000001;
   5471: result <= 12'b010000000001;
   5472: result <= 12'b010000000001;
   5473: result <= 12'b010000000001;
   5474: result <= 12'b010000000010;
   5475: result <= 12'b010000000010;
   5476: result <= 12'b010000000010;
   5477: result <= 12'b010000000010;
   5478: result <= 12'b010000000010;
   5479: result <= 12'b010000000011;
   5480: result <= 12'b010000000011;
   5481: result <= 12'b010000000011;
   5482: result <= 12'b010000000011;
   5483: result <= 12'b010000000011;
   5484: result <= 12'b010000000011;
   5485: result <= 12'b010000000100;
   5486: result <= 12'b010000000100;
   5487: result <= 12'b010000000100;
   5488: result <= 12'b010000000100;
   5489: result <= 12'b010000000100;
   5490: result <= 12'b010000000100;
   5491: result <= 12'b010000000101;
   5492: result <= 12'b010000000101;
   5493: result <= 12'b010000000101;
   5494: result <= 12'b010000000101;
   5495: result <= 12'b010000000101;
   5496: result <= 12'b010000000101;
   5497: result <= 12'b010000000110;
   5498: result <= 12'b010000000110;
   5499: result <= 12'b010000000110;
   5500: result <= 12'b010000000110;
   5501: result <= 12'b010000000110;
   5502: result <= 12'b010000000110;
   5503: result <= 12'b010000000111;
   5504: result <= 12'b010000000111;
   5505: result <= 12'b010000000111;
   5506: result <= 12'b010000000111;
   5507: result <= 12'b010000000111;
   5508: result <= 12'b010000000111;
   5509: result <= 12'b010000001000;
   5510: result <= 12'b010000001000;
   5511: result <= 12'b010000001000;
   5512: result <= 12'b010000001000;
   5513: result <= 12'b010000001000;
   5514: result <= 12'b010000001000;
   5515: result <= 12'b010000001001;
   5516: result <= 12'b010000001001;
   5517: result <= 12'b010000001001;
   5518: result <= 12'b010000001001;
   5519: result <= 12'b010000001001;
   5520: result <= 12'b010000001001;
   5521: result <= 12'b010000001010;
   5522: result <= 12'b010000001010;
   5523: result <= 12'b010000001010;
   5524: result <= 12'b010000001010;
   5525: result <= 12'b010000001010;
   5526: result <= 12'b010000001010;
   5527: result <= 12'b010000001011;
   5528: result <= 12'b010000001011;
   5529: result <= 12'b010000001011;
   5530: result <= 12'b010000001011;
   5531: result <= 12'b010000001011;
   5532: result <= 12'b010000001011;
   5533: result <= 12'b010000001100;
   5534: result <= 12'b010000001100;
   5535: result <= 12'b010000001100;
   5536: result <= 12'b010000001100;
   5537: result <= 12'b010000001100;
   5538: result <= 12'b010000001101;
   5539: result <= 12'b010000001101;
   5540: result <= 12'b010000001101;
   5541: result <= 12'b010000001101;
   5542: result <= 12'b010000001101;
   5543: result <= 12'b010000001101;
   5544: result <= 12'b010000001110;
   5545: result <= 12'b010000001110;
   5546: result <= 12'b010000001110;
   5547: result <= 12'b010000001110;
   5548: result <= 12'b010000001110;
   5549: result <= 12'b010000001110;
   5550: result <= 12'b010000001111;
   5551: result <= 12'b010000001111;
   5552: result <= 12'b010000001111;
   5553: result <= 12'b010000001111;
   5554: result <= 12'b010000001111;
   5555: result <= 12'b010000001111;
   5556: result <= 12'b010000010000;
   5557: result <= 12'b010000010000;
   5558: result <= 12'b010000010000;
   5559: result <= 12'b010000010000;
   5560: result <= 12'b010000010000;
   5561: result <= 12'b010000010000;
   5562: result <= 12'b010000010001;
   5563: result <= 12'b010000010001;
   5564: result <= 12'b010000010001;
   5565: result <= 12'b010000010001;
   5566: result <= 12'b010000010001;
   5567: result <= 12'b010000010001;
   5568: result <= 12'b010000010010;
   5569: result <= 12'b010000010010;
   5570: result <= 12'b010000010010;
   5571: result <= 12'b010000010010;
   5572: result <= 12'b010000010010;
   5573: result <= 12'b010000010010;
   5574: result <= 12'b010000010011;
   5575: result <= 12'b010000010011;
   5576: result <= 12'b010000010011;
   5577: result <= 12'b010000010011;
   5578: result <= 12'b010000010011;
   5579: result <= 12'b010000010011;
   5580: result <= 12'b010000010100;
   5581: result <= 12'b010000010100;
   5582: result <= 12'b010000010100;
   5583: result <= 12'b010000010100;
   5584: result <= 12'b010000010100;
   5585: result <= 12'b010000010100;
   5586: result <= 12'b010000010101;
   5587: result <= 12'b010000010101;
   5588: result <= 12'b010000010101;
   5589: result <= 12'b010000010101;
   5590: result <= 12'b010000010101;
   5591: result <= 12'b010000010101;
   5592: result <= 12'b010000010110;
   5593: result <= 12'b010000010110;
   5594: result <= 12'b010000010110;
   5595: result <= 12'b010000010110;
   5596: result <= 12'b010000010110;
   5597: result <= 12'b010000010110;
   5598: result <= 12'b010000010111;
   5599: result <= 12'b010000010111;
   5600: result <= 12'b010000010111;
   5601: result <= 12'b010000010111;
   5602: result <= 12'b010000010111;
   5603: result <= 12'b010000010111;
   5604: result <= 12'b010000011000;
   5605: result <= 12'b010000011000;
   5606: result <= 12'b010000011000;
   5607: result <= 12'b010000011000;
   5608: result <= 12'b010000011000;
   5609: result <= 12'b010000011001;
   5610: result <= 12'b010000011001;
   5611: result <= 12'b010000011001;
   5612: result <= 12'b010000011001;
   5613: result <= 12'b010000011001;
   5614: result <= 12'b010000011001;
   5615: result <= 12'b010000011010;
   5616: result <= 12'b010000011010;
   5617: result <= 12'b010000011010;
   5618: result <= 12'b010000011010;
   5619: result <= 12'b010000011010;
   5620: result <= 12'b010000011010;
   5621: result <= 12'b010000011011;
   5622: result <= 12'b010000011011;
   5623: result <= 12'b010000011011;
   5624: result <= 12'b010000011011;
   5625: result <= 12'b010000011011;
   5626: result <= 12'b010000011011;
   5627: result <= 12'b010000011100;
   5628: result <= 12'b010000011100;
   5629: result <= 12'b010000011100;
   5630: result <= 12'b010000011100;
   5631: result <= 12'b010000011100;
   5632: result <= 12'b010000011100;
   5633: result <= 12'b010000011101;
   5634: result <= 12'b010000011101;
   5635: result <= 12'b010000011101;
   5636: result <= 12'b010000011101;
   5637: result <= 12'b010000011101;
   5638: result <= 12'b010000011101;
   5639: result <= 12'b010000011110;
   5640: result <= 12'b010000011110;
   5641: result <= 12'b010000011110;
   5642: result <= 12'b010000011110;
   5643: result <= 12'b010000011110;
   5644: result <= 12'b010000011110;
   5645: result <= 12'b010000011111;
   5646: result <= 12'b010000011111;
   5647: result <= 12'b010000011111;
   5648: result <= 12'b010000011111;
   5649: result <= 12'b010000011111;
   5650: result <= 12'b010000011111;
   5651: result <= 12'b010000100000;
   5652: result <= 12'b010000100000;
   5653: result <= 12'b010000100000;
   5654: result <= 12'b010000100000;
   5655: result <= 12'b010000100000;
   5656: result <= 12'b010000100000;
   5657: result <= 12'b010000100001;
   5658: result <= 12'b010000100001;
   5659: result <= 12'b010000100001;
   5660: result <= 12'b010000100001;
   5661: result <= 12'b010000100001;
   5662: result <= 12'b010000100001;
   5663: result <= 12'b010000100010;
   5664: result <= 12'b010000100010;
   5665: result <= 12'b010000100010;
   5666: result <= 12'b010000100010;
   5667: result <= 12'b010000100010;
   5668: result <= 12'b010000100010;
   5669: result <= 12'b010000100011;
   5670: result <= 12'b010000100011;
   5671: result <= 12'b010000100011;
   5672: result <= 12'b010000100011;
   5673: result <= 12'b010000100011;
   5674: result <= 12'b010000100011;
   5675: result <= 12'b010000100100;
   5676: result <= 12'b010000100100;
   5677: result <= 12'b010000100100;
   5678: result <= 12'b010000100100;
   5679: result <= 12'b010000100100;
   5680: result <= 12'b010000100100;
   5681: result <= 12'b010000100101;
   5682: result <= 12'b010000100101;
   5683: result <= 12'b010000100101;
   5684: result <= 12'b010000100101;
   5685: result <= 12'b010000100101;
   5686: result <= 12'b010000100101;
   5687: result <= 12'b010000100110;
   5688: result <= 12'b010000100110;
   5689: result <= 12'b010000100110;
   5690: result <= 12'b010000100110;
   5691: result <= 12'b010000100110;
   5692: result <= 12'b010000100110;
   5693: result <= 12'b010000100111;
   5694: result <= 12'b010000100111;
   5695: result <= 12'b010000100111;
   5696: result <= 12'b010000100111;
   5697: result <= 12'b010000100111;
   5698: result <= 12'b010000100111;
   5699: result <= 12'b010000101000;
   5700: result <= 12'b010000101000;
   5701: result <= 12'b010000101000;
   5702: result <= 12'b010000101000;
   5703: result <= 12'b010000101000;
   5704: result <= 12'b010000101000;
   5705: result <= 12'b010000101001;
   5706: result <= 12'b010000101001;
   5707: result <= 12'b010000101001;
   5708: result <= 12'b010000101001;
   5709: result <= 12'b010000101001;
   5710: result <= 12'b010000101001;
   5711: result <= 12'b010000101010;
   5712: result <= 12'b010000101010;
   5713: result <= 12'b010000101010;
   5714: result <= 12'b010000101010;
   5715: result <= 12'b010000101010;
   5716: result <= 12'b010000101010;
   5717: result <= 12'b010000101011;
   5718: result <= 12'b010000101011;
   5719: result <= 12'b010000101011;
   5720: result <= 12'b010000101011;
   5721: result <= 12'b010000101011;
   5722: result <= 12'b010000101100;
   5723: result <= 12'b010000101100;
   5724: result <= 12'b010000101100;
   5725: result <= 12'b010000101100;
   5726: result <= 12'b010000101100;
   5727: result <= 12'b010000101100;
   5728: result <= 12'b010000101101;
   5729: result <= 12'b010000101101;
   5730: result <= 12'b010000101101;
   5731: result <= 12'b010000101101;
   5732: result <= 12'b010000101101;
   5733: result <= 12'b010000101101;
   5734: result <= 12'b010000101110;
   5735: result <= 12'b010000101110;
   5736: result <= 12'b010000101110;
   5737: result <= 12'b010000101110;
   5738: result <= 12'b010000101110;
   5739: result <= 12'b010000101110;
   5740: result <= 12'b010000101111;
   5741: result <= 12'b010000101111;
   5742: result <= 12'b010000101111;
   5743: result <= 12'b010000101111;
   5744: result <= 12'b010000101111;
   5745: result <= 12'b010000101111;
   5746: result <= 12'b010000110000;
   5747: result <= 12'b010000110000;
   5748: result <= 12'b010000110000;
   5749: result <= 12'b010000110000;
   5750: result <= 12'b010000110000;
   5751: result <= 12'b010000110000;
   5752: result <= 12'b010000110001;
   5753: result <= 12'b010000110001;
   5754: result <= 12'b010000110001;
   5755: result <= 12'b010000110001;
   5756: result <= 12'b010000110001;
   5757: result <= 12'b010000110001;
   5758: result <= 12'b010000110010;
   5759: result <= 12'b010000110010;
   5760: result <= 12'b010000110010;
   5761: result <= 12'b010000110010;
   5762: result <= 12'b010000110010;
   5763: result <= 12'b010000110010;
   5764: result <= 12'b010000110011;
   5765: result <= 12'b010000110011;
   5766: result <= 12'b010000110011;
   5767: result <= 12'b010000110011;
   5768: result <= 12'b010000110011;
   5769: result <= 12'b010000110011;
   5770: result <= 12'b010000110100;
   5771: result <= 12'b010000110100;
   5772: result <= 12'b010000110100;
   5773: result <= 12'b010000110100;
   5774: result <= 12'b010000110100;
   5775: result <= 12'b010000110100;
   5776: result <= 12'b010000110101;
   5777: result <= 12'b010000110101;
   5778: result <= 12'b010000110101;
   5779: result <= 12'b010000110101;
   5780: result <= 12'b010000110101;
   5781: result <= 12'b010000110101;
   5782: result <= 12'b010000110110;
   5783: result <= 12'b010000110110;
   5784: result <= 12'b010000110110;
   5785: result <= 12'b010000110110;
   5786: result <= 12'b010000110110;
   5787: result <= 12'b010000110110;
   5788: result <= 12'b010000110111;
   5789: result <= 12'b010000110111;
   5790: result <= 12'b010000110111;
   5791: result <= 12'b010000110111;
   5792: result <= 12'b010000110111;
   5793: result <= 12'b010000110111;
   5794: result <= 12'b010000111000;
   5795: result <= 12'b010000111000;
   5796: result <= 12'b010000111000;
   5797: result <= 12'b010000111000;
   5798: result <= 12'b010000111000;
   5799: result <= 12'b010000111000;
   5800: result <= 12'b010000111001;
   5801: result <= 12'b010000111001;
   5802: result <= 12'b010000111001;
   5803: result <= 12'b010000111001;
   5804: result <= 12'b010000111001;
   5805: result <= 12'b010000111001;
   5806: result <= 12'b010000111010;
   5807: result <= 12'b010000111010;
   5808: result <= 12'b010000111010;
   5809: result <= 12'b010000111010;
   5810: result <= 12'b010000111010;
   5811: result <= 12'b010000111010;
   5812: result <= 12'b010000111011;
   5813: result <= 12'b010000111011;
   5814: result <= 12'b010000111011;
   5815: result <= 12'b010000111011;
   5816: result <= 12'b010000111011;
   5817: result <= 12'b010000111011;
   5818: result <= 12'b010000111100;
   5819: result <= 12'b010000111100;
   5820: result <= 12'b010000111100;
   5821: result <= 12'b010000111100;
   5822: result <= 12'b010000111100;
   5823: result <= 12'b010000111100;
   5824: result <= 12'b010000111101;
   5825: result <= 12'b010000111101;
   5826: result <= 12'b010000111101;
   5827: result <= 12'b010000111101;
   5828: result <= 12'b010000111101;
   5829: result <= 12'b010000111101;
   5830: result <= 12'b010000111110;
   5831: result <= 12'b010000111110;
   5832: result <= 12'b010000111110;
   5833: result <= 12'b010000111110;
   5834: result <= 12'b010000111110;
   5835: result <= 12'b010000111110;
   5836: result <= 12'b010000111111;
   5837: result <= 12'b010000111111;
   5838: result <= 12'b010000111111;
   5839: result <= 12'b010000111111;
   5840: result <= 12'b010000111111;
   5841: result <= 12'b010000111111;
   5842: result <= 12'b010001000000;
   5843: result <= 12'b010001000000;
   5844: result <= 12'b010001000000;
   5845: result <= 12'b010001000000;
   5846: result <= 12'b010001000000;
   5847: result <= 12'b010001000000;
   5848: result <= 12'b010001000001;
   5849: result <= 12'b010001000001;
   5850: result <= 12'b010001000001;
   5851: result <= 12'b010001000001;
   5852: result <= 12'b010001000001;
   5853: result <= 12'b010001000001;
   5854: result <= 12'b010001000010;
   5855: result <= 12'b010001000010;
   5856: result <= 12'b010001000010;
   5857: result <= 12'b010001000010;
   5858: result <= 12'b010001000010;
   5859: result <= 12'b010001000010;
   5860: result <= 12'b010001000011;
   5861: result <= 12'b010001000011;
   5862: result <= 12'b010001000011;
   5863: result <= 12'b010001000011;
   5864: result <= 12'b010001000011;
   5865: result <= 12'b010001000011;
   5866: result <= 12'b010001000100;
   5867: result <= 12'b010001000100;
   5868: result <= 12'b010001000100;
   5869: result <= 12'b010001000100;
   5870: result <= 12'b010001000100;
   5871: result <= 12'b010001000100;
   5872: result <= 12'b010001000101;
   5873: result <= 12'b010001000101;
   5874: result <= 12'b010001000101;
   5875: result <= 12'b010001000101;
   5876: result <= 12'b010001000101;
   5877: result <= 12'b010001000101;
   5878: result <= 12'b010001000110;
   5879: result <= 12'b010001000110;
   5880: result <= 12'b010001000110;
   5881: result <= 12'b010001000110;
   5882: result <= 12'b010001000110;
   5883: result <= 12'b010001000110;
   5884: result <= 12'b010001000111;
   5885: result <= 12'b010001000111;
   5886: result <= 12'b010001000111;
   5887: result <= 12'b010001000111;
   5888: result <= 12'b010001000111;
   5889: result <= 12'b010001000111;
   5890: result <= 12'b010001001000;
   5891: result <= 12'b010001001000;
   5892: result <= 12'b010001001000;
   5893: result <= 12'b010001001000;
   5894: result <= 12'b010001001000;
   5895: result <= 12'b010001001000;
   5896: result <= 12'b010001001001;
   5897: result <= 12'b010001001001;
   5898: result <= 12'b010001001001;
   5899: result <= 12'b010001001001;
   5900: result <= 12'b010001001001;
   5901: result <= 12'b010001001001;
   5902: result <= 12'b010001001001;
   5903: result <= 12'b010001001010;
   5904: result <= 12'b010001001010;
   5905: result <= 12'b010001001010;
   5906: result <= 12'b010001001010;
   5907: result <= 12'b010001001010;
   5908: result <= 12'b010001001010;
   5909: result <= 12'b010001001011;
   5910: result <= 12'b010001001011;
   5911: result <= 12'b010001001011;
   5912: result <= 12'b010001001011;
   5913: result <= 12'b010001001011;
   5914: result <= 12'b010001001011;
   5915: result <= 12'b010001001100;
   5916: result <= 12'b010001001100;
   5917: result <= 12'b010001001100;
   5918: result <= 12'b010001001100;
   5919: result <= 12'b010001001100;
   5920: result <= 12'b010001001100;
   5921: result <= 12'b010001001101;
   5922: result <= 12'b010001001101;
   5923: result <= 12'b010001001101;
   5924: result <= 12'b010001001101;
   5925: result <= 12'b010001001101;
   5926: result <= 12'b010001001101;
   5927: result <= 12'b010001001110;
   5928: result <= 12'b010001001110;
   5929: result <= 12'b010001001110;
   5930: result <= 12'b010001001110;
   5931: result <= 12'b010001001110;
   5932: result <= 12'b010001001110;
   5933: result <= 12'b010001001111;
   5934: result <= 12'b010001001111;
   5935: result <= 12'b010001001111;
   5936: result <= 12'b010001001111;
   5937: result <= 12'b010001001111;
   5938: result <= 12'b010001001111;
   5939: result <= 12'b010001010000;
   5940: result <= 12'b010001010000;
   5941: result <= 12'b010001010000;
   5942: result <= 12'b010001010000;
   5943: result <= 12'b010001010000;
   5944: result <= 12'b010001010000;
   5945: result <= 12'b010001010001;
   5946: result <= 12'b010001010001;
   5947: result <= 12'b010001010001;
   5948: result <= 12'b010001010001;
   5949: result <= 12'b010001010001;
   5950: result <= 12'b010001010001;
   5951: result <= 12'b010001010010;
   5952: result <= 12'b010001010010;
   5953: result <= 12'b010001010010;
   5954: result <= 12'b010001010010;
   5955: result <= 12'b010001010010;
   5956: result <= 12'b010001010010;
   5957: result <= 12'b010001010011;
   5958: result <= 12'b010001010011;
   5959: result <= 12'b010001010011;
   5960: result <= 12'b010001010011;
   5961: result <= 12'b010001010011;
   5962: result <= 12'b010001010011;
   5963: result <= 12'b010001010100;
   5964: result <= 12'b010001010100;
   5965: result <= 12'b010001010100;
   5966: result <= 12'b010001010100;
   5967: result <= 12'b010001010100;
   5968: result <= 12'b010001010100;
   5969: result <= 12'b010001010101;
   5970: result <= 12'b010001010101;
   5971: result <= 12'b010001010101;
   5972: result <= 12'b010001010101;
   5973: result <= 12'b010001010101;
   5974: result <= 12'b010001010101;
   5975: result <= 12'b010001010110;
   5976: result <= 12'b010001010110;
   5977: result <= 12'b010001010110;
   5978: result <= 12'b010001010110;
   5979: result <= 12'b010001010110;
   5980: result <= 12'b010001010110;
   5981: result <= 12'b010001010111;
   5982: result <= 12'b010001010111;
   5983: result <= 12'b010001010111;
   5984: result <= 12'b010001010111;
   5985: result <= 12'b010001010111;
   5986: result <= 12'b010001010111;
   5987: result <= 12'b010001011000;
   5988: result <= 12'b010001011000;
   5989: result <= 12'b010001011000;
   5990: result <= 12'b010001011000;
   5991: result <= 12'b010001011000;
   5992: result <= 12'b010001011000;
   5993: result <= 12'b010001011001;
   5994: result <= 12'b010001011001;
   5995: result <= 12'b010001011001;
   5996: result <= 12'b010001011001;
   5997: result <= 12'b010001011001;
   5998: result <= 12'b010001011001;
   5999: result <= 12'b010001011010;
   6000: result <= 12'b010001011010;
   6001: result <= 12'b010001011010;
   6002: result <= 12'b010001011010;
   6003: result <= 12'b010001011010;
   6004: result <= 12'b010001011010;
   6005: result <= 12'b010001011011;
   6006: result <= 12'b010001011011;
   6007: result <= 12'b010001011011;
   6008: result <= 12'b010001011011;
   6009: result <= 12'b010001011011;
   6010: result <= 12'b010001011011;
   6011: result <= 12'b010001011100;
   6012: result <= 12'b010001011100;
   6013: result <= 12'b010001011100;
   6014: result <= 12'b010001011100;
   6015: result <= 12'b010001011100;
   6016: result <= 12'b010001011100;
   6017: result <= 12'b010001011100;
   6018: result <= 12'b010001011101;
   6019: result <= 12'b010001011101;
   6020: result <= 12'b010001011101;
   6021: result <= 12'b010001011101;
   6022: result <= 12'b010001011101;
   6023: result <= 12'b010001011101;
   6024: result <= 12'b010001011110;
   6025: result <= 12'b010001011110;
   6026: result <= 12'b010001011110;
   6027: result <= 12'b010001011110;
   6028: result <= 12'b010001011110;
   6029: result <= 12'b010001011110;
   6030: result <= 12'b010001011111;
   6031: result <= 12'b010001011111;
   6032: result <= 12'b010001011111;
   6033: result <= 12'b010001011111;
   6034: result <= 12'b010001011111;
   6035: result <= 12'b010001011111;
   6036: result <= 12'b010001100000;
   6037: result <= 12'b010001100000;
   6038: result <= 12'b010001100000;
   6039: result <= 12'b010001100000;
   6040: result <= 12'b010001100000;
   6041: result <= 12'b010001100000;
   6042: result <= 12'b010001100001;
   6043: result <= 12'b010001100001;
   6044: result <= 12'b010001100001;
   6045: result <= 12'b010001100001;
   6046: result <= 12'b010001100001;
   6047: result <= 12'b010001100001;
   6048: result <= 12'b010001100010;
   6049: result <= 12'b010001100010;
   6050: result <= 12'b010001100010;
   6051: result <= 12'b010001100010;
   6052: result <= 12'b010001100010;
   6053: result <= 12'b010001100010;
   6054: result <= 12'b010001100011;
   6055: result <= 12'b010001100011;
   6056: result <= 12'b010001100011;
   6057: result <= 12'b010001100011;
   6058: result <= 12'b010001100011;
   6059: result <= 12'b010001100011;
   6060: result <= 12'b010001100100;
   6061: result <= 12'b010001100100;
   6062: result <= 12'b010001100100;
   6063: result <= 12'b010001100100;
   6064: result <= 12'b010001100100;
   6065: result <= 12'b010001100100;
   6066: result <= 12'b010001100101;
   6067: result <= 12'b010001100101;
   6068: result <= 12'b010001100101;
   6069: result <= 12'b010001100101;
   6070: result <= 12'b010001100101;
   6071: result <= 12'b010001100101;
   6072: result <= 12'b010001100110;
   6073: result <= 12'b010001100110;
   6074: result <= 12'b010001100110;
   6075: result <= 12'b010001100110;
   6076: result <= 12'b010001100110;
   6077: result <= 12'b010001100110;
   6078: result <= 12'b010001100111;
   6079: result <= 12'b010001100111;
   6080: result <= 12'b010001100111;
   6081: result <= 12'b010001100111;
   6082: result <= 12'b010001100111;
   6083: result <= 12'b010001100111;
   6084: result <= 12'b010001100111;
   6085: result <= 12'b010001101000;
   6086: result <= 12'b010001101000;
   6087: result <= 12'b010001101000;
   6088: result <= 12'b010001101000;
   6089: result <= 12'b010001101000;
   6090: result <= 12'b010001101000;
   6091: result <= 12'b010001101001;
   6092: result <= 12'b010001101001;
   6093: result <= 12'b010001101001;
   6094: result <= 12'b010001101001;
   6095: result <= 12'b010001101001;
   6096: result <= 12'b010001101001;
   6097: result <= 12'b010001101010;
   6098: result <= 12'b010001101010;
   6099: result <= 12'b010001101010;
   6100: result <= 12'b010001101010;
   6101: result <= 12'b010001101010;
   6102: result <= 12'b010001101010;
   6103: result <= 12'b010001101011;
   6104: result <= 12'b010001101011;
   6105: result <= 12'b010001101011;
   6106: result <= 12'b010001101011;
   6107: result <= 12'b010001101011;
   6108: result <= 12'b010001101011;
   6109: result <= 12'b010001101100;
   6110: result <= 12'b010001101100;
   6111: result <= 12'b010001101100;
   6112: result <= 12'b010001101100;
   6113: result <= 12'b010001101100;
   6114: result <= 12'b010001101100;
   6115: result <= 12'b010001101101;
   6116: result <= 12'b010001101101;
   6117: result <= 12'b010001101101;
   6118: result <= 12'b010001101101;
   6119: result <= 12'b010001101101;
   6120: result <= 12'b010001101101;
   6121: result <= 12'b010001101110;
   6122: result <= 12'b010001101110;
   6123: result <= 12'b010001101110;
   6124: result <= 12'b010001101110;
   6125: result <= 12'b010001101110;
   6126: result <= 12'b010001101110;
   6127: result <= 12'b010001101111;
   6128: result <= 12'b010001101111;
   6129: result <= 12'b010001101111;
   6130: result <= 12'b010001101111;
   6131: result <= 12'b010001101111;
   6132: result <= 12'b010001101111;
   6133: result <= 12'b010001110000;
   6134: result <= 12'b010001110000;
   6135: result <= 12'b010001110000;
   6136: result <= 12'b010001110000;
   6137: result <= 12'b010001110000;
   6138: result <= 12'b010001110000;
   6139: result <= 12'b010001110000;
   6140: result <= 12'b010001110001;
   6141: result <= 12'b010001110001;
   6142: result <= 12'b010001110001;
   6143: result <= 12'b010001110001;
   6144: result <= 12'b010001110001;
   6145: result <= 12'b010001110001;
   6146: result <= 12'b010001110010;
   6147: result <= 12'b010001110010;
   6148: result <= 12'b010001110010;
   6149: result <= 12'b010001110010;
   6150: result <= 12'b010001110010;
   6151: result <= 12'b010001110010;
   6152: result <= 12'b010001110011;
   6153: result <= 12'b010001110011;
   6154: result <= 12'b010001110011;
   6155: result <= 12'b010001110011;
   6156: result <= 12'b010001110011;
   6157: result <= 12'b010001110011;
   6158: result <= 12'b010001110100;
   6159: result <= 12'b010001110100;
   6160: result <= 12'b010001110100;
   6161: result <= 12'b010001110100;
   6162: result <= 12'b010001110100;
   6163: result <= 12'b010001110100;
   6164: result <= 12'b010001110101;
   6165: result <= 12'b010001110101;
   6166: result <= 12'b010001110101;
   6167: result <= 12'b010001110101;
   6168: result <= 12'b010001110101;
   6169: result <= 12'b010001110101;
   6170: result <= 12'b010001110110;
   6171: result <= 12'b010001110110;
   6172: result <= 12'b010001110110;
   6173: result <= 12'b010001110110;
   6174: result <= 12'b010001110110;
   6175: result <= 12'b010001110110;
   6176: result <= 12'b010001110111;
   6177: result <= 12'b010001110111;
   6178: result <= 12'b010001110111;
   6179: result <= 12'b010001110111;
   6180: result <= 12'b010001110111;
   6181: result <= 12'b010001110111;
   6182: result <= 12'b010001111000;
   6183: result <= 12'b010001111000;
   6184: result <= 12'b010001111000;
   6185: result <= 12'b010001111000;
   6186: result <= 12'b010001111000;
   6187: result <= 12'b010001111000;
   6188: result <= 12'b010001111000;
   6189: result <= 12'b010001111001;
   6190: result <= 12'b010001111001;
   6191: result <= 12'b010001111001;
   6192: result <= 12'b010001111001;
   6193: result <= 12'b010001111001;
   6194: result <= 12'b010001111001;
   6195: result <= 12'b010001111010;
   6196: result <= 12'b010001111010;
   6197: result <= 12'b010001111010;
   6198: result <= 12'b010001111010;
   6199: result <= 12'b010001111010;
   6200: result <= 12'b010001111010;
   6201: result <= 12'b010001111011;
   6202: result <= 12'b010001111011;
   6203: result <= 12'b010001111011;
   6204: result <= 12'b010001111011;
   6205: result <= 12'b010001111011;
   6206: result <= 12'b010001111011;
   6207: result <= 12'b010001111100;
   6208: result <= 12'b010001111100;
   6209: result <= 12'b010001111100;
   6210: result <= 12'b010001111100;
   6211: result <= 12'b010001111100;
   6212: result <= 12'b010001111100;
   6213: result <= 12'b010001111101;
   6214: result <= 12'b010001111101;
   6215: result <= 12'b010001111101;
   6216: result <= 12'b010001111101;
   6217: result <= 12'b010001111101;
   6218: result <= 12'b010001111101;
   6219: result <= 12'b010001111110;
   6220: result <= 12'b010001111110;
   6221: result <= 12'b010001111110;
   6222: result <= 12'b010001111110;
   6223: result <= 12'b010001111110;
   6224: result <= 12'b010001111110;
   6225: result <= 12'b010001111110;
   6226: result <= 12'b010001111111;
   6227: result <= 12'b010001111111;
   6228: result <= 12'b010001111111;
   6229: result <= 12'b010001111111;
   6230: result <= 12'b010001111111;
   6231: result <= 12'b010001111111;
   6232: result <= 12'b010010000000;
   6233: result <= 12'b010010000000;
   6234: result <= 12'b010010000000;
   6235: result <= 12'b010010000000;
   6236: result <= 12'b010010000000;
   6237: result <= 12'b010010000000;
   6238: result <= 12'b010010000001;
   6239: result <= 12'b010010000001;
   6240: result <= 12'b010010000001;
   6241: result <= 12'b010010000001;
   6242: result <= 12'b010010000001;
   6243: result <= 12'b010010000001;
   6244: result <= 12'b010010000010;
   6245: result <= 12'b010010000010;
   6246: result <= 12'b010010000010;
   6247: result <= 12'b010010000010;
   6248: result <= 12'b010010000010;
   6249: result <= 12'b010010000010;
   6250: result <= 12'b010010000011;
   6251: result <= 12'b010010000011;
   6252: result <= 12'b010010000011;
   6253: result <= 12'b010010000011;
   6254: result <= 12'b010010000011;
   6255: result <= 12'b010010000011;
   6256: result <= 12'b010010000100;
   6257: result <= 12'b010010000100;
   6258: result <= 12'b010010000100;
   6259: result <= 12'b010010000100;
   6260: result <= 12'b010010000100;
   6261: result <= 12'b010010000100;
   6262: result <= 12'b010010000100;
   6263: result <= 12'b010010000101;
   6264: result <= 12'b010010000101;
   6265: result <= 12'b010010000101;
   6266: result <= 12'b010010000101;
   6267: result <= 12'b010010000101;
   6268: result <= 12'b010010000101;
   6269: result <= 12'b010010000110;
   6270: result <= 12'b010010000110;
   6271: result <= 12'b010010000110;
   6272: result <= 12'b010010000110;
   6273: result <= 12'b010010000110;
   6274: result <= 12'b010010000110;
   6275: result <= 12'b010010000111;
   6276: result <= 12'b010010000111;
   6277: result <= 12'b010010000111;
   6278: result <= 12'b010010000111;
   6279: result <= 12'b010010000111;
   6280: result <= 12'b010010000111;
   6281: result <= 12'b010010001000;
   6282: result <= 12'b010010001000;
   6283: result <= 12'b010010001000;
   6284: result <= 12'b010010001000;
   6285: result <= 12'b010010001000;
   6286: result <= 12'b010010001000;
   6287: result <= 12'b010010001001;
   6288: result <= 12'b010010001001;
   6289: result <= 12'b010010001001;
   6290: result <= 12'b010010001001;
   6291: result <= 12'b010010001001;
   6292: result <= 12'b010010001001;
   6293: result <= 12'b010010001010;
   6294: result <= 12'b010010001010;
   6295: result <= 12'b010010001010;
   6296: result <= 12'b010010001010;
   6297: result <= 12'b010010001010;
   6298: result <= 12'b010010001010;
   6299: result <= 12'b010010001010;
   6300: result <= 12'b010010001011;
   6301: result <= 12'b010010001011;
   6302: result <= 12'b010010001011;
   6303: result <= 12'b010010001011;
   6304: result <= 12'b010010001011;
   6305: result <= 12'b010010001011;
   6306: result <= 12'b010010001100;
   6307: result <= 12'b010010001100;
   6308: result <= 12'b010010001100;
   6309: result <= 12'b010010001100;
   6310: result <= 12'b010010001100;
   6311: result <= 12'b010010001100;
   6312: result <= 12'b010010001101;
   6313: result <= 12'b010010001101;
   6314: result <= 12'b010010001101;
   6315: result <= 12'b010010001101;
   6316: result <= 12'b010010001101;
   6317: result <= 12'b010010001101;
   6318: result <= 12'b010010001110;
   6319: result <= 12'b010010001110;
   6320: result <= 12'b010010001110;
   6321: result <= 12'b010010001110;
   6322: result <= 12'b010010001110;
   6323: result <= 12'b010010001110;
   6324: result <= 12'b010010001111;
   6325: result <= 12'b010010001111;
   6326: result <= 12'b010010001111;
   6327: result <= 12'b010010001111;
   6328: result <= 12'b010010001111;
   6329: result <= 12'b010010001111;
   6330: result <= 12'b010010001111;
   6331: result <= 12'b010010010000;
   6332: result <= 12'b010010010000;
   6333: result <= 12'b010010010000;
   6334: result <= 12'b010010010000;
   6335: result <= 12'b010010010000;
   6336: result <= 12'b010010010000;
   6337: result <= 12'b010010010001;
   6338: result <= 12'b010010010001;
   6339: result <= 12'b010010010001;
   6340: result <= 12'b010010010001;
   6341: result <= 12'b010010010001;
   6342: result <= 12'b010010010001;
   6343: result <= 12'b010010010010;
   6344: result <= 12'b010010010010;
   6345: result <= 12'b010010010010;
   6346: result <= 12'b010010010010;
   6347: result <= 12'b010010010010;
   6348: result <= 12'b010010010010;
   6349: result <= 12'b010010010011;
   6350: result <= 12'b010010010011;
   6351: result <= 12'b010010010011;
   6352: result <= 12'b010010010011;
   6353: result <= 12'b010010010011;
   6354: result <= 12'b010010010011;
   6355: result <= 12'b010010010100;
   6356: result <= 12'b010010010100;
   6357: result <= 12'b010010010100;
   6358: result <= 12'b010010010100;
   6359: result <= 12'b010010010100;
   6360: result <= 12'b010010010100;
   6361: result <= 12'b010010010100;
   6362: result <= 12'b010010010101;
   6363: result <= 12'b010010010101;
   6364: result <= 12'b010010010101;
   6365: result <= 12'b010010010101;
   6366: result <= 12'b010010010101;
   6367: result <= 12'b010010010101;
   6368: result <= 12'b010010010110;
   6369: result <= 12'b010010010110;
   6370: result <= 12'b010010010110;
   6371: result <= 12'b010010010110;
   6372: result <= 12'b010010010110;
   6373: result <= 12'b010010010110;
   6374: result <= 12'b010010010111;
   6375: result <= 12'b010010010111;
   6376: result <= 12'b010010010111;
   6377: result <= 12'b010010010111;
   6378: result <= 12'b010010010111;
   6379: result <= 12'b010010010111;
   6380: result <= 12'b010010011000;
   6381: result <= 12'b010010011000;
   6382: result <= 12'b010010011000;
   6383: result <= 12'b010010011000;
   6384: result <= 12'b010010011000;
   6385: result <= 12'b010010011000;
   6386: result <= 12'b010010011001;
   6387: result <= 12'b010010011001;
   6388: result <= 12'b010010011001;
   6389: result <= 12'b010010011001;
   6390: result <= 12'b010010011001;
   6391: result <= 12'b010010011001;
   6392: result <= 12'b010010011001;
   6393: result <= 12'b010010011010;
   6394: result <= 12'b010010011010;
   6395: result <= 12'b010010011010;
   6396: result <= 12'b010010011010;
   6397: result <= 12'b010010011010;
   6398: result <= 12'b010010011010;
   6399: result <= 12'b010010011011;
   6400: result <= 12'b010010011011;
   6401: result <= 12'b010010011011;
   6402: result <= 12'b010010011011;
   6403: result <= 12'b010010011011;
   6404: result <= 12'b010010011011;
   6405: result <= 12'b010010011100;
   6406: result <= 12'b010010011100;
   6407: result <= 12'b010010011100;
   6408: result <= 12'b010010011100;
   6409: result <= 12'b010010011100;
   6410: result <= 12'b010010011100;
   6411: result <= 12'b010010011101;
   6412: result <= 12'b010010011101;
   6413: result <= 12'b010010011101;
   6414: result <= 12'b010010011101;
   6415: result <= 12'b010010011101;
   6416: result <= 12'b010010011101;
   6417: result <= 12'b010010011101;
   6418: result <= 12'b010010011110;
   6419: result <= 12'b010010011110;
   6420: result <= 12'b010010011110;
   6421: result <= 12'b010010011110;
   6422: result <= 12'b010010011110;
   6423: result <= 12'b010010011110;
   6424: result <= 12'b010010011111;
   6425: result <= 12'b010010011111;
   6426: result <= 12'b010010011111;
   6427: result <= 12'b010010011111;
   6428: result <= 12'b010010011111;
   6429: result <= 12'b010010011111;
   6430: result <= 12'b010010100000;
   6431: result <= 12'b010010100000;
   6432: result <= 12'b010010100000;
   6433: result <= 12'b010010100000;
   6434: result <= 12'b010010100000;
   6435: result <= 12'b010010100000;
   6436: result <= 12'b010010100001;
   6437: result <= 12'b010010100001;
   6438: result <= 12'b010010100001;
   6439: result <= 12'b010010100001;
   6440: result <= 12'b010010100001;
   6441: result <= 12'b010010100001;
   6442: result <= 12'b010010100001;
   6443: result <= 12'b010010100010;
   6444: result <= 12'b010010100010;
   6445: result <= 12'b010010100010;
   6446: result <= 12'b010010100010;
   6447: result <= 12'b010010100010;
   6448: result <= 12'b010010100010;
   6449: result <= 12'b010010100011;
   6450: result <= 12'b010010100011;
   6451: result <= 12'b010010100011;
   6452: result <= 12'b010010100011;
   6453: result <= 12'b010010100011;
   6454: result <= 12'b010010100011;
   6455: result <= 12'b010010100100;
   6456: result <= 12'b010010100100;
   6457: result <= 12'b010010100100;
   6458: result <= 12'b010010100100;
   6459: result <= 12'b010010100100;
   6460: result <= 12'b010010100100;
   6461: result <= 12'b010010100101;
   6462: result <= 12'b010010100101;
   6463: result <= 12'b010010100101;
   6464: result <= 12'b010010100101;
   6465: result <= 12'b010010100101;
   6466: result <= 12'b010010100101;
   6467: result <= 12'b010010100101;
   6468: result <= 12'b010010100110;
   6469: result <= 12'b010010100110;
   6470: result <= 12'b010010100110;
   6471: result <= 12'b010010100110;
   6472: result <= 12'b010010100110;
   6473: result <= 12'b010010100110;
   6474: result <= 12'b010010100111;
   6475: result <= 12'b010010100111;
   6476: result <= 12'b010010100111;
   6477: result <= 12'b010010100111;
   6478: result <= 12'b010010100111;
   6479: result <= 12'b010010100111;
   6480: result <= 12'b010010101000;
   6481: result <= 12'b010010101000;
   6482: result <= 12'b010010101000;
   6483: result <= 12'b010010101000;
   6484: result <= 12'b010010101000;
   6485: result <= 12'b010010101000;
   6486: result <= 12'b010010101001;
   6487: result <= 12'b010010101001;
   6488: result <= 12'b010010101001;
   6489: result <= 12'b010010101001;
   6490: result <= 12'b010010101001;
   6491: result <= 12'b010010101001;
   6492: result <= 12'b010010101001;
   6493: result <= 12'b010010101010;
   6494: result <= 12'b010010101010;
   6495: result <= 12'b010010101010;
   6496: result <= 12'b010010101010;
   6497: result <= 12'b010010101010;
   6498: result <= 12'b010010101010;
   6499: result <= 12'b010010101011;
   6500: result <= 12'b010010101011;
   6501: result <= 12'b010010101011;
   6502: result <= 12'b010010101011;
   6503: result <= 12'b010010101011;
   6504: result <= 12'b010010101011;
   6505: result <= 12'b010010101100;
   6506: result <= 12'b010010101100;
   6507: result <= 12'b010010101100;
   6508: result <= 12'b010010101100;
   6509: result <= 12'b010010101100;
   6510: result <= 12'b010010101100;
   6511: result <= 12'b010010101101;
   6512: result <= 12'b010010101101;
   6513: result <= 12'b010010101101;
   6514: result <= 12'b010010101101;
   6515: result <= 12'b010010101101;
   6516: result <= 12'b010010101101;
   6517: result <= 12'b010010101101;
   6518: result <= 12'b010010101110;
   6519: result <= 12'b010010101110;
   6520: result <= 12'b010010101110;
   6521: result <= 12'b010010101110;
   6522: result <= 12'b010010101110;
   6523: result <= 12'b010010101110;
   6524: result <= 12'b010010101111;
   6525: result <= 12'b010010101111;
   6526: result <= 12'b010010101111;
   6527: result <= 12'b010010101111;
   6528: result <= 12'b010010101111;
   6529: result <= 12'b010010101111;
   6530: result <= 12'b010010110000;
   6531: result <= 12'b010010110000;
   6532: result <= 12'b010010110000;
   6533: result <= 12'b010010110000;
   6534: result <= 12'b010010110000;
   6535: result <= 12'b010010110000;
   6536: result <= 12'b010010110000;
   6537: result <= 12'b010010110001;
   6538: result <= 12'b010010110001;
   6539: result <= 12'b010010110001;
   6540: result <= 12'b010010110001;
   6541: result <= 12'b010010110001;
   6542: result <= 12'b010010110001;
   6543: result <= 12'b010010110010;
   6544: result <= 12'b010010110010;
   6545: result <= 12'b010010110010;
   6546: result <= 12'b010010110010;
   6547: result <= 12'b010010110010;
   6548: result <= 12'b010010110010;
   6549: result <= 12'b010010110011;
   6550: result <= 12'b010010110011;
   6551: result <= 12'b010010110011;
   6552: result <= 12'b010010110011;
   6553: result <= 12'b010010110011;
   6554: result <= 12'b010010110011;
   6555: result <= 12'b010010110100;
   6556: result <= 12'b010010110100;
   6557: result <= 12'b010010110100;
   6558: result <= 12'b010010110100;
   6559: result <= 12'b010010110100;
   6560: result <= 12'b010010110100;
   6561: result <= 12'b010010110100;
   6562: result <= 12'b010010110101;
   6563: result <= 12'b010010110101;
   6564: result <= 12'b010010110101;
   6565: result <= 12'b010010110101;
   6566: result <= 12'b010010110101;
   6567: result <= 12'b010010110101;
   6568: result <= 12'b010010110110;
   6569: result <= 12'b010010110110;
   6570: result <= 12'b010010110110;
   6571: result <= 12'b010010110110;
   6572: result <= 12'b010010110110;
   6573: result <= 12'b010010110110;
   6574: result <= 12'b010010110111;
   6575: result <= 12'b010010110111;
   6576: result <= 12'b010010110111;
   6577: result <= 12'b010010110111;
   6578: result <= 12'b010010110111;
   6579: result <= 12'b010010110111;
   6580: result <= 12'b010010110111;
   6581: result <= 12'b010010111000;
   6582: result <= 12'b010010111000;
   6583: result <= 12'b010010111000;
   6584: result <= 12'b010010111000;
   6585: result <= 12'b010010111000;
   6586: result <= 12'b010010111000;
   6587: result <= 12'b010010111001;
   6588: result <= 12'b010010111001;
   6589: result <= 12'b010010111001;
   6590: result <= 12'b010010111001;
   6591: result <= 12'b010010111001;
   6592: result <= 12'b010010111001;
   6593: result <= 12'b010010111010;
   6594: result <= 12'b010010111010;
   6595: result <= 12'b010010111010;
   6596: result <= 12'b010010111010;
   6597: result <= 12'b010010111010;
   6598: result <= 12'b010010111010;
   6599: result <= 12'b010010111010;
   6600: result <= 12'b010010111011;
   6601: result <= 12'b010010111011;
   6602: result <= 12'b010010111011;
   6603: result <= 12'b010010111011;
   6604: result <= 12'b010010111011;
   6605: result <= 12'b010010111011;
   6606: result <= 12'b010010111100;
   6607: result <= 12'b010010111100;
   6608: result <= 12'b010010111100;
   6609: result <= 12'b010010111100;
   6610: result <= 12'b010010111100;
   6611: result <= 12'b010010111100;
   6612: result <= 12'b010010111101;
   6613: result <= 12'b010010111101;
   6614: result <= 12'b010010111101;
   6615: result <= 12'b010010111101;
   6616: result <= 12'b010010111101;
   6617: result <= 12'b010010111101;
   6618: result <= 12'b010010111101;
   6619: result <= 12'b010010111110;
   6620: result <= 12'b010010111110;
   6621: result <= 12'b010010111110;
   6622: result <= 12'b010010111110;
   6623: result <= 12'b010010111110;
   6624: result <= 12'b010010111110;
   6625: result <= 12'b010010111111;
   6626: result <= 12'b010010111111;
   6627: result <= 12'b010010111111;
   6628: result <= 12'b010010111111;
   6629: result <= 12'b010010111111;
   6630: result <= 12'b010010111111;
   6631: result <= 12'b010011000000;
   6632: result <= 12'b010011000000;
   6633: result <= 12'b010011000000;
   6634: result <= 12'b010011000000;
   6635: result <= 12'b010011000000;
   6636: result <= 12'b010011000000;
   6637: result <= 12'b010011000000;
   6638: result <= 12'b010011000001;
   6639: result <= 12'b010011000001;
   6640: result <= 12'b010011000001;
   6641: result <= 12'b010011000001;
   6642: result <= 12'b010011000001;
   6643: result <= 12'b010011000001;
   6644: result <= 12'b010011000010;
   6645: result <= 12'b010011000010;
   6646: result <= 12'b010011000010;
   6647: result <= 12'b010011000010;
   6648: result <= 12'b010011000010;
   6649: result <= 12'b010011000010;
   6650: result <= 12'b010011000011;
   6651: result <= 12'b010011000011;
   6652: result <= 12'b010011000011;
   6653: result <= 12'b010011000011;
   6654: result <= 12'b010011000011;
   6655: result <= 12'b010011000011;
   6656: result <= 12'b010011000011;
   6657: result <= 12'b010011000100;
   6658: result <= 12'b010011000100;
   6659: result <= 12'b010011000100;
   6660: result <= 12'b010011000100;
   6661: result <= 12'b010011000100;
   6662: result <= 12'b010011000100;
   6663: result <= 12'b010011000101;
   6664: result <= 12'b010011000101;
   6665: result <= 12'b010011000101;
   6666: result <= 12'b010011000101;
   6667: result <= 12'b010011000101;
   6668: result <= 12'b010011000101;
   6669: result <= 12'b010011000110;
   6670: result <= 12'b010011000110;
   6671: result <= 12'b010011000110;
   6672: result <= 12'b010011000110;
   6673: result <= 12'b010011000110;
   6674: result <= 12'b010011000110;
   6675: result <= 12'b010011000110;
   6676: result <= 12'b010011000111;
   6677: result <= 12'b010011000111;
   6678: result <= 12'b010011000111;
   6679: result <= 12'b010011000111;
   6680: result <= 12'b010011000111;
   6681: result <= 12'b010011000111;
   6682: result <= 12'b010011001000;
   6683: result <= 12'b010011001000;
   6684: result <= 12'b010011001000;
   6685: result <= 12'b010011001000;
   6686: result <= 12'b010011001000;
   6687: result <= 12'b010011001000;
   6688: result <= 12'b010011001001;
   6689: result <= 12'b010011001001;
   6690: result <= 12'b010011001001;
   6691: result <= 12'b010011001001;
   6692: result <= 12'b010011001001;
   6693: result <= 12'b010011001001;
   6694: result <= 12'b010011001001;
   6695: result <= 12'b010011001010;
   6696: result <= 12'b010011001010;
   6697: result <= 12'b010011001010;
   6698: result <= 12'b010011001010;
   6699: result <= 12'b010011001010;
   6700: result <= 12'b010011001010;
   6701: result <= 12'b010011001011;
   6702: result <= 12'b010011001011;
   6703: result <= 12'b010011001011;
   6704: result <= 12'b010011001011;
   6705: result <= 12'b010011001011;
   6706: result <= 12'b010011001011;
   6707: result <= 12'b010011001100;
   6708: result <= 12'b010011001100;
   6709: result <= 12'b010011001100;
   6710: result <= 12'b010011001100;
   6711: result <= 12'b010011001100;
   6712: result <= 12'b010011001100;
   6713: result <= 12'b010011001100;
   6714: result <= 12'b010011001101;
   6715: result <= 12'b010011001101;
   6716: result <= 12'b010011001101;
   6717: result <= 12'b010011001101;
   6718: result <= 12'b010011001101;
   6719: result <= 12'b010011001101;
   6720: result <= 12'b010011001110;
   6721: result <= 12'b010011001110;
   6722: result <= 12'b010011001110;
   6723: result <= 12'b010011001110;
   6724: result <= 12'b010011001110;
   6725: result <= 12'b010011001110;
   6726: result <= 12'b010011001111;
   6727: result <= 12'b010011001111;
   6728: result <= 12'b010011001111;
   6729: result <= 12'b010011001111;
   6730: result <= 12'b010011001111;
   6731: result <= 12'b010011001111;
   6732: result <= 12'b010011001111;
   6733: result <= 12'b010011010000;
   6734: result <= 12'b010011010000;
   6735: result <= 12'b010011010000;
   6736: result <= 12'b010011010000;
   6737: result <= 12'b010011010000;
   6738: result <= 12'b010011010000;
   6739: result <= 12'b010011010001;
   6740: result <= 12'b010011010001;
   6741: result <= 12'b010011010001;
   6742: result <= 12'b010011010001;
   6743: result <= 12'b010011010001;
   6744: result <= 12'b010011010001;
   6745: result <= 12'b010011010001;
   6746: result <= 12'b010011010010;
   6747: result <= 12'b010011010010;
   6748: result <= 12'b010011010010;
   6749: result <= 12'b010011010010;
   6750: result <= 12'b010011010010;
   6751: result <= 12'b010011010010;
   6752: result <= 12'b010011010011;
   6753: result <= 12'b010011010011;
   6754: result <= 12'b010011010011;
   6755: result <= 12'b010011010011;
   6756: result <= 12'b010011010011;
   6757: result <= 12'b010011010011;
   6758: result <= 12'b010011010100;
   6759: result <= 12'b010011010100;
   6760: result <= 12'b010011010100;
   6761: result <= 12'b010011010100;
   6762: result <= 12'b010011010100;
   6763: result <= 12'b010011010100;
   6764: result <= 12'b010011010100;
   6765: result <= 12'b010011010101;
   6766: result <= 12'b010011010101;
   6767: result <= 12'b010011010101;
   6768: result <= 12'b010011010101;
   6769: result <= 12'b010011010101;
   6770: result <= 12'b010011010101;
   6771: result <= 12'b010011010110;
   6772: result <= 12'b010011010110;
   6773: result <= 12'b010011010110;
   6774: result <= 12'b010011010110;
   6775: result <= 12'b010011010110;
   6776: result <= 12'b010011010110;
   6777: result <= 12'b010011010110;
   6778: result <= 12'b010011010111;
   6779: result <= 12'b010011010111;
   6780: result <= 12'b010011010111;
   6781: result <= 12'b010011010111;
   6782: result <= 12'b010011010111;
   6783: result <= 12'b010011010111;
   6784: result <= 12'b010011011000;
   6785: result <= 12'b010011011000;
   6786: result <= 12'b010011011000;
   6787: result <= 12'b010011011000;
   6788: result <= 12'b010011011000;
   6789: result <= 12'b010011011000;
   6790: result <= 12'b010011011001;
   6791: result <= 12'b010011011001;
   6792: result <= 12'b010011011001;
   6793: result <= 12'b010011011001;
   6794: result <= 12'b010011011001;
   6795: result <= 12'b010011011001;
   6796: result <= 12'b010011011001;
   6797: result <= 12'b010011011010;
   6798: result <= 12'b010011011010;
   6799: result <= 12'b010011011010;
   6800: result <= 12'b010011011010;
   6801: result <= 12'b010011011010;
   6802: result <= 12'b010011011010;
   6803: result <= 12'b010011011011;
   6804: result <= 12'b010011011011;
   6805: result <= 12'b010011011011;
   6806: result <= 12'b010011011011;
   6807: result <= 12'b010011011011;
   6808: result <= 12'b010011011011;
   6809: result <= 12'b010011011011;
   6810: result <= 12'b010011011100;
   6811: result <= 12'b010011011100;
   6812: result <= 12'b010011011100;
   6813: result <= 12'b010011011100;
   6814: result <= 12'b010011011100;
   6815: result <= 12'b010011011100;
   6816: result <= 12'b010011011101;
   6817: result <= 12'b010011011101;
   6818: result <= 12'b010011011101;
   6819: result <= 12'b010011011101;
   6820: result <= 12'b010011011101;
   6821: result <= 12'b010011011101;
   6822: result <= 12'b010011011110;
   6823: result <= 12'b010011011110;
   6824: result <= 12'b010011011110;
   6825: result <= 12'b010011011110;
   6826: result <= 12'b010011011110;
   6827: result <= 12'b010011011110;
   6828: result <= 12'b010011011110;
   6829: result <= 12'b010011011111;
   6830: result <= 12'b010011011111;
   6831: result <= 12'b010011011111;
   6832: result <= 12'b010011011111;
   6833: result <= 12'b010011011111;
   6834: result <= 12'b010011011111;
   6835: result <= 12'b010011100000;
   6836: result <= 12'b010011100000;
   6837: result <= 12'b010011100000;
   6838: result <= 12'b010011100000;
   6839: result <= 12'b010011100000;
   6840: result <= 12'b010011100000;
   6841: result <= 12'b010011100000;
   6842: result <= 12'b010011100001;
   6843: result <= 12'b010011100001;
   6844: result <= 12'b010011100001;
   6845: result <= 12'b010011100001;
   6846: result <= 12'b010011100001;
   6847: result <= 12'b010011100001;
   6848: result <= 12'b010011100010;
   6849: result <= 12'b010011100010;
   6850: result <= 12'b010011100010;
   6851: result <= 12'b010011100010;
   6852: result <= 12'b010011100010;
   6853: result <= 12'b010011100010;
   6854: result <= 12'b010011100010;
   6855: result <= 12'b010011100011;
   6856: result <= 12'b010011100011;
   6857: result <= 12'b010011100011;
   6858: result <= 12'b010011100011;
   6859: result <= 12'b010011100011;
   6860: result <= 12'b010011100011;
   6861: result <= 12'b010011100100;
   6862: result <= 12'b010011100100;
   6863: result <= 12'b010011100100;
   6864: result <= 12'b010011100100;
   6865: result <= 12'b010011100100;
   6866: result <= 12'b010011100100;
   6867: result <= 12'b010011100101;
   6868: result <= 12'b010011100101;
   6869: result <= 12'b010011100101;
   6870: result <= 12'b010011100101;
   6871: result <= 12'b010011100101;
   6872: result <= 12'b010011100101;
   6873: result <= 12'b010011100101;
   6874: result <= 12'b010011100110;
   6875: result <= 12'b010011100110;
   6876: result <= 12'b010011100110;
   6877: result <= 12'b010011100110;
   6878: result <= 12'b010011100110;
   6879: result <= 12'b010011100110;
   6880: result <= 12'b010011100111;
   6881: result <= 12'b010011100111;
   6882: result <= 12'b010011100111;
   6883: result <= 12'b010011100111;
   6884: result <= 12'b010011100111;
   6885: result <= 12'b010011100111;
   6886: result <= 12'b010011100111;
   6887: result <= 12'b010011101000;
   6888: result <= 12'b010011101000;
   6889: result <= 12'b010011101000;
   6890: result <= 12'b010011101000;
   6891: result <= 12'b010011101000;
   6892: result <= 12'b010011101000;
   6893: result <= 12'b010011101001;
   6894: result <= 12'b010011101001;
   6895: result <= 12'b010011101001;
   6896: result <= 12'b010011101001;
   6897: result <= 12'b010011101001;
   6898: result <= 12'b010011101001;
   6899: result <= 12'b010011101001;
   6900: result <= 12'b010011101010;
   6901: result <= 12'b010011101010;
   6902: result <= 12'b010011101010;
   6903: result <= 12'b010011101010;
   6904: result <= 12'b010011101010;
   6905: result <= 12'b010011101010;
   6906: result <= 12'b010011101011;
   6907: result <= 12'b010011101011;
   6908: result <= 12'b010011101011;
   6909: result <= 12'b010011101011;
   6910: result <= 12'b010011101011;
   6911: result <= 12'b010011101011;
   6912: result <= 12'b010011101011;
   6913: result <= 12'b010011101100;
   6914: result <= 12'b010011101100;
   6915: result <= 12'b010011101100;
   6916: result <= 12'b010011101100;
   6917: result <= 12'b010011101100;
   6918: result <= 12'b010011101100;
   6919: result <= 12'b010011101101;
   6920: result <= 12'b010011101101;
   6921: result <= 12'b010011101101;
   6922: result <= 12'b010011101101;
   6923: result <= 12'b010011101101;
   6924: result <= 12'b010011101101;
   6925: result <= 12'b010011101110;
   6926: result <= 12'b010011101110;
   6927: result <= 12'b010011101110;
   6928: result <= 12'b010011101110;
   6929: result <= 12'b010011101110;
   6930: result <= 12'b010011101110;
   6931: result <= 12'b010011101110;
   6932: result <= 12'b010011101111;
   6933: result <= 12'b010011101111;
   6934: result <= 12'b010011101111;
   6935: result <= 12'b010011101111;
   6936: result <= 12'b010011101111;
   6937: result <= 12'b010011101111;
   6938: result <= 12'b010011110000;
   6939: result <= 12'b010011110000;
   6940: result <= 12'b010011110000;
   6941: result <= 12'b010011110000;
   6942: result <= 12'b010011110000;
   6943: result <= 12'b010011110000;
   6944: result <= 12'b010011110000;
   6945: result <= 12'b010011110001;
   6946: result <= 12'b010011110001;
   6947: result <= 12'b010011110001;
   6948: result <= 12'b010011110001;
   6949: result <= 12'b010011110001;
   6950: result <= 12'b010011110001;
   6951: result <= 12'b010011110010;
   6952: result <= 12'b010011110010;
   6953: result <= 12'b010011110010;
   6954: result <= 12'b010011110010;
   6955: result <= 12'b010011110010;
   6956: result <= 12'b010011110010;
   6957: result <= 12'b010011110010;
   6958: result <= 12'b010011110011;
   6959: result <= 12'b010011110011;
   6960: result <= 12'b010011110011;
   6961: result <= 12'b010011110011;
   6962: result <= 12'b010011110011;
   6963: result <= 12'b010011110011;
   6964: result <= 12'b010011110100;
   6965: result <= 12'b010011110100;
   6966: result <= 12'b010011110100;
   6967: result <= 12'b010011110100;
   6968: result <= 12'b010011110100;
   6969: result <= 12'b010011110100;
   6970: result <= 12'b010011110100;
   6971: result <= 12'b010011110101;
   6972: result <= 12'b010011110101;
   6973: result <= 12'b010011110101;
   6974: result <= 12'b010011110101;
   6975: result <= 12'b010011110101;
   6976: result <= 12'b010011110101;
   6977: result <= 12'b010011110110;
   6978: result <= 12'b010011110110;
   6979: result <= 12'b010011110110;
   6980: result <= 12'b010011110110;
   6981: result <= 12'b010011110110;
   6982: result <= 12'b010011110110;
   6983: result <= 12'b010011110110;
   6984: result <= 12'b010011110111;
   6985: result <= 12'b010011110111;
   6986: result <= 12'b010011110111;
   6987: result <= 12'b010011110111;
   6988: result <= 12'b010011110111;
   6989: result <= 12'b010011110111;
   6990: result <= 12'b010011111000;
   6991: result <= 12'b010011111000;
   6992: result <= 12'b010011111000;
   6993: result <= 12'b010011111000;
   6994: result <= 12'b010011111000;
   6995: result <= 12'b010011111000;
   6996: result <= 12'b010011111000;
   6997: result <= 12'b010011111001;
   6998: result <= 12'b010011111001;
   6999: result <= 12'b010011111001;
   7000: result <= 12'b010011111001;
   7001: result <= 12'b010011111001;
   7002: result <= 12'b010011111001;
   7003: result <= 12'b010011111010;
   7004: result <= 12'b010011111010;
   7005: result <= 12'b010011111010;
   7006: result <= 12'b010011111010;
   7007: result <= 12'b010011111010;
   7008: result <= 12'b010011111010;
   7009: result <= 12'b010011111010;
   7010: result <= 12'b010011111011;
   7011: result <= 12'b010011111011;
   7012: result <= 12'b010011111011;
   7013: result <= 12'b010011111011;
   7014: result <= 12'b010011111011;
   7015: result <= 12'b010011111011;
   7016: result <= 12'b010011111100;
   7017: result <= 12'b010011111100;
   7018: result <= 12'b010011111100;
   7019: result <= 12'b010011111100;
   7020: result <= 12'b010011111100;
   7021: result <= 12'b010011111100;
   7022: result <= 12'b010011111100;
   7023: result <= 12'b010011111101;
   7024: result <= 12'b010011111101;
   7025: result <= 12'b010011111101;
   7026: result <= 12'b010011111101;
   7027: result <= 12'b010011111101;
   7028: result <= 12'b010011111101;
   7029: result <= 12'b010011111110;
   7030: result <= 12'b010011111110;
   7031: result <= 12'b010011111110;
   7032: result <= 12'b010011111110;
   7033: result <= 12'b010011111110;
   7034: result <= 12'b010011111110;
   7035: result <= 12'b010011111110;
   7036: result <= 12'b010011111111;
   7037: result <= 12'b010011111111;
   7038: result <= 12'b010011111111;
   7039: result <= 12'b010011111111;
   7040: result <= 12'b010011111111;
   7041: result <= 12'b010011111111;
   7042: result <= 12'b010100000000;
   7043: result <= 12'b010100000000;
   7044: result <= 12'b010100000000;
   7045: result <= 12'b010100000000;
   7046: result <= 12'b010100000000;
   7047: result <= 12'b010100000000;
   7048: result <= 12'b010100000000;
   7049: result <= 12'b010100000001;
   7050: result <= 12'b010100000001;
   7051: result <= 12'b010100000001;
   7052: result <= 12'b010100000001;
   7053: result <= 12'b010100000001;
   7054: result <= 12'b010100000001;
   7055: result <= 12'b010100000010;
   7056: result <= 12'b010100000010;
   7057: result <= 12'b010100000010;
   7058: result <= 12'b010100000010;
   7059: result <= 12'b010100000010;
   7060: result <= 12'b010100000010;
   7061: result <= 12'b010100000010;
   7062: result <= 12'b010100000011;
   7063: result <= 12'b010100000011;
   7064: result <= 12'b010100000011;
   7065: result <= 12'b010100000011;
   7066: result <= 12'b010100000011;
   7067: result <= 12'b010100000011;
   7068: result <= 12'b010100000011;
   7069: result <= 12'b010100000100;
   7070: result <= 12'b010100000100;
   7071: result <= 12'b010100000100;
   7072: result <= 12'b010100000100;
   7073: result <= 12'b010100000100;
   7074: result <= 12'b010100000100;
   7075: result <= 12'b010100000101;
   7076: result <= 12'b010100000101;
   7077: result <= 12'b010100000101;
   7078: result <= 12'b010100000101;
   7079: result <= 12'b010100000101;
   7080: result <= 12'b010100000101;
   7081: result <= 12'b010100000101;
   7082: result <= 12'b010100000110;
   7083: result <= 12'b010100000110;
   7084: result <= 12'b010100000110;
   7085: result <= 12'b010100000110;
   7086: result <= 12'b010100000110;
   7087: result <= 12'b010100000110;
   7088: result <= 12'b010100000111;
   7089: result <= 12'b010100000111;
   7090: result <= 12'b010100000111;
   7091: result <= 12'b010100000111;
   7092: result <= 12'b010100000111;
   7093: result <= 12'b010100000111;
   7094: result <= 12'b010100000111;
   7095: result <= 12'b010100001000;
   7096: result <= 12'b010100001000;
   7097: result <= 12'b010100001000;
   7098: result <= 12'b010100001000;
   7099: result <= 12'b010100001000;
   7100: result <= 12'b010100001000;
   7101: result <= 12'b010100001001;
   7102: result <= 12'b010100001001;
   7103: result <= 12'b010100001001;
   7104: result <= 12'b010100001001;
   7105: result <= 12'b010100001001;
   7106: result <= 12'b010100001001;
   7107: result <= 12'b010100001001;
   7108: result <= 12'b010100001010;
   7109: result <= 12'b010100001010;
   7110: result <= 12'b010100001010;
   7111: result <= 12'b010100001010;
   7112: result <= 12'b010100001010;
   7113: result <= 12'b010100001010;
   7114: result <= 12'b010100001011;
   7115: result <= 12'b010100001011;
   7116: result <= 12'b010100001011;
   7117: result <= 12'b010100001011;
   7118: result <= 12'b010100001011;
   7119: result <= 12'b010100001011;
   7120: result <= 12'b010100001011;
   7121: result <= 12'b010100001100;
   7122: result <= 12'b010100001100;
   7123: result <= 12'b010100001100;
   7124: result <= 12'b010100001100;
   7125: result <= 12'b010100001100;
   7126: result <= 12'b010100001100;
   7127: result <= 12'b010100001101;
   7128: result <= 12'b010100001101;
   7129: result <= 12'b010100001101;
   7130: result <= 12'b010100001101;
   7131: result <= 12'b010100001101;
   7132: result <= 12'b010100001101;
   7133: result <= 12'b010100001101;
   7134: result <= 12'b010100001110;
   7135: result <= 12'b010100001110;
   7136: result <= 12'b010100001110;
   7137: result <= 12'b010100001110;
   7138: result <= 12'b010100001110;
   7139: result <= 12'b010100001110;
   7140: result <= 12'b010100001110;
   7141: result <= 12'b010100001111;
   7142: result <= 12'b010100001111;
   7143: result <= 12'b010100001111;
   7144: result <= 12'b010100001111;
   7145: result <= 12'b010100001111;
   7146: result <= 12'b010100001111;
   7147: result <= 12'b010100010000;
   7148: result <= 12'b010100010000;
   7149: result <= 12'b010100010000;
   7150: result <= 12'b010100010000;
   7151: result <= 12'b010100010000;
   7152: result <= 12'b010100010000;
   7153: result <= 12'b010100010000;
   7154: result <= 12'b010100010001;
   7155: result <= 12'b010100010001;
   7156: result <= 12'b010100010001;
   7157: result <= 12'b010100010001;
   7158: result <= 12'b010100010001;
   7159: result <= 12'b010100010001;
   7160: result <= 12'b010100010010;
   7161: result <= 12'b010100010010;
   7162: result <= 12'b010100010010;
   7163: result <= 12'b010100010010;
   7164: result <= 12'b010100010010;
   7165: result <= 12'b010100010010;
   7166: result <= 12'b010100010010;
   7167: result <= 12'b010100010011;
   7168: result <= 12'b010100010011;
   7169: result <= 12'b010100010011;
   7170: result <= 12'b010100010011;
   7171: result <= 12'b010100010011;
   7172: result <= 12'b010100010011;
   7173: result <= 12'b010100010011;
   7174: result <= 12'b010100010100;
   7175: result <= 12'b010100010100;
   7176: result <= 12'b010100010100;
   7177: result <= 12'b010100010100;
   7178: result <= 12'b010100010100;
   7179: result <= 12'b010100010100;
   7180: result <= 12'b010100010101;
   7181: result <= 12'b010100010101;
   7182: result <= 12'b010100010101;
   7183: result <= 12'b010100010101;
   7184: result <= 12'b010100010101;
   7185: result <= 12'b010100010101;
   7186: result <= 12'b010100010101;
   7187: result <= 12'b010100010110;
   7188: result <= 12'b010100010110;
   7189: result <= 12'b010100010110;
   7190: result <= 12'b010100010110;
   7191: result <= 12'b010100010110;
   7192: result <= 12'b010100010110;
   7193: result <= 12'b010100010111;
   7194: result <= 12'b010100010111;
   7195: result <= 12'b010100010111;
   7196: result <= 12'b010100010111;
   7197: result <= 12'b010100010111;
   7198: result <= 12'b010100010111;
   7199: result <= 12'b010100010111;
   7200: result <= 12'b010100011000;
   7201: result <= 12'b010100011000;
   7202: result <= 12'b010100011000;
   7203: result <= 12'b010100011000;
   7204: result <= 12'b010100011000;
   7205: result <= 12'b010100011000;
   7206: result <= 12'b010100011000;
   7207: result <= 12'b010100011001;
   7208: result <= 12'b010100011001;
   7209: result <= 12'b010100011001;
   7210: result <= 12'b010100011001;
   7211: result <= 12'b010100011001;
   7212: result <= 12'b010100011001;
   7213: result <= 12'b010100011010;
   7214: result <= 12'b010100011010;
   7215: result <= 12'b010100011010;
   7216: result <= 12'b010100011010;
   7217: result <= 12'b010100011010;
   7218: result <= 12'b010100011010;
   7219: result <= 12'b010100011010;
   7220: result <= 12'b010100011011;
   7221: result <= 12'b010100011011;
   7222: result <= 12'b010100011011;
   7223: result <= 12'b010100011011;
   7224: result <= 12'b010100011011;
   7225: result <= 12'b010100011011;
   7226: result <= 12'b010100011100;
   7227: result <= 12'b010100011100;
   7228: result <= 12'b010100011100;
   7229: result <= 12'b010100011100;
   7230: result <= 12'b010100011100;
   7231: result <= 12'b010100011100;
   7232: result <= 12'b010100011100;
   7233: result <= 12'b010100011101;
   7234: result <= 12'b010100011101;
   7235: result <= 12'b010100011101;
   7236: result <= 12'b010100011101;
   7237: result <= 12'b010100011101;
   7238: result <= 12'b010100011101;
   7239: result <= 12'b010100011101;
   7240: result <= 12'b010100011110;
   7241: result <= 12'b010100011110;
   7242: result <= 12'b010100011110;
   7243: result <= 12'b010100011110;
   7244: result <= 12'b010100011110;
   7245: result <= 12'b010100011110;
   7246: result <= 12'b010100011111;
   7247: result <= 12'b010100011111;
   7248: result <= 12'b010100011111;
   7249: result <= 12'b010100011111;
   7250: result <= 12'b010100011111;
   7251: result <= 12'b010100011111;
   7252: result <= 12'b010100011111;
   7253: result <= 12'b010100100000;
   7254: result <= 12'b010100100000;
   7255: result <= 12'b010100100000;
   7256: result <= 12'b010100100000;
   7257: result <= 12'b010100100000;
   7258: result <= 12'b010100100000;
   7259: result <= 12'b010100100000;
   7260: result <= 12'b010100100001;
   7261: result <= 12'b010100100001;
   7262: result <= 12'b010100100001;
   7263: result <= 12'b010100100001;
   7264: result <= 12'b010100100001;
   7265: result <= 12'b010100100001;
   7266: result <= 12'b010100100010;
   7267: result <= 12'b010100100010;
   7268: result <= 12'b010100100010;
   7269: result <= 12'b010100100010;
   7270: result <= 12'b010100100010;
   7271: result <= 12'b010100100010;
   7272: result <= 12'b010100100010;
   7273: result <= 12'b010100100011;
   7274: result <= 12'b010100100011;
   7275: result <= 12'b010100100011;
   7276: result <= 12'b010100100011;
   7277: result <= 12'b010100100011;
   7278: result <= 12'b010100100011;
   7279: result <= 12'b010100100100;
   7280: result <= 12'b010100100100;
   7281: result <= 12'b010100100100;
   7282: result <= 12'b010100100100;
   7283: result <= 12'b010100100100;
   7284: result <= 12'b010100100100;
   7285: result <= 12'b010100100100;
   7286: result <= 12'b010100100101;
   7287: result <= 12'b010100100101;
   7288: result <= 12'b010100100101;
   7289: result <= 12'b010100100101;
   7290: result <= 12'b010100100101;
   7291: result <= 12'b010100100101;
   7292: result <= 12'b010100100101;
   7293: result <= 12'b010100100110;
   7294: result <= 12'b010100100110;
   7295: result <= 12'b010100100110;
   7296: result <= 12'b010100100110;
   7297: result <= 12'b010100100110;
   7298: result <= 12'b010100100110;
   7299: result <= 12'b010100100111;
   7300: result <= 12'b010100100111;
   7301: result <= 12'b010100100111;
   7302: result <= 12'b010100100111;
   7303: result <= 12'b010100100111;
   7304: result <= 12'b010100100111;
   7305: result <= 12'b010100100111;
   7306: result <= 12'b010100101000;
   7307: result <= 12'b010100101000;
   7308: result <= 12'b010100101000;
   7309: result <= 12'b010100101000;
   7310: result <= 12'b010100101000;
   7311: result <= 12'b010100101000;
   7312: result <= 12'b010100101000;
   7313: result <= 12'b010100101001;
   7314: result <= 12'b010100101001;
   7315: result <= 12'b010100101001;
   7316: result <= 12'b010100101001;
   7317: result <= 12'b010100101001;
   7318: result <= 12'b010100101001;
   7319: result <= 12'b010100101010;
   7320: result <= 12'b010100101010;
   7321: result <= 12'b010100101010;
   7322: result <= 12'b010100101010;
   7323: result <= 12'b010100101010;
   7324: result <= 12'b010100101010;
   7325: result <= 12'b010100101010;
   7326: result <= 12'b010100101011;
   7327: result <= 12'b010100101011;
   7328: result <= 12'b010100101011;
   7329: result <= 12'b010100101011;
   7330: result <= 12'b010100101011;
   7331: result <= 12'b010100101011;
   7332: result <= 12'b010100101011;
   7333: result <= 12'b010100101100;
   7334: result <= 12'b010100101100;
   7335: result <= 12'b010100101100;
   7336: result <= 12'b010100101100;
   7337: result <= 12'b010100101100;
   7338: result <= 12'b010100101100;
   7339: result <= 12'b010100101101;
   7340: result <= 12'b010100101101;
   7341: result <= 12'b010100101101;
   7342: result <= 12'b010100101101;
   7343: result <= 12'b010100101101;
   7344: result <= 12'b010100101101;
   7345: result <= 12'b010100101101;
   7346: result <= 12'b010100101110;
   7347: result <= 12'b010100101110;
   7348: result <= 12'b010100101110;
   7349: result <= 12'b010100101110;
   7350: result <= 12'b010100101110;
   7351: result <= 12'b010100101110;
   7352: result <= 12'b010100101110;
   7353: result <= 12'b010100101111;
   7354: result <= 12'b010100101111;
   7355: result <= 12'b010100101111;
   7356: result <= 12'b010100101111;
   7357: result <= 12'b010100101111;
   7358: result <= 12'b010100101111;
   7359: result <= 12'b010100110000;
   7360: result <= 12'b010100110000;
   7361: result <= 12'b010100110000;
   7362: result <= 12'b010100110000;
   7363: result <= 12'b010100110000;
   7364: result <= 12'b010100110000;
   7365: result <= 12'b010100110000;
   7366: result <= 12'b010100110001;
   7367: result <= 12'b010100110001;
   7368: result <= 12'b010100110001;
   7369: result <= 12'b010100110001;
   7370: result <= 12'b010100110001;
   7371: result <= 12'b010100110001;
   7372: result <= 12'b010100110001;
   7373: result <= 12'b010100110010;
   7374: result <= 12'b010100110010;
   7375: result <= 12'b010100110010;
   7376: result <= 12'b010100110010;
   7377: result <= 12'b010100110010;
   7378: result <= 12'b010100110010;
   7379: result <= 12'b010100110010;
   7380: result <= 12'b010100110011;
   7381: result <= 12'b010100110011;
   7382: result <= 12'b010100110011;
   7383: result <= 12'b010100110011;
   7384: result <= 12'b010100110011;
   7385: result <= 12'b010100110011;
   7386: result <= 12'b010100110100;
   7387: result <= 12'b010100110100;
   7388: result <= 12'b010100110100;
   7389: result <= 12'b010100110100;
   7390: result <= 12'b010100110100;
   7391: result <= 12'b010100110100;
   7392: result <= 12'b010100110100;
   7393: result <= 12'b010100110101;
   7394: result <= 12'b010100110101;
   7395: result <= 12'b010100110101;
   7396: result <= 12'b010100110101;
   7397: result <= 12'b010100110101;
   7398: result <= 12'b010100110101;
   7399: result <= 12'b010100110101;
   7400: result <= 12'b010100110110;
   7401: result <= 12'b010100110110;
   7402: result <= 12'b010100110110;
   7403: result <= 12'b010100110110;
   7404: result <= 12'b010100110110;
   7405: result <= 12'b010100110110;
   7406: result <= 12'b010100110111;
   7407: result <= 12'b010100110111;
   7408: result <= 12'b010100110111;
   7409: result <= 12'b010100110111;
   7410: result <= 12'b010100110111;
   7411: result <= 12'b010100110111;
   7412: result <= 12'b010100110111;
   7413: result <= 12'b010100111000;
   7414: result <= 12'b010100111000;
   7415: result <= 12'b010100111000;
   7416: result <= 12'b010100111000;
   7417: result <= 12'b010100111000;
   7418: result <= 12'b010100111000;
   7419: result <= 12'b010100111000;
   7420: result <= 12'b010100111001;
   7421: result <= 12'b010100111001;
   7422: result <= 12'b010100111001;
   7423: result <= 12'b010100111001;
   7424: result <= 12'b010100111001;
   7425: result <= 12'b010100111001;
   7426: result <= 12'b010100111001;
   7427: result <= 12'b010100111010;
   7428: result <= 12'b010100111010;
   7429: result <= 12'b010100111010;
   7430: result <= 12'b010100111010;
   7431: result <= 12'b010100111010;
   7432: result <= 12'b010100111010;
   7433: result <= 12'b010100111011;
   7434: result <= 12'b010100111011;
   7435: result <= 12'b010100111011;
   7436: result <= 12'b010100111011;
   7437: result <= 12'b010100111011;
   7438: result <= 12'b010100111011;
   7439: result <= 12'b010100111011;
   7440: result <= 12'b010100111100;
   7441: result <= 12'b010100111100;
   7442: result <= 12'b010100111100;
   7443: result <= 12'b010100111100;
   7444: result <= 12'b010100111100;
   7445: result <= 12'b010100111100;
   7446: result <= 12'b010100111100;
   7447: result <= 12'b010100111101;
   7448: result <= 12'b010100111101;
   7449: result <= 12'b010100111101;
   7450: result <= 12'b010100111101;
   7451: result <= 12'b010100111101;
   7452: result <= 12'b010100111101;
   7453: result <= 12'b010100111110;
   7454: result <= 12'b010100111110;
   7455: result <= 12'b010100111110;
   7456: result <= 12'b010100111110;
   7457: result <= 12'b010100111110;
   7458: result <= 12'b010100111110;
   7459: result <= 12'b010100111110;
   7460: result <= 12'b010100111111;
   7461: result <= 12'b010100111111;
   7462: result <= 12'b010100111111;
   7463: result <= 12'b010100111111;
   7464: result <= 12'b010100111111;
   7465: result <= 12'b010100111111;
   7466: result <= 12'b010100111111;
   7467: result <= 12'b010101000000;
   7468: result <= 12'b010101000000;
   7469: result <= 12'b010101000000;
   7470: result <= 12'b010101000000;
   7471: result <= 12'b010101000000;
   7472: result <= 12'b010101000000;
   7473: result <= 12'b010101000000;
   7474: result <= 12'b010101000001;
   7475: result <= 12'b010101000001;
   7476: result <= 12'b010101000001;
   7477: result <= 12'b010101000001;
   7478: result <= 12'b010101000001;
   7479: result <= 12'b010101000001;
   7480: result <= 12'b010101000010;
   7481: result <= 12'b010101000010;
   7482: result <= 12'b010101000010;
   7483: result <= 12'b010101000010;
   7484: result <= 12'b010101000010;
   7485: result <= 12'b010101000010;
   7486: result <= 12'b010101000010;
   7487: result <= 12'b010101000011;
   7488: result <= 12'b010101000011;
   7489: result <= 12'b010101000011;
   7490: result <= 12'b010101000011;
   7491: result <= 12'b010101000011;
   7492: result <= 12'b010101000011;
   7493: result <= 12'b010101000011;
   7494: result <= 12'b010101000100;
   7495: result <= 12'b010101000100;
   7496: result <= 12'b010101000100;
   7497: result <= 12'b010101000100;
   7498: result <= 12'b010101000100;
   7499: result <= 12'b010101000100;
   7500: result <= 12'b010101000100;
   7501: result <= 12'b010101000101;
   7502: result <= 12'b010101000101;
   7503: result <= 12'b010101000101;
   7504: result <= 12'b010101000101;
   7505: result <= 12'b010101000101;
   7506: result <= 12'b010101000101;
   7507: result <= 12'b010101000101;
   7508: result <= 12'b010101000110;
   7509: result <= 12'b010101000110;
   7510: result <= 12'b010101000110;
   7511: result <= 12'b010101000110;
   7512: result <= 12'b010101000110;
   7513: result <= 12'b010101000110;
   7514: result <= 12'b010101000111;
   7515: result <= 12'b010101000111;
   7516: result <= 12'b010101000111;
   7517: result <= 12'b010101000111;
   7518: result <= 12'b010101000111;
   7519: result <= 12'b010101000111;
   7520: result <= 12'b010101000111;
   7521: result <= 12'b010101001000;
   7522: result <= 12'b010101001000;
   7523: result <= 12'b010101001000;
   7524: result <= 12'b010101001000;
   7525: result <= 12'b010101001000;
   7526: result <= 12'b010101001000;
   7527: result <= 12'b010101001000;
   7528: result <= 12'b010101001001;
   7529: result <= 12'b010101001001;
   7530: result <= 12'b010101001001;
   7531: result <= 12'b010101001001;
   7532: result <= 12'b010101001001;
   7533: result <= 12'b010101001001;
   7534: result <= 12'b010101001001;
   7535: result <= 12'b010101001010;
   7536: result <= 12'b010101001010;
   7537: result <= 12'b010101001010;
   7538: result <= 12'b010101001010;
   7539: result <= 12'b010101001010;
   7540: result <= 12'b010101001010;
   7541: result <= 12'b010101001011;
   7542: result <= 12'b010101001011;
   7543: result <= 12'b010101001011;
   7544: result <= 12'b010101001011;
   7545: result <= 12'b010101001011;
   7546: result <= 12'b010101001011;
   7547: result <= 12'b010101001011;
   7548: result <= 12'b010101001100;
   7549: result <= 12'b010101001100;
   7550: result <= 12'b010101001100;
   7551: result <= 12'b010101001100;
   7552: result <= 12'b010101001100;
   7553: result <= 12'b010101001100;
   7554: result <= 12'b010101001100;
   7555: result <= 12'b010101001101;
   7556: result <= 12'b010101001101;
   7557: result <= 12'b010101001101;
   7558: result <= 12'b010101001101;
   7559: result <= 12'b010101001101;
   7560: result <= 12'b010101001101;
   7561: result <= 12'b010101001101;
   7562: result <= 12'b010101001110;
   7563: result <= 12'b010101001110;
   7564: result <= 12'b010101001110;
   7565: result <= 12'b010101001110;
   7566: result <= 12'b010101001110;
   7567: result <= 12'b010101001110;
   7568: result <= 12'b010101001110;
   7569: result <= 12'b010101001111;
   7570: result <= 12'b010101001111;
   7571: result <= 12'b010101001111;
   7572: result <= 12'b010101001111;
   7573: result <= 12'b010101001111;
   7574: result <= 12'b010101001111;
   7575: result <= 12'b010101010000;
   7576: result <= 12'b010101010000;
   7577: result <= 12'b010101010000;
   7578: result <= 12'b010101010000;
   7579: result <= 12'b010101010000;
   7580: result <= 12'b010101010000;
   7581: result <= 12'b010101010000;
   7582: result <= 12'b010101010001;
   7583: result <= 12'b010101010001;
   7584: result <= 12'b010101010001;
   7585: result <= 12'b010101010001;
   7586: result <= 12'b010101010001;
   7587: result <= 12'b010101010001;
   7588: result <= 12'b010101010001;
   7589: result <= 12'b010101010010;
   7590: result <= 12'b010101010010;
   7591: result <= 12'b010101010010;
   7592: result <= 12'b010101010010;
   7593: result <= 12'b010101010010;
   7594: result <= 12'b010101010010;
   7595: result <= 12'b010101010010;
   7596: result <= 12'b010101010011;
   7597: result <= 12'b010101010011;
   7598: result <= 12'b010101010011;
   7599: result <= 12'b010101010011;
   7600: result <= 12'b010101010011;
   7601: result <= 12'b010101010011;
   7602: result <= 12'b010101010011;
   7603: result <= 12'b010101010100;
   7604: result <= 12'b010101010100;
   7605: result <= 12'b010101010100;
   7606: result <= 12'b010101010100;
   7607: result <= 12'b010101010100;
   7608: result <= 12'b010101010100;
   7609: result <= 12'b010101010100;
   7610: result <= 12'b010101010101;
   7611: result <= 12'b010101010101;
   7612: result <= 12'b010101010101;
   7613: result <= 12'b010101010101;
   7614: result <= 12'b010101010101;
   7615: result <= 12'b010101010101;
   7616: result <= 12'b010101010110;
   7617: result <= 12'b010101010110;
   7618: result <= 12'b010101010110;
   7619: result <= 12'b010101010110;
   7620: result <= 12'b010101010110;
   7621: result <= 12'b010101010110;
   7622: result <= 12'b010101010110;
   7623: result <= 12'b010101010111;
   7624: result <= 12'b010101010111;
   7625: result <= 12'b010101010111;
   7626: result <= 12'b010101010111;
   7627: result <= 12'b010101010111;
   7628: result <= 12'b010101010111;
   7629: result <= 12'b010101010111;
   7630: result <= 12'b010101011000;
   7631: result <= 12'b010101011000;
   7632: result <= 12'b010101011000;
   7633: result <= 12'b010101011000;
   7634: result <= 12'b010101011000;
   7635: result <= 12'b010101011000;
   7636: result <= 12'b010101011000;
   7637: result <= 12'b010101011001;
   7638: result <= 12'b010101011001;
   7639: result <= 12'b010101011001;
   7640: result <= 12'b010101011001;
   7641: result <= 12'b010101011001;
   7642: result <= 12'b010101011001;
   7643: result <= 12'b010101011001;
   7644: result <= 12'b010101011010;
   7645: result <= 12'b010101011010;
   7646: result <= 12'b010101011010;
   7647: result <= 12'b010101011010;
   7648: result <= 12'b010101011010;
   7649: result <= 12'b010101011010;
   7650: result <= 12'b010101011010;
   7651: result <= 12'b010101011011;
   7652: result <= 12'b010101011011;
   7653: result <= 12'b010101011011;
   7654: result <= 12'b010101011011;
   7655: result <= 12'b010101011011;
   7656: result <= 12'b010101011011;
   7657: result <= 12'b010101011100;
   7658: result <= 12'b010101011100;
   7659: result <= 12'b010101011100;
   7660: result <= 12'b010101011100;
   7661: result <= 12'b010101011100;
   7662: result <= 12'b010101011100;
   7663: result <= 12'b010101011100;
   7664: result <= 12'b010101011101;
   7665: result <= 12'b010101011101;
   7666: result <= 12'b010101011101;
   7667: result <= 12'b010101011101;
   7668: result <= 12'b010101011101;
   7669: result <= 12'b010101011101;
   7670: result <= 12'b010101011101;
   7671: result <= 12'b010101011110;
   7672: result <= 12'b010101011110;
   7673: result <= 12'b010101011110;
   7674: result <= 12'b010101011110;
   7675: result <= 12'b010101011110;
   7676: result <= 12'b010101011110;
   7677: result <= 12'b010101011110;
   7678: result <= 12'b010101011111;
   7679: result <= 12'b010101011111;
   7680: result <= 12'b010101011111;
   7681: result <= 12'b010101011111;
   7682: result <= 12'b010101011111;
   7683: result <= 12'b010101011111;
   7684: result <= 12'b010101011111;
   7685: result <= 12'b010101100000;
   7686: result <= 12'b010101100000;
   7687: result <= 12'b010101100000;
   7688: result <= 12'b010101100000;
   7689: result <= 12'b010101100000;
   7690: result <= 12'b010101100000;
   7691: result <= 12'b010101100000;
   7692: result <= 12'b010101100001;
   7693: result <= 12'b010101100001;
   7694: result <= 12'b010101100001;
   7695: result <= 12'b010101100001;
   7696: result <= 12'b010101100001;
   7697: result <= 12'b010101100001;
   7698: result <= 12'b010101100001;
   7699: result <= 12'b010101100010;
   7700: result <= 12'b010101100010;
   7701: result <= 12'b010101100010;
   7702: result <= 12'b010101100010;
   7703: result <= 12'b010101100010;
   7704: result <= 12'b010101100010;
   7705: result <= 12'b010101100010;
   7706: result <= 12'b010101100011;
   7707: result <= 12'b010101100011;
   7708: result <= 12'b010101100011;
   7709: result <= 12'b010101100011;
   7710: result <= 12'b010101100011;
   7711: result <= 12'b010101100011;
   7712: result <= 12'b010101100100;
   7713: result <= 12'b010101100100;
   7714: result <= 12'b010101100100;
   7715: result <= 12'b010101100100;
   7716: result <= 12'b010101100100;
   7717: result <= 12'b010101100100;
   7718: result <= 12'b010101100100;
   7719: result <= 12'b010101100101;
   7720: result <= 12'b010101100101;
   7721: result <= 12'b010101100101;
   7722: result <= 12'b010101100101;
   7723: result <= 12'b010101100101;
   7724: result <= 12'b010101100101;
   7725: result <= 12'b010101100101;
   7726: result <= 12'b010101100110;
   7727: result <= 12'b010101100110;
   7728: result <= 12'b010101100110;
   7729: result <= 12'b010101100110;
   7730: result <= 12'b010101100110;
   7731: result <= 12'b010101100110;
   7732: result <= 12'b010101100110;
   7733: result <= 12'b010101100111;
   7734: result <= 12'b010101100111;
   7735: result <= 12'b010101100111;
   7736: result <= 12'b010101100111;
   7737: result <= 12'b010101100111;
   7738: result <= 12'b010101100111;
   7739: result <= 12'b010101100111;
   7740: result <= 12'b010101101000;
   7741: result <= 12'b010101101000;
   7742: result <= 12'b010101101000;
   7743: result <= 12'b010101101000;
   7744: result <= 12'b010101101000;
   7745: result <= 12'b010101101000;
   7746: result <= 12'b010101101000;
   7747: result <= 12'b010101101001;
   7748: result <= 12'b010101101001;
   7749: result <= 12'b010101101001;
   7750: result <= 12'b010101101001;
   7751: result <= 12'b010101101001;
   7752: result <= 12'b010101101001;
   7753: result <= 12'b010101101001;
   7754: result <= 12'b010101101010;
   7755: result <= 12'b010101101010;
   7756: result <= 12'b010101101010;
   7757: result <= 12'b010101101010;
   7758: result <= 12'b010101101010;
   7759: result <= 12'b010101101010;
   7760: result <= 12'b010101101010;
   7761: result <= 12'b010101101011;
   7762: result <= 12'b010101101011;
   7763: result <= 12'b010101101011;
   7764: result <= 12'b010101101011;
   7765: result <= 12'b010101101011;
   7766: result <= 12'b010101101011;
   7767: result <= 12'b010101101011;
   7768: result <= 12'b010101101100;
   7769: result <= 12'b010101101100;
   7770: result <= 12'b010101101100;
   7771: result <= 12'b010101101100;
   7772: result <= 12'b010101101100;
   7773: result <= 12'b010101101100;
   7774: result <= 12'b010101101100;
   7775: result <= 12'b010101101101;
   7776: result <= 12'b010101101101;
   7777: result <= 12'b010101101101;
   7778: result <= 12'b010101101101;
   7779: result <= 12'b010101101101;
   7780: result <= 12'b010101101101;
   7781: result <= 12'b010101101101;
   7782: result <= 12'b010101101110;
   7783: result <= 12'b010101101110;
   7784: result <= 12'b010101101110;
   7785: result <= 12'b010101101110;
   7786: result <= 12'b010101101110;
   7787: result <= 12'b010101101110;
   7788: result <= 12'b010101101110;
   7789: result <= 12'b010101101111;
   7790: result <= 12'b010101101111;
   7791: result <= 12'b010101101111;
   7792: result <= 12'b010101101111;
   7793: result <= 12'b010101101111;
   7794: result <= 12'b010101101111;
   7795: result <= 12'b010101101111;
   7796: result <= 12'b010101110000;
   7797: result <= 12'b010101110000;
   7798: result <= 12'b010101110000;
   7799: result <= 12'b010101110000;
   7800: result <= 12'b010101110000;
   7801: result <= 12'b010101110000;
   7802: result <= 12'b010101110001;
   7803: result <= 12'b010101110001;
   7804: result <= 12'b010101110001;
   7805: result <= 12'b010101110001;
   7806: result <= 12'b010101110001;
   7807: result <= 12'b010101110001;
   7808: result <= 12'b010101110001;
   7809: result <= 12'b010101110010;
   7810: result <= 12'b010101110010;
   7811: result <= 12'b010101110010;
   7812: result <= 12'b010101110010;
   7813: result <= 12'b010101110010;
   7814: result <= 12'b010101110010;
   7815: result <= 12'b010101110010;
   7816: result <= 12'b010101110011;
   7817: result <= 12'b010101110011;
   7818: result <= 12'b010101110011;
   7819: result <= 12'b010101110011;
   7820: result <= 12'b010101110011;
   7821: result <= 12'b010101110011;
   7822: result <= 12'b010101110011;
   7823: result <= 12'b010101110100;
   7824: result <= 12'b010101110100;
   7825: result <= 12'b010101110100;
   7826: result <= 12'b010101110100;
   7827: result <= 12'b010101110100;
   7828: result <= 12'b010101110100;
   7829: result <= 12'b010101110100;
   7830: result <= 12'b010101110101;
   7831: result <= 12'b010101110101;
   7832: result <= 12'b010101110101;
   7833: result <= 12'b010101110101;
   7834: result <= 12'b010101110101;
   7835: result <= 12'b010101110101;
   7836: result <= 12'b010101110101;
   7837: result <= 12'b010101110110;
   7838: result <= 12'b010101110110;
   7839: result <= 12'b010101110110;
   7840: result <= 12'b010101110110;
   7841: result <= 12'b010101110110;
   7842: result <= 12'b010101110110;
   7843: result <= 12'b010101110110;
   7844: result <= 12'b010101110111;
   7845: result <= 12'b010101110111;
   7846: result <= 12'b010101110111;
   7847: result <= 12'b010101110111;
   7848: result <= 12'b010101110111;
   7849: result <= 12'b010101110111;
   7850: result <= 12'b010101110111;
   7851: result <= 12'b010101111000;
   7852: result <= 12'b010101111000;
   7853: result <= 12'b010101111000;
   7854: result <= 12'b010101111000;
   7855: result <= 12'b010101111000;
   7856: result <= 12'b010101111000;
   7857: result <= 12'b010101111000;
   7858: result <= 12'b010101111001;
   7859: result <= 12'b010101111001;
   7860: result <= 12'b010101111001;
   7861: result <= 12'b010101111001;
   7862: result <= 12'b010101111001;
   7863: result <= 12'b010101111001;
   7864: result <= 12'b010101111001;
   7865: result <= 12'b010101111010;
   7866: result <= 12'b010101111010;
   7867: result <= 12'b010101111010;
   7868: result <= 12'b010101111010;
   7869: result <= 12'b010101111010;
   7870: result <= 12'b010101111010;
   7871: result <= 12'b010101111010;
   7872: result <= 12'b010101111011;
   7873: result <= 12'b010101111011;
   7874: result <= 12'b010101111011;
   7875: result <= 12'b010101111011;
   7876: result <= 12'b010101111011;
   7877: result <= 12'b010101111011;
   7878: result <= 12'b010101111011;
   7879: result <= 12'b010101111100;
   7880: result <= 12'b010101111100;
   7881: result <= 12'b010101111100;
   7882: result <= 12'b010101111100;
   7883: result <= 12'b010101111100;
   7884: result <= 12'b010101111100;
   7885: result <= 12'b010101111100;
   7886: result <= 12'b010101111101;
   7887: result <= 12'b010101111101;
   7888: result <= 12'b010101111101;
   7889: result <= 12'b010101111101;
   7890: result <= 12'b010101111101;
   7891: result <= 12'b010101111101;
   7892: result <= 12'b010101111101;
   7893: result <= 12'b010101111110;
   7894: result <= 12'b010101111110;
   7895: result <= 12'b010101111110;
   7896: result <= 12'b010101111110;
   7897: result <= 12'b010101111110;
   7898: result <= 12'b010101111110;
   7899: result <= 12'b010101111110;
   7900: result <= 12'b010101111111;
   7901: result <= 12'b010101111111;
   7902: result <= 12'b010101111111;
   7903: result <= 12'b010101111111;
   7904: result <= 12'b010101111111;
   7905: result <= 12'b010101111111;
   7906: result <= 12'b010101111111;
   7907: result <= 12'b010110000000;
   7908: result <= 12'b010110000000;
   7909: result <= 12'b010110000000;
   7910: result <= 12'b010110000000;
   7911: result <= 12'b010110000000;
   7912: result <= 12'b010110000000;
   7913: result <= 12'b010110000000;
   7914: result <= 12'b010110000001;
   7915: result <= 12'b010110000001;
   7916: result <= 12'b010110000001;
   7917: result <= 12'b010110000001;
   7918: result <= 12'b010110000001;
   7919: result <= 12'b010110000001;
   7920: result <= 12'b010110000001;
   7921: result <= 12'b010110000010;
   7922: result <= 12'b010110000010;
   7923: result <= 12'b010110000010;
   7924: result <= 12'b010110000010;
   7925: result <= 12'b010110000010;
   7926: result <= 12'b010110000010;
   7927: result <= 12'b010110000010;
   7928: result <= 12'b010110000011;
   7929: result <= 12'b010110000011;
   7930: result <= 12'b010110000011;
   7931: result <= 12'b010110000011;
   7932: result <= 12'b010110000011;
   7933: result <= 12'b010110000011;
   7934: result <= 12'b010110000011;
   7935: result <= 12'b010110000100;
   7936: result <= 12'b010110000100;
   7937: result <= 12'b010110000100;
   7938: result <= 12'b010110000100;
   7939: result <= 12'b010110000100;
   7940: result <= 12'b010110000100;
   7941: result <= 12'b010110000100;
   7942: result <= 12'b010110000101;
   7943: result <= 12'b010110000101;
   7944: result <= 12'b010110000101;
   7945: result <= 12'b010110000101;
   7946: result <= 12'b010110000101;
   7947: result <= 12'b010110000101;
   7948: result <= 12'b010110000101;
   7949: result <= 12'b010110000110;
   7950: result <= 12'b010110000110;
   7951: result <= 12'b010110000110;
   7952: result <= 12'b010110000110;
   7953: result <= 12'b010110000110;
   7954: result <= 12'b010110000110;
   7955: result <= 12'b010110000110;
   7956: result <= 12'b010110000111;
   7957: result <= 12'b010110000111;
   7958: result <= 12'b010110000111;
   7959: result <= 12'b010110000111;
   7960: result <= 12'b010110000111;
   7961: result <= 12'b010110000111;
   7962: result <= 12'b010110000111;
   7963: result <= 12'b010110001000;
   7964: result <= 12'b010110001000;
   7965: result <= 12'b010110001000;
   7966: result <= 12'b010110001000;
   7967: result <= 12'b010110001000;
   7968: result <= 12'b010110001000;
   7969: result <= 12'b010110001000;
   7970: result <= 12'b010110001001;
   7971: result <= 12'b010110001001;
   7972: result <= 12'b010110001001;
   7973: result <= 12'b010110001001;
   7974: result <= 12'b010110001001;
   7975: result <= 12'b010110001001;
   7976: result <= 12'b010110001001;
   7977: result <= 12'b010110001001;
   7978: result <= 12'b010110001010;
   7979: result <= 12'b010110001010;
   7980: result <= 12'b010110001010;
   7981: result <= 12'b010110001010;
   7982: result <= 12'b010110001010;
   7983: result <= 12'b010110001010;
   7984: result <= 12'b010110001010;
   7985: result <= 12'b010110001011;
   7986: result <= 12'b010110001011;
   7987: result <= 12'b010110001011;
   7988: result <= 12'b010110001011;
   7989: result <= 12'b010110001011;
   7990: result <= 12'b010110001011;
   7991: result <= 12'b010110001011;
   7992: result <= 12'b010110001100;
   7993: result <= 12'b010110001100;
   7994: result <= 12'b010110001100;
   7995: result <= 12'b010110001100;
   7996: result <= 12'b010110001100;
   7997: result <= 12'b010110001100;
   7998: result <= 12'b010110001100;
   7999: result <= 12'b010110001101;
   8000: result <= 12'b010110001101;
   8001: result <= 12'b010110001101;
   8002: result <= 12'b010110001101;
   8003: result <= 12'b010110001101;
   8004: result <= 12'b010110001101;
   8005: result <= 12'b010110001101;
   8006: result <= 12'b010110001110;
   8007: result <= 12'b010110001110;
   8008: result <= 12'b010110001110;
   8009: result <= 12'b010110001110;
   8010: result <= 12'b010110001110;
   8011: result <= 12'b010110001110;
   8012: result <= 12'b010110001110;
   8013: result <= 12'b010110001111;
   8014: result <= 12'b010110001111;
   8015: result <= 12'b010110001111;
   8016: result <= 12'b010110001111;
   8017: result <= 12'b010110001111;
   8018: result <= 12'b010110001111;
   8019: result <= 12'b010110001111;
   8020: result <= 12'b010110010000;
   8021: result <= 12'b010110010000;
   8022: result <= 12'b010110010000;
   8023: result <= 12'b010110010000;
   8024: result <= 12'b010110010000;
   8025: result <= 12'b010110010000;
   8026: result <= 12'b010110010000;
   8027: result <= 12'b010110010001;
   8028: result <= 12'b010110010001;
   8029: result <= 12'b010110010001;
   8030: result <= 12'b010110010001;
   8031: result <= 12'b010110010001;
   8032: result <= 12'b010110010001;
   8033: result <= 12'b010110010001;
   8034: result <= 12'b010110010010;
   8035: result <= 12'b010110010010;
   8036: result <= 12'b010110010010;
   8037: result <= 12'b010110010010;
   8038: result <= 12'b010110010010;
   8039: result <= 12'b010110010010;
   8040: result <= 12'b010110010010;
   8041: result <= 12'b010110010011;
   8042: result <= 12'b010110010011;
   8043: result <= 12'b010110010011;
   8044: result <= 12'b010110010011;
   8045: result <= 12'b010110010011;
   8046: result <= 12'b010110010011;
   8047: result <= 12'b010110010011;
   8048: result <= 12'b010110010100;
   8049: result <= 12'b010110010100;
   8050: result <= 12'b010110010100;
   8051: result <= 12'b010110010100;
   8052: result <= 12'b010110010100;
   8053: result <= 12'b010110010100;
   8054: result <= 12'b010110010100;
   8055: result <= 12'b010110010101;
   8056: result <= 12'b010110010101;
   8057: result <= 12'b010110010101;
   8058: result <= 12'b010110010101;
   8059: result <= 12'b010110010101;
   8060: result <= 12'b010110010101;
   8061: result <= 12'b010110010101;
   8062: result <= 12'b010110010101;
   8063: result <= 12'b010110010110;
   8064: result <= 12'b010110010110;
   8065: result <= 12'b010110010110;
   8066: result <= 12'b010110010110;
   8067: result <= 12'b010110010110;
   8068: result <= 12'b010110010110;
   8069: result <= 12'b010110010110;
   8070: result <= 12'b010110010111;
   8071: result <= 12'b010110010111;
   8072: result <= 12'b010110010111;
   8073: result <= 12'b010110010111;
   8074: result <= 12'b010110010111;
   8075: result <= 12'b010110010111;
   8076: result <= 12'b010110010111;
   8077: result <= 12'b010110011000;
   8078: result <= 12'b010110011000;
   8079: result <= 12'b010110011000;
   8080: result <= 12'b010110011000;
   8081: result <= 12'b010110011000;
   8082: result <= 12'b010110011000;
   8083: result <= 12'b010110011000;
   8084: result <= 12'b010110011001;
   8085: result <= 12'b010110011001;
   8086: result <= 12'b010110011001;
   8087: result <= 12'b010110011001;
   8088: result <= 12'b010110011001;
   8089: result <= 12'b010110011001;
   8090: result <= 12'b010110011001;
   8091: result <= 12'b010110011010;
   8092: result <= 12'b010110011010;
   8093: result <= 12'b010110011010;
   8094: result <= 12'b010110011010;
   8095: result <= 12'b010110011010;
   8096: result <= 12'b010110011010;
   8097: result <= 12'b010110011010;
   8098: result <= 12'b010110011011;
   8099: result <= 12'b010110011011;
   8100: result <= 12'b010110011011;
   8101: result <= 12'b010110011011;
   8102: result <= 12'b010110011011;
   8103: result <= 12'b010110011011;
   8104: result <= 12'b010110011011;
   8105: result <= 12'b010110011100;
   8106: result <= 12'b010110011100;
   8107: result <= 12'b010110011100;
   8108: result <= 12'b010110011100;
   8109: result <= 12'b010110011100;
   8110: result <= 12'b010110011100;
   8111: result <= 12'b010110011100;
   8112: result <= 12'b010110011101;
   8113: result <= 12'b010110011101;
   8114: result <= 12'b010110011101;
   8115: result <= 12'b010110011101;
   8116: result <= 12'b010110011101;
   8117: result <= 12'b010110011101;
   8118: result <= 12'b010110011101;
   8119: result <= 12'b010110011101;
   8120: result <= 12'b010110011110;
   8121: result <= 12'b010110011110;
   8122: result <= 12'b010110011110;
   8123: result <= 12'b010110011110;
   8124: result <= 12'b010110011110;
   8125: result <= 12'b010110011110;
   8126: result <= 12'b010110011110;
   8127: result <= 12'b010110011111;
   8128: result <= 12'b010110011111;
   8129: result <= 12'b010110011111;
   8130: result <= 12'b010110011111;
   8131: result <= 12'b010110011111;
   8132: result <= 12'b010110011111;
   8133: result <= 12'b010110011111;
   8134: result <= 12'b010110100000;
   8135: result <= 12'b010110100000;
   8136: result <= 12'b010110100000;
   8137: result <= 12'b010110100000;
   8138: result <= 12'b010110100000;
   8139: result <= 12'b010110100000;
   8140: result <= 12'b010110100000;
   8141: result <= 12'b010110100001;
   8142: result <= 12'b010110100001;
   8143: result <= 12'b010110100001;
   8144: result <= 12'b010110100001;
   8145: result <= 12'b010110100001;
   8146: result <= 12'b010110100001;
   8147: result <= 12'b010110100001;
   8148: result <= 12'b010110100010;
   8149: result <= 12'b010110100010;
   8150: result <= 12'b010110100010;
   8151: result <= 12'b010110100010;
   8152: result <= 12'b010110100010;
   8153: result <= 12'b010110100010;
   8154: result <= 12'b010110100010;
   8155: result <= 12'b010110100011;
   8156: result <= 12'b010110100011;
   8157: result <= 12'b010110100011;
   8158: result <= 12'b010110100011;
   8159: result <= 12'b010110100011;
   8160: result <= 12'b010110100011;
   8161: result <= 12'b010110100011;
   8162: result <= 12'b010110100011;
   8163: result <= 12'b010110100100;
   8164: result <= 12'b010110100100;
   8165: result <= 12'b010110100100;
   8166: result <= 12'b010110100100;
   8167: result <= 12'b010110100100;
   8168: result <= 12'b010110100100;
   8169: result <= 12'b010110100100;
   8170: result <= 12'b010110100101;
   8171: result <= 12'b010110100101;
   8172: result <= 12'b010110100101;
   8173: result <= 12'b010110100101;
   8174: result <= 12'b010110100101;
   8175: result <= 12'b010110100101;
   8176: result <= 12'b010110100101;
   8177: result <= 12'b010110100110;
   8178: result <= 12'b010110100110;
   8179: result <= 12'b010110100110;
   8180: result <= 12'b010110100110;
   8181: result <= 12'b010110100110;
   8182: result <= 12'b010110100110;
   8183: result <= 12'b010110100110;
   8184: result <= 12'b010110100111;
   8185: result <= 12'b010110100111;
   8186: result <= 12'b010110100111;
   8187: result <= 12'b010110100111;
   8188: result <= 12'b010110100111;
   8189: result <= 12'b010110100111;
   8190: result <= 12'b010110100111;
   8191: result <= 12'b010110101000;
   8192: result <= 12'b010110101000;
   8193: result <= 12'b010110101000;
   8194: result <= 12'b010110101000;
   8195: result <= 12'b010110101000;
   8196: result <= 12'b010110101000;
   8197: result <= 12'b010110101000;
   8198: result <= 12'b010110101000;
   8199: result <= 12'b010110101001;
   8200: result <= 12'b010110101001;
   8201: result <= 12'b010110101001;
   8202: result <= 12'b010110101001;
   8203: result <= 12'b010110101001;
   8204: result <= 12'b010110101001;
   8205: result <= 12'b010110101001;
   8206: result <= 12'b010110101010;
   8207: result <= 12'b010110101010;
   8208: result <= 12'b010110101010;
   8209: result <= 12'b010110101010;
   8210: result <= 12'b010110101010;
   8211: result <= 12'b010110101010;
   8212: result <= 12'b010110101010;
   8213: result <= 12'b010110101011;
   8214: result <= 12'b010110101011;
   8215: result <= 12'b010110101011;
   8216: result <= 12'b010110101011;
   8217: result <= 12'b010110101011;
   8218: result <= 12'b010110101011;
   8219: result <= 12'b010110101011;
   8220: result <= 12'b010110101100;
   8221: result <= 12'b010110101100;
   8222: result <= 12'b010110101100;
   8223: result <= 12'b010110101100;
   8224: result <= 12'b010110101100;
   8225: result <= 12'b010110101100;
   8226: result <= 12'b010110101100;
   8227: result <= 12'b010110101101;
   8228: result <= 12'b010110101101;
   8229: result <= 12'b010110101101;
   8230: result <= 12'b010110101101;
   8231: result <= 12'b010110101101;
   8232: result <= 12'b010110101101;
   8233: result <= 12'b010110101101;
   8234: result <= 12'b010110101101;
   8235: result <= 12'b010110101110;
   8236: result <= 12'b010110101110;
   8237: result <= 12'b010110101110;
   8238: result <= 12'b010110101110;
   8239: result <= 12'b010110101110;
   8240: result <= 12'b010110101110;
   8241: result <= 12'b010110101110;
   8242: result <= 12'b010110101111;
   8243: result <= 12'b010110101111;
   8244: result <= 12'b010110101111;
   8245: result <= 12'b010110101111;
   8246: result <= 12'b010110101111;
   8247: result <= 12'b010110101111;
   8248: result <= 12'b010110101111;
   8249: result <= 12'b010110110000;
   8250: result <= 12'b010110110000;
   8251: result <= 12'b010110110000;
   8252: result <= 12'b010110110000;
   8253: result <= 12'b010110110000;
   8254: result <= 12'b010110110000;
   8255: result <= 12'b010110110000;
   8256: result <= 12'b010110110001;
   8257: result <= 12'b010110110001;
   8258: result <= 12'b010110110001;
   8259: result <= 12'b010110110001;
   8260: result <= 12'b010110110001;
   8261: result <= 12'b010110110001;
   8262: result <= 12'b010110110001;
   8263: result <= 12'b010110110001;
   8264: result <= 12'b010110110010;
   8265: result <= 12'b010110110010;
   8266: result <= 12'b010110110010;
   8267: result <= 12'b010110110010;
   8268: result <= 12'b010110110010;
   8269: result <= 12'b010110110010;
   8270: result <= 12'b010110110010;
   8271: result <= 12'b010110110011;
   8272: result <= 12'b010110110011;
   8273: result <= 12'b010110110011;
   8274: result <= 12'b010110110011;
   8275: result <= 12'b010110110011;
   8276: result <= 12'b010110110011;
   8277: result <= 12'b010110110011;
   8278: result <= 12'b010110110100;
   8279: result <= 12'b010110110100;
   8280: result <= 12'b010110110100;
   8281: result <= 12'b010110110100;
   8282: result <= 12'b010110110100;
   8283: result <= 12'b010110110100;
   8284: result <= 12'b010110110100;
   8285: result <= 12'b010110110101;
   8286: result <= 12'b010110110101;
   8287: result <= 12'b010110110101;
   8288: result <= 12'b010110110101;
   8289: result <= 12'b010110110101;
   8290: result <= 12'b010110110101;
   8291: result <= 12'b010110110101;
   8292: result <= 12'b010110110101;
   8293: result <= 12'b010110110110;
   8294: result <= 12'b010110110110;
   8295: result <= 12'b010110110110;
   8296: result <= 12'b010110110110;
   8297: result <= 12'b010110110110;
   8298: result <= 12'b010110110110;
   8299: result <= 12'b010110110110;
   8300: result <= 12'b010110110111;
   8301: result <= 12'b010110110111;
   8302: result <= 12'b010110110111;
   8303: result <= 12'b010110110111;
   8304: result <= 12'b010110110111;
   8305: result <= 12'b010110110111;
   8306: result <= 12'b010110110111;
   8307: result <= 12'b010110111000;
   8308: result <= 12'b010110111000;
   8309: result <= 12'b010110111000;
   8310: result <= 12'b010110111000;
   8311: result <= 12'b010110111000;
   8312: result <= 12'b010110111000;
   8313: result <= 12'b010110111000;
   8314: result <= 12'b010110111000;
   8315: result <= 12'b010110111001;
   8316: result <= 12'b010110111001;
   8317: result <= 12'b010110111001;
   8318: result <= 12'b010110111001;
   8319: result <= 12'b010110111001;
   8320: result <= 12'b010110111001;
   8321: result <= 12'b010110111001;
   8322: result <= 12'b010110111010;
   8323: result <= 12'b010110111010;
   8324: result <= 12'b010110111010;
   8325: result <= 12'b010110111010;
   8326: result <= 12'b010110111010;
   8327: result <= 12'b010110111010;
   8328: result <= 12'b010110111010;
   8329: result <= 12'b010110111011;
   8330: result <= 12'b010110111011;
   8331: result <= 12'b010110111011;
   8332: result <= 12'b010110111011;
   8333: result <= 12'b010110111011;
   8334: result <= 12'b010110111011;
   8335: result <= 12'b010110111011;
   8336: result <= 12'b010110111100;
   8337: result <= 12'b010110111100;
   8338: result <= 12'b010110111100;
   8339: result <= 12'b010110111100;
   8340: result <= 12'b010110111100;
   8341: result <= 12'b010110111100;
   8342: result <= 12'b010110111100;
   8343: result <= 12'b010110111100;
   8344: result <= 12'b010110111101;
   8345: result <= 12'b010110111101;
   8346: result <= 12'b010110111101;
   8347: result <= 12'b010110111101;
   8348: result <= 12'b010110111101;
   8349: result <= 12'b010110111101;
   8350: result <= 12'b010110111101;
   8351: result <= 12'b010110111110;
   8352: result <= 12'b010110111110;
   8353: result <= 12'b010110111110;
   8354: result <= 12'b010110111110;
   8355: result <= 12'b010110111110;
   8356: result <= 12'b010110111110;
   8357: result <= 12'b010110111110;
   8358: result <= 12'b010110111111;
   8359: result <= 12'b010110111111;
   8360: result <= 12'b010110111111;
   8361: result <= 12'b010110111111;
   8362: result <= 12'b010110111111;
   8363: result <= 12'b010110111111;
   8364: result <= 12'b010110111111;
   8365: result <= 12'b010110111111;
   8366: result <= 12'b010111000000;
   8367: result <= 12'b010111000000;
   8368: result <= 12'b010111000000;
   8369: result <= 12'b010111000000;
   8370: result <= 12'b010111000000;
   8371: result <= 12'b010111000000;
   8372: result <= 12'b010111000000;
   8373: result <= 12'b010111000001;
   8374: result <= 12'b010111000001;
   8375: result <= 12'b010111000001;
   8376: result <= 12'b010111000001;
   8377: result <= 12'b010111000001;
   8378: result <= 12'b010111000001;
   8379: result <= 12'b010111000001;
   8380: result <= 12'b010111000010;
   8381: result <= 12'b010111000010;
   8382: result <= 12'b010111000010;
   8383: result <= 12'b010111000010;
   8384: result <= 12'b010111000010;
   8385: result <= 12'b010111000010;
   8386: result <= 12'b010111000010;
   8387: result <= 12'b010111000010;
   8388: result <= 12'b010111000011;
   8389: result <= 12'b010111000011;
   8390: result <= 12'b010111000011;
   8391: result <= 12'b010111000011;
   8392: result <= 12'b010111000011;
   8393: result <= 12'b010111000011;
   8394: result <= 12'b010111000011;
   8395: result <= 12'b010111000100;
   8396: result <= 12'b010111000100;
   8397: result <= 12'b010111000100;
   8398: result <= 12'b010111000100;
   8399: result <= 12'b010111000100;
   8400: result <= 12'b010111000100;
   8401: result <= 12'b010111000100;
   8402: result <= 12'b010111000101;
   8403: result <= 12'b010111000101;
   8404: result <= 12'b010111000101;
   8405: result <= 12'b010111000101;
   8406: result <= 12'b010111000101;
   8407: result <= 12'b010111000101;
   8408: result <= 12'b010111000101;
   8409: result <= 12'b010111000101;
   8410: result <= 12'b010111000110;
   8411: result <= 12'b010111000110;
   8412: result <= 12'b010111000110;
   8413: result <= 12'b010111000110;
   8414: result <= 12'b010111000110;
   8415: result <= 12'b010111000110;
   8416: result <= 12'b010111000110;
   8417: result <= 12'b010111000111;
   8418: result <= 12'b010111000111;
   8419: result <= 12'b010111000111;
   8420: result <= 12'b010111000111;
   8421: result <= 12'b010111000111;
   8422: result <= 12'b010111000111;
   8423: result <= 12'b010111000111;
   8424: result <= 12'b010111001000;
   8425: result <= 12'b010111001000;
   8426: result <= 12'b010111001000;
   8427: result <= 12'b010111001000;
   8428: result <= 12'b010111001000;
   8429: result <= 12'b010111001000;
   8430: result <= 12'b010111001000;
   8431: result <= 12'b010111001000;
   8432: result <= 12'b010111001001;
   8433: result <= 12'b010111001001;
   8434: result <= 12'b010111001001;
   8435: result <= 12'b010111001001;
   8436: result <= 12'b010111001001;
   8437: result <= 12'b010111001001;
   8438: result <= 12'b010111001001;
   8439: result <= 12'b010111001010;
   8440: result <= 12'b010111001010;
   8441: result <= 12'b010111001010;
   8442: result <= 12'b010111001010;
   8443: result <= 12'b010111001010;
   8444: result <= 12'b010111001010;
   8445: result <= 12'b010111001010;
   8446: result <= 12'b010111001010;
   8447: result <= 12'b010111001011;
   8448: result <= 12'b010111001011;
   8449: result <= 12'b010111001011;
   8450: result <= 12'b010111001011;
   8451: result <= 12'b010111001011;
   8452: result <= 12'b010111001011;
   8453: result <= 12'b010111001011;
   8454: result <= 12'b010111001100;
   8455: result <= 12'b010111001100;
   8456: result <= 12'b010111001100;
   8457: result <= 12'b010111001100;
   8458: result <= 12'b010111001100;
   8459: result <= 12'b010111001100;
   8460: result <= 12'b010111001100;
   8461: result <= 12'b010111001101;
   8462: result <= 12'b010111001101;
   8463: result <= 12'b010111001101;
   8464: result <= 12'b010111001101;
   8465: result <= 12'b010111001101;
   8466: result <= 12'b010111001101;
   8467: result <= 12'b010111001101;
   8468: result <= 12'b010111001101;
   8469: result <= 12'b010111001110;
   8470: result <= 12'b010111001110;
   8471: result <= 12'b010111001110;
   8472: result <= 12'b010111001110;
   8473: result <= 12'b010111001110;
   8474: result <= 12'b010111001110;
   8475: result <= 12'b010111001110;
   8476: result <= 12'b010111001111;
   8477: result <= 12'b010111001111;
   8478: result <= 12'b010111001111;
   8479: result <= 12'b010111001111;
   8480: result <= 12'b010111001111;
   8481: result <= 12'b010111001111;
   8482: result <= 12'b010111001111;
   8483: result <= 12'b010111001111;
   8484: result <= 12'b010111010000;
   8485: result <= 12'b010111010000;
   8486: result <= 12'b010111010000;
   8487: result <= 12'b010111010000;
   8488: result <= 12'b010111010000;
   8489: result <= 12'b010111010000;
   8490: result <= 12'b010111010000;
   8491: result <= 12'b010111010001;
   8492: result <= 12'b010111010001;
   8493: result <= 12'b010111010001;
   8494: result <= 12'b010111010001;
   8495: result <= 12'b010111010001;
   8496: result <= 12'b010111010001;
   8497: result <= 12'b010111010001;
   8498: result <= 12'b010111010010;
   8499: result <= 12'b010111010010;
   8500: result <= 12'b010111010010;
   8501: result <= 12'b010111010010;
   8502: result <= 12'b010111010010;
   8503: result <= 12'b010111010010;
   8504: result <= 12'b010111010010;
   8505: result <= 12'b010111010010;
   8506: result <= 12'b010111010011;
   8507: result <= 12'b010111010011;
   8508: result <= 12'b010111010011;
   8509: result <= 12'b010111010011;
   8510: result <= 12'b010111010011;
   8511: result <= 12'b010111010011;
   8512: result <= 12'b010111010011;
   8513: result <= 12'b010111010100;
   8514: result <= 12'b010111010100;
   8515: result <= 12'b010111010100;
   8516: result <= 12'b010111010100;
   8517: result <= 12'b010111010100;
   8518: result <= 12'b010111010100;
   8519: result <= 12'b010111010100;
   8520: result <= 12'b010111010100;
   8521: result <= 12'b010111010101;
   8522: result <= 12'b010111010101;
   8523: result <= 12'b010111010101;
   8524: result <= 12'b010111010101;
   8525: result <= 12'b010111010101;
   8526: result <= 12'b010111010101;
   8527: result <= 12'b010111010101;
   8528: result <= 12'b010111010110;
   8529: result <= 12'b010111010110;
   8530: result <= 12'b010111010110;
   8531: result <= 12'b010111010110;
   8532: result <= 12'b010111010110;
   8533: result <= 12'b010111010110;
   8534: result <= 12'b010111010110;
   8535: result <= 12'b010111010110;
   8536: result <= 12'b010111010111;
   8537: result <= 12'b010111010111;
   8538: result <= 12'b010111010111;
   8539: result <= 12'b010111010111;
   8540: result <= 12'b010111010111;
   8541: result <= 12'b010111010111;
   8542: result <= 12'b010111010111;
   8543: result <= 12'b010111011000;
   8544: result <= 12'b010111011000;
   8545: result <= 12'b010111011000;
   8546: result <= 12'b010111011000;
   8547: result <= 12'b010111011000;
   8548: result <= 12'b010111011000;
   8549: result <= 12'b010111011000;
   8550: result <= 12'b010111011000;
   8551: result <= 12'b010111011001;
   8552: result <= 12'b010111011001;
   8553: result <= 12'b010111011001;
   8554: result <= 12'b010111011001;
   8555: result <= 12'b010111011001;
   8556: result <= 12'b010111011001;
   8557: result <= 12'b010111011001;
   8558: result <= 12'b010111011010;
   8559: result <= 12'b010111011010;
   8560: result <= 12'b010111011010;
   8561: result <= 12'b010111011010;
   8562: result <= 12'b010111011010;
   8563: result <= 12'b010111011010;
   8564: result <= 12'b010111011010;
   8565: result <= 12'b010111011011;
   8566: result <= 12'b010111011011;
   8567: result <= 12'b010111011011;
   8568: result <= 12'b010111011011;
   8569: result <= 12'b010111011011;
   8570: result <= 12'b010111011011;
   8571: result <= 12'b010111011011;
   8572: result <= 12'b010111011011;
   8573: result <= 12'b010111011100;
   8574: result <= 12'b010111011100;
   8575: result <= 12'b010111011100;
   8576: result <= 12'b010111011100;
   8577: result <= 12'b010111011100;
   8578: result <= 12'b010111011100;
   8579: result <= 12'b010111011100;
   8580: result <= 12'b010111011101;
   8581: result <= 12'b010111011101;
   8582: result <= 12'b010111011101;
   8583: result <= 12'b010111011101;
   8584: result <= 12'b010111011101;
   8585: result <= 12'b010111011101;
   8586: result <= 12'b010111011101;
   8587: result <= 12'b010111011101;
   8588: result <= 12'b010111011110;
   8589: result <= 12'b010111011110;
   8590: result <= 12'b010111011110;
   8591: result <= 12'b010111011110;
   8592: result <= 12'b010111011110;
   8593: result <= 12'b010111011110;
   8594: result <= 12'b010111011110;
   8595: result <= 12'b010111011111;
   8596: result <= 12'b010111011111;
   8597: result <= 12'b010111011111;
   8598: result <= 12'b010111011111;
   8599: result <= 12'b010111011111;
   8600: result <= 12'b010111011111;
   8601: result <= 12'b010111011111;
   8602: result <= 12'b010111011111;
   8603: result <= 12'b010111100000;
   8604: result <= 12'b010111100000;
   8605: result <= 12'b010111100000;
   8606: result <= 12'b010111100000;
   8607: result <= 12'b010111100000;
   8608: result <= 12'b010111100000;
   8609: result <= 12'b010111100000;
   8610: result <= 12'b010111100001;
   8611: result <= 12'b010111100001;
   8612: result <= 12'b010111100001;
   8613: result <= 12'b010111100001;
   8614: result <= 12'b010111100001;
   8615: result <= 12'b010111100001;
   8616: result <= 12'b010111100001;
   8617: result <= 12'b010111100001;
   8618: result <= 12'b010111100010;
   8619: result <= 12'b010111100010;
   8620: result <= 12'b010111100010;
   8621: result <= 12'b010111100010;
   8622: result <= 12'b010111100010;
   8623: result <= 12'b010111100010;
   8624: result <= 12'b010111100010;
   8625: result <= 12'b010111100011;
   8626: result <= 12'b010111100011;
   8627: result <= 12'b010111100011;
   8628: result <= 12'b010111100011;
   8629: result <= 12'b010111100011;
   8630: result <= 12'b010111100011;
   8631: result <= 12'b010111100011;
   8632: result <= 12'b010111100011;
   8633: result <= 12'b010111100100;
   8634: result <= 12'b010111100100;
   8635: result <= 12'b010111100100;
   8636: result <= 12'b010111100100;
   8637: result <= 12'b010111100100;
   8638: result <= 12'b010111100100;
   8639: result <= 12'b010111100100;
   8640: result <= 12'b010111100101;
   8641: result <= 12'b010111100101;
   8642: result <= 12'b010111100101;
   8643: result <= 12'b010111100101;
   8644: result <= 12'b010111100101;
   8645: result <= 12'b010111100101;
   8646: result <= 12'b010111100101;
   8647: result <= 12'b010111100101;
   8648: result <= 12'b010111100110;
   8649: result <= 12'b010111100110;
   8650: result <= 12'b010111100110;
   8651: result <= 12'b010111100110;
   8652: result <= 12'b010111100110;
   8653: result <= 12'b010111100110;
   8654: result <= 12'b010111100110;
   8655: result <= 12'b010111100110;
   8656: result <= 12'b010111100111;
   8657: result <= 12'b010111100111;
   8658: result <= 12'b010111100111;
   8659: result <= 12'b010111100111;
   8660: result <= 12'b010111100111;
   8661: result <= 12'b010111100111;
   8662: result <= 12'b010111100111;
   8663: result <= 12'b010111101000;
   8664: result <= 12'b010111101000;
   8665: result <= 12'b010111101000;
   8666: result <= 12'b010111101000;
   8667: result <= 12'b010111101000;
   8668: result <= 12'b010111101000;
   8669: result <= 12'b010111101000;
   8670: result <= 12'b010111101000;
   8671: result <= 12'b010111101001;
   8672: result <= 12'b010111101001;
   8673: result <= 12'b010111101001;
   8674: result <= 12'b010111101001;
   8675: result <= 12'b010111101001;
   8676: result <= 12'b010111101001;
   8677: result <= 12'b010111101001;
   8678: result <= 12'b010111101010;
   8679: result <= 12'b010111101010;
   8680: result <= 12'b010111101010;
   8681: result <= 12'b010111101010;
   8682: result <= 12'b010111101010;
   8683: result <= 12'b010111101010;
   8684: result <= 12'b010111101010;
   8685: result <= 12'b010111101010;
   8686: result <= 12'b010111101011;
   8687: result <= 12'b010111101011;
   8688: result <= 12'b010111101011;
   8689: result <= 12'b010111101011;
   8690: result <= 12'b010111101011;
   8691: result <= 12'b010111101011;
   8692: result <= 12'b010111101011;
   8693: result <= 12'b010111101100;
   8694: result <= 12'b010111101100;
   8695: result <= 12'b010111101100;
   8696: result <= 12'b010111101100;
   8697: result <= 12'b010111101100;
   8698: result <= 12'b010111101100;
   8699: result <= 12'b010111101100;
   8700: result <= 12'b010111101100;
   8701: result <= 12'b010111101101;
   8702: result <= 12'b010111101101;
   8703: result <= 12'b010111101101;
   8704: result <= 12'b010111101101;
   8705: result <= 12'b010111101101;
   8706: result <= 12'b010111101101;
   8707: result <= 12'b010111101101;
   8708: result <= 12'b010111101101;
   8709: result <= 12'b010111101110;
   8710: result <= 12'b010111101110;
   8711: result <= 12'b010111101110;
   8712: result <= 12'b010111101110;
   8713: result <= 12'b010111101110;
   8714: result <= 12'b010111101110;
   8715: result <= 12'b010111101110;
   8716: result <= 12'b010111101111;
   8717: result <= 12'b010111101111;
   8718: result <= 12'b010111101111;
   8719: result <= 12'b010111101111;
   8720: result <= 12'b010111101111;
   8721: result <= 12'b010111101111;
   8722: result <= 12'b010111101111;
   8723: result <= 12'b010111101111;
   8724: result <= 12'b010111110000;
   8725: result <= 12'b010111110000;
   8726: result <= 12'b010111110000;
   8727: result <= 12'b010111110000;
   8728: result <= 12'b010111110000;
   8729: result <= 12'b010111110000;
   8730: result <= 12'b010111110000;
   8731: result <= 12'b010111110001;
   8732: result <= 12'b010111110001;
   8733: result <= 12'b010111110001;
   8734: result <= 12'b010111110001;
   8735: result <= 12'b010111110001;
   8736: result <= 12'b010111110001;
   8737: result <= 12'b010111110001;
   8738: result <= 12'b010111110001;
   8739: result <= 12'b010111110010;
   8740: result <= 12'b010111110010;
   8741: result <= 12'b010111110010;
   8742: result <= 12'b010111110010;
   8743: result <= 12'b010111110010;
   8744: result <= 12'b010111110010;
   8745: result <= 12'b010111110010;
   8746: result <= 12'b010111110010;
   8747: result <= 12'b010111110011;
   8748: result <= 12'b010111110011;
   8749: result <= 12'b010111110011;
   8750: result <= 12'b010111110011;
   8751: result <= 12'b010111110011;
   8752: result <= 12'b010111110011;
   8753: result <= 12'b010111110011;
   8754: result <= 12'b010111110100;
   8755: result <= 12'b010111110100;
   8756: result <= 12'b010111110100;
   8757: result <= 12'b010111110100;
   8758: result <= 12'b010111110100;
   8759: result <= 12'b010111110100;
   8760: result <= 12'b010111110100;
   8761: result <= 12'b010111110100;
   8762: result <= 12'b010111110101;
   8763: result <= 12'b010111110101;
   8764: result <= 12'b010111110101;
   8765: result <= 12'b010111110101;
   8766: result <= 12'b010111110101;
   8767: result <= 12'b010111110101;
   8768: result <= 12'b010111110101;
   8769: result <= 12'b010111110110;
   8770: result <= 12'b010111110110;
   8771: result <= 12'b010111110110;
   8772: result <= 12'b010111110110;
   8773: result <= 12'b010111110110;
   8774: result <= 12'b010111110110;
   8775: result <= 12'b010111110110;
   8776: result <= 12'b010111110110;
   8777: result <= 12'b010111110111;
   8778: result <= 12'b010111110111;
   8779: result <= 12'b010111110111;
   8780: result <= 12'b010111110111;
   8781: result <= 12'b010111110111;
   8782: result <= 12'b010111110111;
   8783: result <= 12'b010111110111;
   8784: result <= 12'b010111110111;
   8785: result <= 12'b010111111000;
   8786: result <= 12'b010111111000;
   8787: result <= 12'b010111111000;
   8788: result <= 12'b010111111000;
   8789: result <= 12'b010111111000;
   8790: result <= 12'b010111111000;
   8791: result <= 12'b010111111000;
   8792: result <= 12'b010111111001;
   8793: result <= 12'b010111111001;
   8794: result <= 12'b010111111001;
   8795: result <= 12'b010111111001;
   8796: result <= 12'b010111111001;
   8797: result <= 12'b010111111001;
   8798: result <= 12'b010111111001;
   8799: result <= 12'b010111111001;
   8800: result <= 12'b010111111010;
   8801: result <= 12'b010111111010;
   8802: result <= 12'b010111111010;
   8803: result <= 12'b010111111010;
   8804: result <= 12'b010111111010;
   8805: result <= 12'b010111111010;
   8806: result <= 12'b010111111010;
   8807: result <= 12'b010111111010;
   8808: result <= 12'b010111111011;
   8809: result <= 12'b010111111011;
   8810: result <= 12'b010111111011;
   8811: result <= 12'b010111111011;
   8812: result <= 12'b010111111011;
   8813: result <= 12'b010111111011;
   8814: result <= 12'b010111111011;
   8815: result <= 12'b010111111100;
   8816: result <= 12'b010111111100;
   8817: result <= 12'b010111111100;
   8818: result <= 12'b010111111100;
   8819: result <= 12'b010111111100;
   8820: result <= 12'b010111111100;
   8821: result <= 12'b010111111100;
   8822: result <= 12'b010111111100;
   8823: result <= 12'b010111111101;
   8824: result <= 12'b010111111101;
   8825: result <= 12'b010111111101;
   8826: result <= 12'b010111111101;
   8827: result <= 12'b010111111101;
   8828: result <= 12'b010111111101;
   8829: result <= 12'b010111111101;
   8830: result <= 12'b010111111101;
   8831: result <= 12'b010111111110;
   8832: result <= 12'b010111111110;
   8833: result <= 12'b010111111110;
   8834: result <= 12'b010111111110;
   8835: result <= 12'b010111111110;
   8836: result <= 12'b010111111110;
   8837: result <= 12'b010111111110;
   8838: result <= 12'b010111111111;
   8839: result <= 12'b010111111111;
   8840: result <= 12'b010111111111;
   8841: result <= 12'b010111111111;
   8842: result <= 12'b010111111111;
   8843: result <= 12'b010111111111;
   8844: result <= 12'b010111111111;
   8845: result <= 12'b010111111111;
   8846: result <= 12'b011000000000;
   8847: result <= 12'b011000000000;
   8848: result <= 12'b011000000000;
   8849: result <= 12'b011000000000;
   8850: result <= 12'b011000000000;
   8851: result <= 12'b011000000000;
   8852: result <= 12'b011000000000;
   8853: result <= 12'b011000000000;
   8854: result <= 12'b011000000001;
   8855: result <= 12'b011000000001;
   8856: result <= 12'b011000000001;
   8857: result <= 12'b011000000001;
   8858: result <= 12'b011000000001;
   8859: result <= 12'b011000000001;
   8860: result <= 12'b011000000001;
   8861: result <= 12'b011000000001;
   8862: result <= 12'b011000000010;
   8863: result <= 12'b011000000010;
   8864: result <= 12'b011000000010;
   8865: result <= 12'b011000000010;
   8866: result <= 12'b011000000010;
   8867: result <= 12'b011000000010;
   8868: result <= 12'b011000000010;
   8869: result <= 12'b011000000011;
   8870: result <= 12'b011000000011;
   8871: result <= 12'b011000000011;
   8872: result <= 12'b011000000011;
   8873: result <= 12'b011000000011;
   8874: result <= 12'b011000000011;
   8875: result <= 12'b011000000011;
   8876: result <= 12'b011000000011;
   8877: result <= 12'b011000000100;
   8878: result <= 12'b011000000100;
   8879: result <= 12'b011000000100;
   8880: result <= 12'b011000000100;
   8881: result <= 12'b011000000100;
   8882: result <= 12'b011000000100;
   8883: result <= 12'b011000000100;
   8884: result <= 12'b011000000100;
   8885: result <= 12'b011000000101;
   8886: result <= 12'b011000000101;
   8887: result <= 12'b011000000101;
   8888: result <= 12'b011000000101;
   8889: result <= 12'b011000000101;
   8890: result <= 12'b011000000101;
   8891: result <= 12'b011000000101;
   8892: result <= 12'b011000000110;
   8893: result <= 12'b011000000110;
   8894: result <= 12'b011000000110;
   8895: result <= 12'b011000000110;
   8896: result <= 12'b011000000110;
   8897: result <= 12'b011000000110;
   8898: result <= 12'b011000000110;
   8899: result <= 12'b011000000110;
   8900: result <= 12'b011000000111;
   8901: result <= 12'b011000000111;
   8902: result <= 12'b011000000111;
   8903: result <= 12'b011000000111;
   8904: result <= 12'b011000000111;
   8905: result <= 12'b011000000111;
   8906: result <= 12'b011000000111;
   8907: result <= 12'b011000000111;
   8908: result <= 12'b011000001000;
   8909: result <= 12'b011000001000;
   8910: result <= 12'b011000001000;
   8911: result <= 12'b011000001000;
   8912: result <= 12'b011000001000;
   8913: result <= 12'b011000001000;
   8914: result <= 12'b011000001000;
   8915: result <= 12'b011000001000;
   8916: result <= 12'b011000001001;
   8917: result <= 12'b011000001001;
   8918: result <= 12'b011000001001;
   8919: result <= 12'b011000001001;
   8920: result <= 12'b011000001001;
   8921: result <= 12'b011000001001;
   8922: result <= 12'b011000001001;
   8923: result <= 12'b011000001010;
   8924: result <= 12'b011000001010;
   8925: result <= 12'b011000001010;
   8926: result <= 12'b011000001010;
   8927: result <= 12'b011000001010;
   8928: result <= 12'b011000001010;
   8929: result <= 12'b011000001010;
   8930: result <= 12'b011000001010;
   8931: result <= 12'b011000001011;
   8932: result <= 12'b011000001011;
   8933: result <= 12'b011000001011;
   8934: result <= 12'b011000001011;
   8935: result <= 12'b011000001011;
   8936: result <= 12'b011000001011;
   8937: result <= 12'b011000001011;
   8938: result <= 12'b011000001011;
   8939: result <= 12'b011000001100;
   8940: result <= 12'b011000001100;
   8941: result <= 12'b011000001100;
   8942: result <= 12'b011000001100;
   8943: result <= 12'b011000001100;
   8944: result <= 12'b011000001100;
   8945: result <= 12'b011000001100;
   8946: result <= 12'b011000001100;
   8947: result <= 12'b011000001101;
   8948: result <= 12'b011000001101;
   8949: result <= 12'b011000001101;
   8950: result <= 12'b011000001101;
   8951: result <= 12'b011000001101;
   8952: result <= 12'b011000001101;
   8953: result <= 12'b011000001101;
   8954: result <= 12'b011000001101;
   8955: result <= 12'b011000001110;
   8956: result <= 12'b011000001110;
   8957: result <= 12'b011000001110;
   8958: result <= 12'b011000001110;
   8959: result <= 12'b011000001110;
   8960: result <= 12'b011000001110;
   8961: result <= 12'b011000001110;
   8962: result <= 12'b011000001111;
   8963: result <= 12'b011000001111;
   8964: result <= 12'b011000001111;
   8965: result <= 12'b011000001111;
   8966: result <= 12'b011000001111;
   8967: result <= 12'b011000001111;
   8968: result <= 12'b011000001111;
   8969: result <= 12'b011000001111;
   8970: result <= 12'b011000010000;
   8971: result <= 12'b011000010000;
   8972: result <= 12'b011000010000;
   8973: result <= 12'b011000010000;
   8974: result <= 12'b011000010000;
   8975: result <= 12'b011000010000;
   8976: result <= 12'b011000010000;
   8977: result <= 12'b011000010000;
   8978: result <= 12'b011000010001;
   8979: result <= 12'b011000010001;
   8980: result <= 12'b011000010001;
   8981: result <= 12'b011000010001;
   8982: result <= 12'b011000010001;
   8983: result <= 12'b011000010001;
   8984: result <= 12'b011000010001;
   8985: result <= 12'b011000010001;
   8986: result <= 12'b011000010010;
   8987: result <= 12'b011000010010;
   8988: result <= 12'b011000010010;
   8989: result <= 12'b011000010010;
   8990: result <= 12'b011000010010;
   8991: result <= 12'b011000010010;
   8992: result <= 12'b011000010010;
   8993: result <= 12'b011000010010;
   8994: result <= 12'b011000010011;
   8995: result <= 12'b011000010011;
   8996: result <= 12'b011000010011;
   8997: result <= 12'b011000010011;
   8998: result <= 12'b011000010011;
   8999: result <= 12'b011000010011;
   9000: result <= 12'b011000010011;
   9001: result <= 12'b011000010100;
   9002: result <= 12'b011000010100;
   9003: result <= 12'b011000010100;
   9004: result <= 12'b011000010100;
   9005: result <= 12'b011000010100;
   9006: result <= 12'b011000010100;
   9007: result <= 12'b011000010100;
   9008: result <= 12'b011000010100;
   9009: result <= 12'b011000010101;
   9010: result <= 12'b011000010101;
   9011: result <= 12'b011000010101;
   9012: result <= 12'b011000010101;
   9013: result <= 12'b011000010101;
   9014: result <= 12'b011000010101;
   9015: result <= 12'b011000010101;
   9016: result <= 12'b011000010101;
   9017: result <= 12'b011000010110;
   9018: result <= 12'b011000010110;
   9019: result <= 12'b011000010110;
   9020: result <= 12'b011000010110;
   9021: result <= 12'b011000010110;
   9022: result <= 12'b011000010110;
   9023: result <= 12'b011000010110;
   9024: result <= 12'b011000010110;
   9025: result <= 12'b011000010111;
   9026: result <= 12'b011000010111;
   9027: result <= 12'b011000010111;
   9028: result <= 12'b011000010111;
   9029: result <= 12'b011000010111;
   9030: result <= 12'b011000010111;
   9031: result <= 12'b011000010111;
   9032: result <= 12'b011000010111;
   9033: result <= 12'b011000011000;
   9034: result <= 12'b011000011000;
   9035: result <= 12'b011000011000;
   9036: result <= 12'b011000011000;
   9037: result <= 12'b011000011000;
   9038: result <= 12'b011000011000;
   9039: result <= 12'b011000011000;
   9040: result <= 12'b011000011000;
   9041: result <= 12'b011000011001;
   9042: result <= 12'b011000011001;
   9043: result <= 12'b011000011001;
   9044: result <= 12'b011000011001;
   9045: result <= 12'b011000011001;
   9046: result <= 12'b011000011001;
   9047: result <= 12'b011000011001;
   9048: result <= 12'b011000011001;
   9049: result <= 12'b011000011010;
   9050: result <= 12'b011000011010;
   9051: result <= 12'b011000011010;
   9052: result <= 12'b011000011010;
   9053: result <= 12'b011000011010;
   9054: result <= 12'b011000011010;
   9055: result <= 12'b011000011010;
   9056: result <= 12'b011000011011;
   9057: result <= 12'b011000011011;
   9058: result <= 12'b011000011011;
   9059: result <= 12'b011000011011;
   9060: result <= 12'b011000011011;
   9061: result <= 12'b011000011011;
   9062: result <= 12'b011000011011;
   9063: result <= 12'b011000011011;
   9064: result <= 12'b011000011100;
   9065: result <= 12'b011000011100;
   9066: result <= 12'b011000011100;
   9067: result <= 12'b011000011100;
   9068: result <= 12'b011000011100;
   9069: result <= 12'b011000011100;
   9070: result <= 12'b011000011100;
   9071: result <= 12'b011000011100;
   9072: result <= 12'b011000011101;
   9073: result <= 12'b011000011101;
   9074: result <= 12'b011000011101;
   9075: result <= 12'b011000011101;
   9076: result <= 12'b011000011101;
   9077: result <= 12'b011000011101;
   9078: result <= 12'b011000011101;
   9079: result <= 12'b011000011101;
   9080: result <= 12'b011000011110;
   9081: result <= 12'b011000011110;
   9082: result <= 12'b011000011110;
   9083: result <= 12'b011000011110;
   9084: result <= 12'b011000011110;
   9085: result <= 12'b011000011110;
   9086: result <= 12'b011000011110;
   9087: result <= 12'b011000011110;
   9088: result <= 12'b011000011111;
   9089: result <= 12'b011000011111;
   9090: result <= 12'b011000011111;
   9091: result <= 12'b011000011111;
   9092: result <= 12'b011000011111;
   9093: result <= 12'b011000011111;
   9094: result <= 12'b011000011111;
   9095: result <= 12'b011000011111;
   9096: result <= 12'b011000100000;
   9097: result <= 12'b011000100000;
   9098: result <= 12'b011000100000;
   9099: result <= 12'b011000100000;
   9100: result <= 12'b011000100000;
   9101: result <= 12'b011000100000;
   9102: result <= 12'b011000100000;
   9103: result <= 12'b011000100000;
   9104: result <= 12'b011000100001;
   9105: result <= 12'b011000100001;
   9106: result <= 12'b011000100001;
   9107: result <= 12'b011000100001;
   9108: result <= 12'b011000100001;
   9109: result <= 12'b011000100001;
   9110: result <= 12'b011000100001;
   9111: result <= 12'b011000100001;
   9112: result <= 12'b011000100010;
   9113: result <= 12'b011000100010;
   9114: result <= 12'b011000100010;
   9115: result <= 12'b011000100010;
   9116: result <= 12'b011000100010;
   9117: result <= 12'b011000100010;
   9118: result <= 12'b011000100010;
   9119: result <= 12'b011000100010;
   9120: result <= 12'b011000100011;
   9121: result <= 12'b011000100011;
   9122: result <= 12'b011000100011;
   9123: result <= 12'b011000100011;
   9124: result <= 12'b011000100011;
   9125: result <= 12'b011000100011;
   9126: result <= 12'b011000100011;
   9127: result <= 12'b011000100011;
   9128: result <= 12'b011000100100;
   9129: result <= 12'b011000100100;
   9130: result <= 12'b011000100100;
   9131: result <= 12'b011000100100;
   9132: result <= 12'b011000100100;
   9133: result <= 12'b011000100100;
   9134: result <= 12'b011000100100;
   9135: result <= 12'b011000100100;
   9136: result <= 12'b011000100101;
   9137: result <= 12'b011000100101;
   9138: result <= 12'b011000100101;
   9139: result <= 12'b011000100101;
   9140: result <= 12'b011000100101;
   9141: result <= 12'b011000100101;
   9142: result <= 12'b011000100101;
   9143: result <= 12'b011000100101;
   9144: result <= 12'b011000100110;
   9145: result <= 12'b011000100110;
   9146: result <= 12'b011000100110;
   9147: result <= 12'b011000100110;
   9148: result <= 12'b011000100110;
   9149: result <= 12'b011000100110;
   9150: result <= 12'b011000100110;
   9151: result <= 12'b011000100110;
   9152: result <= 12'b011000100111;
   9153: result <= 12'b011000100111;
   9154: result <= 12'b011000100111;
   9155: result <= 12'b011000100111;
   9156: result <= 12'b011000100111;
   9157: result <= 12'b011000100111;
   9158: result <= 12'b011000100111;
   9159: result <= 12'b011000101000;
   9160: result <= 12'b011000101000;
   9161: result <= 12'b011000101000;
   9162: result <= 12'b011000101000;
   9163: result <= 12'b011000101000;
   9164: result <= 12'b011000101000;
   9165: result <= 12'b011000101000;
   9166: result <= 12'b011000101000;
   9167: result <= 12'b011000101001;
   9168: result <= 12'b011000101001;
   9169: result <= 12'b011000101001;
   9170: result <= 12'b011000101001;
   9171: result <= 12'b011000101001;
   9172: result <= 12'b011000101001;
   9173: result <= 12'b011000101001;
   9174: result <= 12'b011000101001;
   9175: result <= 12'b011000101010;
   9176: result <= 12'b011000101010;
   9177: result <= 12'b011000101010;
   9178: result <= 12'b011000101010;
   9179: result <= 12'b011000101010;
   9180: result <= 12'b011000101010;
   9181: result <= 12'b011000101010;
   9182: result <= 12'b011000101010;
   9183: result <= 12'b011000101011;
   9184: result <= 12'b011000101011;
   9185: result <= 12'b011000101011;
   9186: result <= 12'b011000101011;
   9187: result <= 12'b011000101011;
   9188: result <= 12'b011000101011;
   9189: result <= 12'b011000101011;
   9190: result <= 12'b011000101011;
   9191: result <= 12'b011000101100;
   9192: result <= 12'b011000101100;
   9193: result <= 12'b011000101100;
   9194: result <= 12'b011000101100;
   9195: result <= 12'b011000101100;
   9196: result <= 12'b011000101100;
   9197: result <= 12'b011000101100;
   9198: result <= 12'b011000101100;
   9199: result <= 12'b011000101101;
   9200: result <= 12'b011000101101;
   9201: result <= 12'b011000101101;
   9202: result <= 12'b011000101101;
   9203: result <= 12'b011000101101;
   9204: result <= 12'b011000101101;
   9205: result <= 12'b011000101101;
   9206: result <= 12'b011000101101;
   9207: result <= 12'b011000101110;
   9208: result <= 12'b011000101110;
   9209: result <= 12'b011000101110;
   9210: result <= 12'b011000101110;
   9211: result <= 12'b011000101110;
   9212: result <= 12'b011000101110;
   9213: result <= 12'b011000101110;
   9214: result <= 12'b011000101110;
   9215: result <= 12'b011000101111;
   9216: result <= 12'b011000101111;
   9217: result <= 12'b011000101111;
   9218: result <= 12'b011000101111;
   9219: result <= 12'b011000101111;
   9220: result <= 12'b011000101111;
   9221: result <= 12'b011000101111;
   9222: result <= 12'b011000101111;
   9223: result <= 12'b011000101111;
   9224: result <= 12'b011000110000;
   9225: result <= 12'b011000110000;
   9226: result <= 12'b011000110000;
   9227: result <= 12'b011000110000;
   9228: result <= 12'b011000110000;
   9229: result <= 12'b011000110000;
   9230: result <= 12'b011000110000;
   9231: result <= 12'b011000110000;
   9232: result <= 12'b011000110001;
   9233: result <= 12'b011000110001;
   9234: result <= 12'b011000110001;
   9235: result <= 12'b011000110001;
   9236: result <= 12'b011000110001;
   9237: result <= 12'b011000110001;
   9238: result <= 12'b011000110001;
   9239: result <= 12'b011000110001;
   9240: result <= 12'b011000110010;
   9241: result <= 12'b011000110010;
   9242: result <= 12'b011000110010;
   9243: result <= 12'b011000110010;
   9244: result <= 12'b011000110010;
   9245: result <= 12'b011000110010;
   9246: result <= 12'b011000110010;
   9247: result <= 12'b011000110010;
   9248: result <= 12'b011000110011;
   9249: result <= 12'b011000110011;
   9250: result <= 12'b011000110011;
   9251: result <= 12'b011000110011;
   9252: result <= 12'b011000110011;
   9253: result <= 12'b011000110011;
   9254: result <= 12'b011000110011;
   9255: result <= 12'b011000110011;
   9256: result <= 12'b011000110100;
   9257: result <= 12'b011000110100;
   9258: result <= 12'b011000110100;
   9259: result <= 12'b011000110100;
   9260: result <= 12'b011000110100;
   9261: result <= 12'b011000110100;
   9262: result <= 12'b011000110100;
   9263: result <= 12'b011000110100;
   9264: result <= 12'b011000110101;
   9265: result <= 12'b011000110101;
   9266: result <= 12'b011000110101;
   9267: result <= 12'b011000110101;
   9268: result <= 12'b011000110101;
   9269: result <= 12'b011000110101;
   9270: result <= 12'b011000110101;
   9271: result <= 12'b011000110101;
   9272: result <= 12'b011000110110;
   9273: result <= 12'b011000110110;
   9274: result <= 12'b011000110110;
   9275: result <= 12'b011000110110;
   9276: result <= 12'b011000110110;
   9277: result <= 12'b011000110110;
   9278: result <= 12'b011000110110;
   9279: result <= 12'b011000110110;
   9280: result <= 12'b011000110111;
   9281: result <= 12'b011000110111;
   9282: result <= 12'b011000110111;
   9283: result <= 12'b011000110111;
   9284: result <= 12'b011000110111;
   9285: result <= 12'b011000110111;
   9286: result <= 12'b011000110111;
   9287: result <= 12'b011000110111;
   9288: result <= 12'b011000111000;
   9289: result <= 12'b011000111000;
   9290: result <= 12'b011000111000;
   9291: result <= 12'b011000111000;
   9292: result <= 12'b011000111000;
   9293: result <= 12'b011000111000;
   9294: result <= 12'b011000111000;
   9295: result <= 12'b011000111000;
   9296: result <= 12'b011000111001;
   9297: result <= 12'b011000111001;
   9298: result <= 12'b011000111001;
   9299: result <= 12'b011000111001;
   9300: result <= 12'b011000111001;
   9301: result <= 12'b011000111001;
   9302: result <= 12'b011000111001;
   9303: result <= 12'b011000111001;
   9304: result <= 12'b011000111010;
   9305: result <= 12'b011000111010;
   9306: result <= 12'b011000111010;
   9307: result <= 12'b011000111010;
   9308: result <= 12'b011000111010;
   9309: result <= 12'b011000111010;
   9310: result <= 12'b011000111010;
   9311: result <= 12'b011000111010;
   9312: result <= 12'b011000111011;
   9313: result <= 12'b011000111011;
   9314: result <= 12'b011000111011;
   9315: result <= 12'b011000111011;
   9316: result <= 12'b011000111011;
   9317: result <= 12'b011000111011;
   9318: result <= 12'b011000111011;
   9319: result <= 12'b011000111011;
   9320: result <= 12'b011000111100;
   9321: result <= 12'b011000111100;
   9322: result <= 12'b011000111100;
   9323: result <= 12'b011000111100;
   9324: result <= 12'b011000111100;
   9325: result <= 12'b011000111100;
   9326: result <= 12'b011000111100;
   9327: result <= 12'b011000111100;
   9328: result <= 12'b011000111100;
   9329: result <= 12'b011000111101;
   9330: result <= 12'b011000111101;
   9331: result <= 12'b011000111101;
   9332: result <= 12'b011000111101;
   9333: result <= 12'b011000111101;
   9334: result <= 12'b011000111101;
   9335: result <= 12'b011000111101;
   9336: result <= 12'b011000111101;
   9337: result <= 12'b011000111110;
   9338: result <= 12'b011000111110;
   9339: result <= 12'b011000111110;
   9340: result <= 12'b011000111110;
   9341: result <= 12'b011000111110;
   9342: result <= 12'b011000111110;
   9343: result <= 12'b011000111110;
   9344: result <= 12'b011000111110;
   9345: result <= 12'b011000111111;
   9346: result <= 12'b011000111111;
   9347: result <= 12'b011000111111;
   9348: result <= 12'b011000111111;
   9349: result <= 12'b011000111111;
   9350: result <= 12'b011000111111;
   9351: result <= 12'b011000111111;
   9352: result <= 12'b011000111111;
   9353: result <= 12'b011001000000;
   9354: result <= 12'b011001000000;
   9355: result <= 12'b011001000000;
   9356: result <= 12'b011001000000;
   9357: result <= 12'b011001000000;
   9358: result <= 12'b011001000000;
   9359: result <= 12'b011001000000;
   9360: result <= 12'b011001000000;
   9361: result <= 12'b011001000001;
   9362: result <= 12'b011001000001;
   9363: result <= 12'b011001000001;
   9364: result <= 12'b011001000001;
   9365: result <= 12'b011001000001;
   9366: result <= 12'b011001000001;
   9367: result <= 12'b011001000001;
   9368: result <= 12'b011001000001;
   9369: result <= 12'b011001000010;
   9370: result <= 12'b011001000010;
   9371: result <= 12'b011001000010;
   9372: result <= 12'b011001000010;
   9373: result <= 12'b011001000010;
   9374: result <= 12'b011001000010;
   9375: result <= 12'b011001000010;
   9376: result <= 12'b011001000010;
   9377: result <= 12'b011001000010;
   9378: result <= 12'b011001000011;
   9379: result <= 12'b011001000011;
   9380: result <= 12'b011001000011;
   9381: result <= 12'b011001000011;
   9382: result <= 12'b011001000011;
   9383: result <= 12'b011001000011;
   9384: result <= 12'b011001000011;
   9385: result <= 12'b011001000011;
   9386: result <= 12'b011001000100;
   9387: result <= 12'b011001000100;
   9388: result <= 12'b011001000100;
   9389: result <= 12'b011001000100;
   9390: result <= 12'b011001000100;
   9391: result <= 12'b011001000100;
   9392: result <= 12'b011001000100;
   9393: result <= 12'b011001000100;
   9394: result <= 12'b011001000101;
   9395: result <= 12'b011001000101;
   9396: result <= 12'b011001000101;
   9397: result <= 12'b011001000101;
   9398: result <= 12'b011001000101;
   9399: result <= 12'b011001000101;
   9400: result <= 12'b011001000101;
   9401: result <= 12'b011001000101;
   9402: result <= 12'b011001000110;
   9403: result <= 12'b011001000110;
   9404: result <= 12'b011001000110;
   9405: result <= 12'b011001000110;
   9406: result <= 12'b011001000110;
   9407: result <= 12'b011001000110;
   9408: result <= 12'b011001000110;
   9409: result <= 12'b011001000110;
   9410: result <= 12'b011001000111;
   9411: result <= 12'b011001000111;
   9412: result <= 12'b011001000111;
   9413: result <= 12'b011001000111;
   9414: result <= 12'b011001000111;
   9415: result <= 12'b011001000111;
   9416: result <= 12'b011001000111;
   9417: result <= 12'b011001000111;
   9418: result <= 12'b011001000111;
   9419: result <= 12'b011001001000;
   9420: result <= 12'b011001001000;
   9421: result <= 12'b011001001000;
   9422: result <= 12'b011001001000;
   9423: result <= 12'b011001001000;
   9424: result <= 12'b011001001000;
   9425: result <= 12'b011001001000;
   9426: result <= 12'b011001001000;
   9427: result <= 12'b011001001001;
   9428: result <= 12'b011001001001;
   9429: result <= 12'b011001001001;
   9430: result <= 12'b011001001001;
   9431: result <= 12'b011001001001;
   9432: result <= 12'b011001001001;
   9433: result <= 12'b011001001001;
   9434: result <= 12'b011001001001;
   9435: result <= 12'b011001001010;
   9436: result <= 12'b011001001010;
   9437: result <= 12'b011001001010;
   9438: result <= 12'b011001001010;
   9439: result <= 12'b011001001010;
   9440: result <= 12'b011001001010;
   9441: result <= 12'b011001001010;
   9442: result <= 12'b011001001010;
   9443: result <= 12'b011001001011;
   9444: result <= 12'b011001001011;
   9445: result <= 12'b011001001011;
   9446: result <= 12'b011001001011;
   9447: result <= 12'b011001001011;
   9448: result <= 12'b011001001011;
   9449: result <= 12'b011001001011;
   9450: result <= 12'b011001001011;
   9451: result <= 12'b011001001011;
   9452: result <= 12'b011001001100;
   9453: result <= 12'b011001001100;
   9454: result <= 12'b011001001100;
   9455: result <= 12'b011001001100;
   9456: result <= 12'b011001001100;
   9457: result <= 12'b011001001100;
   9458: result <= 12'b011001001100;
   9459: result <= 12'b011001001100;
   9460: result <= 12'b011001001101;
   9461: result <= 12'b011001001101;
   9462: result <= 12'b011001001101;
   9463: result <= 12'b011001001101;
   9464: result <= 12'b011001001101;
   9465: result <= 12'b011001001101;
   9466: result <= 12'b011001001101;
   9467: result <= 12'b011001001101;
   9468: result <= 12'b011001001110;
   9469: result <= 12'b011001001110;
   9470: result <= 12'b011001001110;
   9471: result <= 12'b011001001110;
   9472: result <= 12'b011001001110;
   9473: result <= 12'b011001001110;
   9474: result <= 12'b011001001110;
   9475: result <= 12'b011001001110;
   9476: result <= 12'b011001001111;
   9477: result <= 12'b011001001111;
   9478: result <= 12'b011001001111;
   9479: result <= 12'b011001001111;
   9480: result <= 12'b011001001111;
   9481: result <= 12'b011001001111;
   9482: result <= 12'b011001001111;
   9483: result <= 12'b011001001111;
   9484: result <= 12'b011001001111;
   9485: result <= 12'b011001010000;
   9486: result <= 12'b011001010000;
   9487: result <= 12'b011001010000;
   9488: result <= 12'b011001010000;
   9489: result <= 12'b011001010000;
   9490: result <= 12'b011001010000;
   9491: result <= 12'b011001010000;
   9492: result <= 12'b011001010000;
   9493: result <= 12'b011001010001;
   9494: result <= 12'b011001010001;
   9495: result <= 12'b011001010001;
   9496: result <= 12'b011001010001;
   9497: result <= 12'b011001010001;
   9498: result <= 12'b011001010001;
   9499: result <= 12'b011001010001;
   9500: result <= 12'b011001010001;
   9501: result <= 12'b011001010010;
   9502: result <= 12'b011001010010;
   9503: result <= 12'b011001010010;
   9504: result <= 12'b011001010010;
   9505: result <= 12'b011001010010;
   9506: result <= 12'b011001010010;
   9507: result <= 12'b011001010010;
   9508: result <= 12'b011001010010;
   9509: result <= 12'b011001010010;
   9510: result <= 12'b011001010011;
   9511: result <= 12'b011001010011;
   9512: result <= 12'b011001010011;
   9513: result <= 12'b011001010011;
   9514: result <= 12'b011001010011;
   9515: result <= 12'b011001010011;
   9516: result <= 12'b011001010011;
   9517: result <= 12'b011001010011;
   9518: result <= 12'b011001010100;
   9519: result <= 12'b011001010100;
   9520: result <= 12'b011001010100;
   9521: result <= 12'b011001010100;
   9522: result <= 12'b011001010100;
   9523: result <= 12'b011001010100;
   9524: result <= 12'b011001010100;
   9525: result <= 12'b011001010100;
   9526: result <= 12'b011001010101;
   9527: result <= 12'b011001010101;
   9528: result <= 12'b011001010101;
   9529: result <= 12'b011001010101;
   9530: result <= 12'b011001010101;
   9531: result <= 12'b011001010101;
   9532: result <= 12'b011001010101;
   9533: result <= 12'b011001010101;
   9534: result <= 12'b011001010101;
   9535: result <= 12'b011001010110;
   9536: result <= 12'b011001010110;
   9537: result <= 12'b011001010110;
   9538: result <= 12'b011001010110;
   9539: result <= 12'b011001010110;
   9540: result <= 12'b011001010110;
   9541: result <= 12'b011001010110;
   9542: result <= 12'b011001010110;
   9543: result <= 12'b011001010111;
   9544: result <= 12'b011001010111;
   9545: result <= 12'b011001010111;
   9546: result <= 12'b011001010111;
   9547: result <= 12'b011001010111;
   9548: result <= 12'b011001010111;
   9549: result <= 12'b011001010111;
   9550: result <= 12'b011001010111;
   9551: result <= 12'b011001011000;
   9552: result <= 12'b011001011000;
   9553: result <= 12'b011001011000;
   9554: result <= 12'b011001011000;
   9555: result <= 12'b011001011000;
   9556: result <= 12'b011001011000;
   9557: result <= 12'b011001011000;
   9558: result <= 12'b011001011000;
   9559: result <= 12'b011001011000;
   9560: result <= 12'b011001011001;
   9561: result <= 12'b011001011001;
   9562: result <= 12'b011001011001;
   9563: result <= 12'b011001011001;
   9564: result <= 12'b011001011001;
   9565: result <= 12'b011001011001;
   9566: result <= 12'b011001011001;
   9567: result <= 12'b011001011001;
   9568: result <= 12'b011001011010;
   9569: result <= 12'b011001011010;
   9570: result <= 12'b011001011010;
   9571: result <= 12'b011001011010;
   9572: result <= 12'b011001011010;
   9573: result <= 12'b011001011010;
   9574: result <= 12'b011001011010;
   9575: result <= 12'b011001011010;
   9576: result <= 12'b011001011011;
   9577: result <= 12'b011001011011;
   9578: result <= 12'b011001011011;
   9579: result <= 12'b011001011011;
   9580: result <= 12'b011001011011;
   9581: result <= 12'b011001011011;
   9582: result <= 12'b011001011011;
   9583: result <= 12'b011001011011;
   9584: result <= 12'b011001011011;
   9585: result <= 12'b011001011100;
   9586: result <= 12'b011001011100;
   9587: result <= 12'b011001011100;
   9588: result <= 12'b011001011100;
   9589: result <= 12'b011001011100;
   9590: result <= 12'b011001011100;
   9591: result <= 12'b011001011100;
   9592: result <= 12'b011001011100;
   9593: result <= 12'b011001011101;
   9594: result <= 12'b011001011101;
   9595: result <= 12'b011001011101;
   9596: result <= 12'b011001011101;
   9597: result <= 12'b011001011101;
   9598: result <= 12'b011001011101;
   9599: result <= 12'b011001011101;
   9600: result <= 12'b011001011101;
   9601: result <= 12'b011001011101;
   9602: result <= 12'b011001011110;
   9603: result <= 12'b011001011110;
   9604: result <= 12'b011001011110;
   9605: result <= 12'b011001011110;
   9606: result <= 12'b011001011110;
   9607: result <= 12'b011001011110;
   9608: result <= 12'b011001011110;
   9609: result <= 12'b011001011110;
   9610: result <= 12'b011001011111;
   9611: result <= 12'b011001011111;
   9612: result <= 12'b011001011111;
   9613: result <= 12'b011001011111;
   9614: result <= 12'b011001011111;
   9615: result <= 12'b011001011111;
   9616: result <= 12'b011001011111;
   9617: result <= 12'b011001011111;
   9618: result <= 12'b011001100000;
   9619: result <= 12'b011001100000;
   9620: result <= 12'b011001100000;
   9621: result <= 12'b011001100000;
   9622: result <= 12'b011001100000;
   9623: result <= 12'b011001100000;
   9624: result <= 12'b011001100000;
   9625: result <= 12'b011001100000;
   9626: result <= 12'b011001100000;
   9627: result <= 12'b011001100001;
   9628: result <= 12'b011001100001;
   9629: result <= 12'b011001100001;
   9630: result <= 12'b011001100001;
   9631: result <= 12'b011001100001;
   9632: result <= 12'b011001100001;
   9633: result <= 12'b011001100001;
   9634: result <= 12'b011001100001;
   9635: result <= 12'b011001100010;
   9636: result <= 12'b011001100010;
   9637: result <= 12'b011001100010;
   9638: result <= 12'b011001100010;
   9639: result <= 12'b011001100010;
   9640: result <= 12'b011001100010;
   9641: result <= 12'b011001100010;
   9642: result <= 12'b011001100010;
   9643: result <= 12'b011001100010;
   9644: result <= 12'b011001100011;
   9645: result <= 12'b011001100011;
   9646: result <= 12'b011001100011;
   9647: result <= 12'b011001100011;
   9648: result <= 12'b011001100011;
   9649: result <= 12'b011001100011;
   9650: result <= 12'b011001100011;
   9651: result <= 12'b011001100011;
   9652: result <= 12'b011001100100;
   9653: result <= 12'b011001100100;
   9654: result <= 12'b011001100100;
   9655: result <= 12'b011001100100;
   9656: result <= 12'b011001100100;
   9657: result <= 12'b011001100100;
   9658: result <= 12'b011001100100;
   9659: result <= 12'b011001100100;
   9660: result <= 12'b011001100100;
   9661: result <= 12'b011001100101;
   9662: result <= 12'b011001100101;
   9663: result <= 12'b011001100101;
   9664: result <= 12'b011001100101;
   9665: result <= 12'b011001100101;
   9666: result <= 12'b011001100101;
   9667: result <= 12'b011001100101;
   9668: result <= 12'b011001100101;
   9669: result <= 12'b011001100110;
   9670: result <= 12'b011001100110;
   9671: result <= 12'b011001100110;
   9672: result <= 12'b011001100110;
   9673: result <= 12'b011001100110;
   9674: result <= 12'b011001100110;
   9675: result <= 12'b011001100110;
   9676: result <= 12'b011001100110;
   9677: result <= 12'b011001100110;
   9678: result <= 12'b011001100111;
   9679: result <= 12'b011001100111;
   9680: result <= 12'b011001100111;
   9681: result <= 12'b011001100111;
   9682: result <= 12'b011001100111;
   9683: result <= 12'b011001100111;
   9684: result <= 12'b011001100111;
   9685: result <= 12'b011001100111;
   9686: result <= 12'b011001101000;
   9687: result <= 12'b011001101000;
   9688: result <= 12'b011001101000;
   9689: result <= 12'b011001101000;
   9690: result <= 12'b011001101000;
   9691: result <= 12'b011001101000;
   9692: result <= 12'b011001101000;
   9693: result <= 12'b011001101000;
   9694: result <= 12'b011001101000;
   9695: result <= 12'b011001101001;
   9696: result <= 12'b011001101001;
   9697: result <= 12'b011001101001;
   9698: result <= 12'b011001101001;
   9699: result <= 12'b011001101001;
   9700: result <= 12'b011001101001;
   9701: result <= 12'b011001101001;
   9702: result <= 12'b011001101001;
   9703: result <= 12'b011001101010;
   9704: result <= 12'b011001101010;
   9705: result <= 12'b011001101010;
   9706: result <= 12'b011001101010;
   9707: result <= 12'b011001101010;
   9708: result <= 12'b011001101010;
   9709: result <= 12'b011001101010;
   9710: result <= 12'b011001101010;
   9711: result <= 12'b011001101010;
   9712: result <= 12'b011001101011;
   9713: result <= 12'b011001101011;
   9714: result <= 12'b011001101011;
   9715: result <= 12'b011001101011;
   9716: result <= 12'b011001101011;
   9717: result <= 12'b011001101011;
   9718: result <= 12'b011001101011;
   9719: result <= 12'b011001101011;
   9720: result <= 12'b011001101100;
   9721: result <= 12'b011001101100;
   9722: result <= 12'b011001101100;
   9723: result <= 12'b011001101100;
   9724: result <= 12'b011001101100;
   9725: result <= 12'b011001101100;
   9726: result <= 12'b011001101100;
   9727: result <= 12'b011001101100;
   9728: result <= 12'b011001101100;
   9729: result <= 12'b011001101101;
   9730: result <= 12'b011001101101;
   9731: result <= 12'b011001101101;
   9732: result <= 12'b011001101101;
   9733: result <= 12'b011001101101;
   9734: result <= 12'b011001101101;
   9735: result <= 12'b011001101101;
   9736: result <= 12'b011001101101;
   9737: result <= 12'b011001101110;
   9738: result <= 12'b011001101110;
   9739: result <= 12'b011001101110;
   9740: result <= 12'b011001101110;
   9741: result <= 12'b011001101110;
   9742: result <= 12'b011001101110;
   9743: result <= 12'b011001101110;
   9744: result <= 12'b011001101110;
   9745: result <= 12'b011001101110;
   9746: result <= 12'b011001101111;
   9747: result <= 12'b011001101111;
   9748: result <= 12'b011001101111;
   9749: result <= 12'b011001101111;
   9750: result <= 12'b011001101111;
   9751: result <= 12'b011001101111;
   9752: result <= 12'b011001101111;
   9753: result <= 12'b011001101111;
   9754: result <= 12'b011001110000;
   9755: result <= 12'b011001110000;
   9756: result <= 12'b011001110000;
   9757: result <= 12'b011001110000;
   9758: result <= 12'b011001110000;
   9759: result <= 12'b011001110000;
   9760: result <= 12'b011001110000;
   9761: result <= 12'b011001110000;
   9762: result <= 12'b011001110000;
   9763: result <= 12'b011001110001;
   9764: result <= 12'b011001110001;
   9765: result <= 12'b011001110001;
   9766: result <= 12'b011001110001;
   9767: result <= 12'b011001110001;
   9768: result <= 12'b011001110001;
   9769: result <= 12'b011001110001;
   9770: result <= 12'b011001110001;
   9771: result <= 12'b011001110001;
   9772: result <= 12'b011001110010;
   9773: result <= 12'b011001110010;
   9774: result <= 12'b011001110010;
   9775: result <= 12'b011001110010;
   9776: result <= 12'b011001110010;
   9777: result <= 12'b011001110010;
   9778: result <= 12'b011001110010;
   9779: result <= 12'b011001110010;
   9780: result <= 12'b011001110011;
   9781: result <= 12'b011001110011;
   9782: result <= 12'b011001110011;
   9783: result <= 12'b011001110011;
   9784: result <= 12'b011001110011;
   9785: result <= 12'b011001110011;
   9786: result <= 12'b011001110011;
   9787: result <= 12'b011001110011;
   9788: result <= 12'b011001110011;
   9789: result <= 12'b011001110100;
   9790: result <= 12'b011001110100;
   9791: result <= 12'b011001110100;
   9792: result <= 12'b011001110100;
   9793: result <= 12'b011001110100;
   9794: result <= 12'b011001110100;
   9795: result <= 12'b011001110100;
   9796: result <= 12'b011001110100;
   9797: result <= 12'b011001110101;
   9798: result <= 12'b011001110101;
   9799: result <= 12'b011001110101;
   9800: result <= 12'b011001110101;
   9801: result <= 12'b011001110101;
   9802: result <= 12'b011001110101;
   9803: result <= 12'b011001110101;
   9804: result <= 12'b011001110101;
   9805: result <= 12'b011001110101;
   9806: result <= 12'b011001110110;
   9807: result <= 12'b011001110110;
   9808: result <= 12'b011001110110;
   9809: result <= 12'b011001110110;
   9810: result <= 12'b011001110110;
   9811: result <= 12'b011001110110;
   9812: result <= 12'b011001110110;
   9813: result <= 12'b011001110110;
   9814: result <= 12'b011001110110;
   9815: result <= 12'b011001110111;
   9816: result <= 12'b011001110111;
   9817: result <= 12'b011001110111;
   9818: result <= 12'b011001110111;
   9819: result <= 12'b011001110111;
   9820: result <= 12'b011001110111;
   9821: result <= 12'b011001110111;
   9822: result <= 12'b011001110111;
   9823: result <= 12'b011001111000;
   9824: result <= 12'b011001111000;
   9825: result <= 12'b011001111000;
   9826: result <= 12'b011001111000;
   9827: result <= 12'b011001111000;
   9828: result <= 12'b011001111000;
   9829: result <= 12'b011001111000;
   9830: result <= 12'b011001111000;
   9831: result <= 12'b011001111000;
   9832: result <= 12'b011001111001;
   9833: result <= 12'b011001111001;
   9834: result <= 12'b011001111001;
   9835: result <= 12'b011001111001;
   9836: result <= 12'b011001111001;
   9837: result <= 12'b011001111001;
   9838: result <= 12'b011001111001;
   9839: result <= 12'b011001111001;
   9840: result <= 12'b011001111001;
   9841: result <= 12'b011001111010;
   9842: result <= 12'b011001111010;
   9843: result <= 12'b011001111010;
   9844: result <= 12'b011001111010;
   9845: result <= 12'b011001111010;
   9846: result <= 12'b011001111010;
   9847: result <= 12'b011001111010;
   9848: result <= 12'b011001111010;
   9849: result <= 12'b011001111011;
   9850: result <= 12'b011001111011;
   9851: result <= 12'b011001111011;
   9852: result <= 12'b011001111011;
   9853: result <= 12'b011001111011;
   9854: result <= 12'b011001111011;
   9855: result <= 12'b011001111011;
   9856: result <= 12'b011001111011;
   9857: result <= 12'b011001111011;
   9858: result <= 12'b011001111100;
   9859: result <= 12'b011001111100;
   9860: result <= 12'b011001111100;
   9861: result <= 12'b011001111100;
   9862: result <= 12'b011001111100;
   9863: result <= 12'b011001111100;
   9864: result <= 12'b011001111100;
   9865: result <= 12'b011001111100;
   9866: result <= 12'b011001111100;
   9867: result <= 12'b011001111101;
   9868: result <= 12'b011001111101;
   9869: result <= 12'b011001111101;
   9870: result <= 12'b011001111101;
   9871: result <= 12'b011001111101;
   9872: result <= 12'b011001111101;
   9873: result <= 12'b011001111101;
   9874: result <= 12'b011001111101;
   9875: result <= 12'b011001111101;
   9876: result <= 12'b011001111110;
   9877: result <= 12'b011001111110;
   9878: result <= 12'b011001111110;
   9879: result <= 12'b011001111110;
   9880: result <= 12'b011001111110;
   9881: result <= 12'b011001111110;
   9882: result <= 12'b011001111110;
   9883: result <= 12'b011001111110;
   9884: result <= 12'b011001111111;
   9885: result <= 12'b011001111111;
   9886: result <= 12'b011001111111;
   9887: result <= 12'b011001111111;
   9888: result <= 12'b011001111111;
   9889: result <= 12'b011001111111;
   9890: result <= 12'b011001111111;
   9891: result <= 12'b011001111111;
   9892: result <= 12'b011001111111;
   9893: result <= 12'b011010000000;
   9894: result <= 12'b011010000000;
   9895: result <= 12'b011010000000;
   9896: result <= 12'b011010000000;
   9897: result <= 12'b011010000000;
   9898: result <= 12'b011010000000;
   9899: result <= 12'b011010000000;
   9900: result <= 12'b011010000000;
   9901: result <= 12'b011010000000;
   9902: result <= 12'b011010000001;
   9903: result <= 12'b011010000001;
   9904: result <= 12'b011010000001;
   9905: result <= 12'b011010000001;
   9906: result <= 12'b011010000001;
   9907: result <= 12'b011010000001;
   9908: result <= 12'b011010000001;
   9909: result <= 12'b011010000001;
   9910: result <= 12'b011010000010;
   9911: result <= 12'b011010000010;
   9912: result <= 12'b011010000010;
   9913: result <= 12'b011010000010;
   9914: result <= 12'b011010000010;
   9915: result <= 12'b011010000010;
   9916: result <= 12'b011010000010;
   9917: result <= 12'b011010000010;
   9918: result <= 12'b011010000010;
   9919: result <= 12'b011010000011;
   9920: result <= 12'b011010000011;
   9921: result <= 12'b011010000011;
   9922: result <= 12'b011010000011;
   9923: result <= 12'b011010000011;
   9924: result <= 12'b011010000011;
   9925: result <= 12'b011010000011;
   9926: result <= 12'b011010000011;
   9927: result <= 12'b011010000011;
   9928: result <= 12'b011010000100;
   9929: result <= 12'b011010000100;
   9930: result <= 12'b011010000100;
   9931: result <= 12'b011010000100;
   9932: result <= 12'b011010000100;
   9933: result <= 12'b011010000100;
   9934: result <= 12'b011010000100;
   9935: result <= 12'b011010000100;
   9936: result <= 12'b011010000100;
   9937: result <= 12'b011010000101;
   9938: result <= 12'b011010000101;
   9939: result <= 12'b011010000101;
   9940: result <= 12'b011010000101;
   9941: result <= 12'b011010000101;
   9942: result <= 12'b011010000101;
   9943: result <= 12'b011010000101;
   9944: result <= 12'b011010000101;
   9945: result <= 12'b011010000101;
   9946: result <= 12'b011010000110;
   9947: result <= 12'b011010000110;
   9948: result <= 12'b011010000110;
   9949: result <= 12'b011010000110;
   9950: result <= 12'b011010000110;
   9951: result <= 12'b011010000110;
   9952: result <= 12'b011010000110;
   9953: result <= 12'b011010000110;
   9954: result <= 12'b011010000111;
   9955: result <= 12'b011010000111;
   9956: result <= 12'b011010000111;
   9957: result <= 12'b011010000111;
   9958: result <= 12'b011010000111;
   9959: result <= 12'b011010000111;
   9960: result <= 12'b011010000111;
   9961: result <= 12'b011010000111;
   9962: result <= 12'b011010000111;
   9963: result <= 12'b011010001000;
   9964: result <= 12'b011010001000;
   9965: result <= 12'b011010001000;
   9966: result <= 12'b011010001000;
   9967: result <= 12'b011010001000;
   9968: result <= 12'b011010001000;
   9969: result <= 12'b011010001000;
   9970: result <= 12'b011010001000;
   9971: result <= 12'b011010001000;
   9972: result <= 12'b011010001001;
   9973: result <= 12'b011010001001;
   9974: result <= 12'b011010001001;
   9975: result <= 12'b011010001001;
   9976: result <= 12'b011010001001;
   9977: result <= 12'b011010001001;
   9978: result <= 12'b011010001001;
   9979: result <= 12'b011010001001;
   9980: result <= 12'b011010001001;
   9981: result <= 12'b011010001010;
   9982: result <= 12'b011010001010;
   9983: result <= 12'b011010001010;
   9984: result <= 12'b011010001010;
   9985: result <= 12'b011010001010;
   9986: result <= 12'b011010001010;
   9987: result <= 12'b011010001010;
   9988: result <= 12'b011010001010;
   9989: result <= 12'b011010001010;
   9990: result <= 12'b011010001011;
   9991: result <= 12'b011010001011;
   9992: result <= 12'b011010001011;
   9993: result <= 12'b011010001011;
   9994: result <= 12'b011010001011;
   9995: result <= 12'b011010001011;
   9996: result <= 12'b011010001011;
   9997: result <= 12'b011010001011;
   9998: result <= 12'b011010001011;
   9999: result <= 12'b011010001100;
   10000: result <= 12'b011010001100;
   10001: result <= 12'b011010001100;
   10002: result <= 12'b011010001100;
   10003: result <= 12'b011010001100;
   10004: result <= 12'b011010001100;
   10005: result <= 12'b011010001100;
   10006: result <= 12'b011010001100;
   10007: result <= 12'b011010001101;
   10008: result <= 12'b011010001101;
   10009: result <= 12'b011010001101;
   10010: result <= 12'b011010001101;
   10011: result <= 12'b011010001101;
   10012: result <= 12'b011010001101;
   10013: result <= 12'b011010001101;
   10014: result <= 12'b011010001101;
   10015: result <= 12'b011010001101;
   10016: result <= 12'b011010001110;
   10017: result <= 12'b011010001110;
   10018: result <= 12'b011010001110;
   10019: result <= 12'b011010001110;
   10020: result <= 12'b011010001110;
   10021: result <= 12'b011010001110;
   10022: result <= 12'b011010001110;
   10023: result <= 12'b011010001110;
   10024: result <= 12'b011010001110;
   10025: result <= 12'b011010001111;
   10026: result <= 12'b011010001111;
   10027: result <= 12'b011010001111;
   10028: result <= 12'b011010001111;
   10029: result <= 12'b011010001111;
   10030: result <= 12'b011010001111;
   10031: result <= 12'b011010001111;
   10032: result <= 12'b011010001111;
   10033: result <= 12'b011010001111;
   10034: result <= 12'b011010010000;
   10035: result <= 12'b011010010000;
   10036: result <= 12'b011010010000;
   10037: result <= 12'b011010010000;
   10038: result <= 12'b011010010000;
   10039: result <= 12'b011010010000;
   10040: result <= 12'b011010010000;
   10041: result <= 12'b011010010000;
   10042: result <= 12'b011010010000;
   10043: result <= 12'b011010010001;
   10044: result <= 12'b011010010001;
   10045: result <= 12'b011010010001;
   10046: result <= 12'b011010010001;
   10047: result <= 12'b011010010001;
   10048: result <= 12'b011010010001;
   10049: result <= 12'b011010010001;
   10050: result <= 12'b011010010001;
   10051: result <= 12'b011010010001;
   10052: result <= 12'b011010010010;
   10053: result <= 12'b011010010010;
   10054: result <= 12'b011010010010;
   10055: result <= 12'b011010010010;
   10056: result <= 12'b011010010010;
   10057: result <= 12'b011010010010;
   10058: result <= 12'b011010010010;
   10059: result <= 12'b011010010010;
   10060: result <= 12'b011010010010;
   10061: result <= 12'b011010010011;
   10062: result <= 12'b011010010011;
   10063: result <= 12'b011010010011;
   10064: result <= 12'b011010010011;
   10065: result <= 12'b011010010011;
   10066: result <= 12'b011010010011;
   10067: result <= 12'b011010010011;
   10068: result <= 12'b011010010011;
   10069: result <= 12'b011010010011;
   10070: result <= 12'b011010010100;
   10071: result <= 12'b011010010100;
   10072: result <= 12'b011010010100;
   10073: result <= 12'b011010010100;
   10074: result <= 12'b011010010100;
   10075: result <= 12'b011010010100;
   10076: result <= 12'b011010010100;
   10077: result <= 12'b011010010100;
   10078: result <= 12'b011010010100;
   10079: result <= 12'b011010010101;
   10080: result <= 12'b011010010101;
   10081: result <= 12'b011010010101;
   10082: result <= 12'b011010010101;
   10083: result <= 12'b011010010101;
   10084: result <= 12'b011010010101;
   10085: result <= 12'b011010010101;
   10086: result <= 12'b011010010101;
   10087: result <= 12'b011010010101;
   10088: result <= 12'b011010010110;
   10089: result <= 12'b011010010110;
   10090: result <= 12'b011010010110;
   10091: result <= 12'b011010010110;
   10092: result <= 12'b011010010110;
   10093: result <= 12'b011010010110;
   10094: result <= 12'b011010010110;
   10095: result <= 12'b011010010110;
   10096: result <= 12'b011010010110;
   10097: result <= 12'b011010010111;
   10098: result <= 12'b011010010111;
   10099: result <= 12'b011010010111;
   10100: result <= 12'b011010010111;
   10101: result <= 12'b011010010111;
   10102: result <= 12'b011010010111;
   10103: result <= 12'b011010010111;
   10104: result <= 12'b011010010111;
   10105: result <= 12'b011010010111;
   10106: result <= 12'b011010011000;
   10107: result <= 12'b011010011000;
   10108: result <= 12'b011010011000;
   10109: result <= 12'b011010011000;
   10110: result <= 12'b011010011000;
   10111: result <= 12'b011010011000;
   10112: result <= 12'b011010011000;
   10113: result <= 12'b011010011000;
   10114: result <= 12'b011010011000;
   10115: result <= 12'b011010011001;
   10116: result <= 12'b011010011001;
   10117: result <= 12'b011010011001;
   10118: result <= 12'b011010011001;
   10119: result <= 12'b011010011001;
   10120: result <= 12'b011010011001;
   10121: result <= 12'b011010011001;
   10122: result <= 12'b011010011001;
   10123: result <= 12'b011010011001;
   10124: result <= 12'b011010011010;
   10125: result <= 12'b011010011010;
   10126: result <= 12'b011010011010;
   10127: result <= 12'b011010011010;
   10128: result <= 12'b011010011010;
   10129: result <= 12'b011010011010;
   10130: result <= 12'b011010011010;
   10131: result <= 12'b011010011010;
   10132: result <= 12'b011010011010;
   10133: result <= 12'b011010011011;
   10134: result <= 12'b011010011011;
   10135: result <= 12'b011010011011;
   10136: result <= 12'b011010011011;
   10137: result <= 12'b011010011011;
   10138: result <= 12'b011010011011;
   10139: result <= 12'b011010011011;
   10140: result <= 12'b011010011011;
   10141: result <= 12'b011010011011;
   10142: result <= 12'b011010011100;
   10143: result <= 12'b011010011100;
   10144: result <= 12'b011010011100;
   10145: result <= 12'b011010011100;
   10146: result <= 12'b011010011100;
   10147: result <= 12'b011010011100;
   10148: result <= 12'b011010011100;
   10149: result <= 12'b011010011100;
   10150: result <= 12'b011010011100;
   10151: result <= 12'b011010011101;
   10152: result <= 12'b011010011101;
   10153: result <= 12'b011010011101;
   10154: result <= 12'b011010011101;
   10155: result <= 12'b011010011101;
   10156: result <= 12'b011010011101;
   10157: result <= 12'b011010011101;
   10158: result <= 12'b011010011101;
   10159: result <= 12'b011010011101;
   10160: result <= 12'b011010011110;
   10161: result <= 12'b011010011110;
   10162: result <= 12'b011010011110;
   10163: result <= 12'b011010011110;
   10164: result <= 12'b011010011110;
   10165: result <= 12'b011010011110;
   10166: result <= 12'b011010011110;
   10167: result <= 12'b011010011110;
   10168: result <= 12'b011010011110;
   10169: result <= 12'b011010011111;
   10170: result <= 12'b011010011111;
   10171: result <= 12'b011010011111;
   10172: result <= 12'b011010011111;
   10173: result <= 12'b011010011111;
   10174: result <= 12'b011010011111;
   10175: result <= 12'b011010011111;
   10176: result <= 12'b011010011111;
   10177: result <= 12'b011010011111;
   10178: result <= 12'b011010100000;
   10179: result <= 12'b011010100000;
   10180: result <= 12'b011010100000;
   10181: result <= 12'b011010100000;
   10182: result <= 12'b011010100000;
   10183: result <= 12'b011010100000;
   10184: result <= 12'b011010100000;
   10185: result <= 12'b011010100000;
   10186: result <= 12'b011010100000;
   10187: result <= 12'b011010100001;
   10188: result <= 12'b011010100001;
   10189: result <= 12'b011010100001;
   10190: result <= 12'b011010100001;
   10191: result <= 12'b011010100001;
   10192: result <= 12'b011010100001;
   10193: result <= 12'b011010100001;
   10194: result <= 12'b011010100001;
   10195: result <= 12'b011010100001;
   10196: result <= 12'b011010100010;
   10197: result <= 12'b011010100010;
   10198: result <= 12'b011010100010;
   10199: result <= 12'b011010100010;
   10200: result <= 12'b011010100010;
   10201: result <= 12'b011010100010;
   10202: result <= 12'b011010100010;
   10203: result <= 12'b011010100010;
   10204: result <= 12'b011010100010;
   10205: result <= 12'b011010100011;
   10206: result <= 12'b011010100011;
   10207: result <= 12'b011010100011;
   10208: result <= 12'b011010100011;
   10209: result <= 12'b011010100011;
   10210: result <= 12'b011010100011;
   10211: result <= 12'b011010100011;
   10212: result <= 12'b011010100011;
   10213: result <= 12'b011010100011;
   10214: result <= 12'b011010100100;
   10215: result <= 12'b011010100100;
   10216: result <= 12'b011010100100;
   10217: result <= 12'b011010100100;
   10218: result <= 12'b011010100100;
   10219: result <= 12'b011010100100;
   10220: result <= 12'b011010100100;
   10221: result <= 12'b011010100100;
   10222: result <= 12'b011010100100;
   10223: result <= 12'b011010100100;
   10224: result <= 12'b011010100101;
   10225: result <= 12'b011010100101;
   10226: result <= 12'b011010100101;
   10227: result <= 12'b011010100101;
   10228: result <= 12'b011010100101;
   10229: result <= 12'b011010100101;
   10230: result <= 12'b011010100101;
   10231: result <= 12'b011010100101;
   10232: result <= 12'b011010100101;
   10233: result <= 12'b011010100110;
   10234: result <= 12'b011010100110;
   10235: result <= 12'b011010100110;
   10236: result <= 12'b011010100110;
   10237: result <= 12'b011010100110;
   10238: result <= 12'b011010100110;
   10239: result <= 12'b011010100110;
   10240: result <= 12'b011010100110;
   10241: result <= 12'b011010100110;
   10242: result <= 12'b011010100111;
   10243: result <= 12'b011010100111;
   10244: result <= 12'b011010100111;
   10245: result <= 12'b011010100111;
   10246: result <= 12'b011010100111;
   10247: result <= 12'b011010100111;
   10248: result <= 12'b011010100111;
   10249: result <= 12'b011010100111;
   10250: result <= 12'b011010100111;
   10251: result <= 12'b011010101000;
   10252: result <= 12'b011010101000;
   10253: result <= 12'b011010101000;
   10254: result <= 12'b011010101000;
   10255: result <= 12'b011010101000;
   10256: result <= 12'b011010101000;
   10257: result <= 12'b011010101000;
   10258: result <= 12'b011010101000;
   10259: result <= 12'b011010101000;
   10260: result <= 12'b011010101001;
   10261: result <= 12'b011010101001;
   10262: result <= 12'b011010101001;
   10263: result <= 12'b011010101001;
   10264: result <= 12'b011010101001;
   10265: result <= 12'b011010101001;
   10266: result <= 12'b011010101001;
   10267: result <= 12'b011010101001;
   10268: result <= 12'b011010101001;
   10269: result <= 12'b011010101010;
   10270: result <= 12'b011010101010;
   10271: result <= 12'b011010101010;
   10272: result <= 12'b011010101010;
   10273: result <= 12'b011010101010;
   10274: result <= 12'b011010101010;
   10275: result <= 12'b011010101010;
   10276: result <= 12'b011010101010;
   10277: result <= 12'b011010101010;
   10278: result <= 12'b011010101010;
   10279: result <= 12'b011010101011;
   10280: result <= 12'b011010101011;
   10281: result <= 12'b011010101011;
   10282: result <= 12'b011010101011;
   10283: result <= 12'b011010101011;
   10284: result <= 12'b011010101011;
   10285: result <= 12'b011010101011;
   10286: result <= 12'b011010101011;
   10287: result <= 12'b011010101011;
   10288: result <= 12'b011010101100;
   10289: result <= 12'b011010101100;
   10290: result <= 12'b011010101100;
   10291: result <= 12'b011010101100;
   10292: result <= 12'b011010101100;
   10293: result <= 12'b011010101100;
   10294: result <= 12'b011010101100;
   10295: result <= 12'b011010101100;
   10296: result <= 12'b011010101100;
   10297: result <= 12'b011010101101;
   10298: result <= 12'b011010101101;
   10299: result <= 12'b011010101101;
   10300: result <= 12'b011010101101;
   10301: result <= 12'b011010101101;
   10302: result <= 12'b011010101101;
   10303: result <= 12'b011010101101;
   10304: result <= 12'b011010101101;
   10305: result <= 12'b011010101101;
   10306: result <= 12'b011010101110;
   10307: result <= 12'b011010101110;
   10308: result <= 12'b011010101110;
   10309: result <= 12'b011010101110;
   10310: result <= 12'b011010101110;
   10311: result <= 12'b011010101110;
   10312: result <= 12'b011010101110;
   10313: result <= 12'b011010101110;
   10314: result <= 12'b011010101110;
   10315: result <= 12'b011010101110;
   10316: result <= 12'b011010101111;
   10317: result <= 12'b011010101111;
   10318: result <= 12'b011010101111;
   10319: result <= 12'b011010101111;
   10320: result <= 12'b011010101111;
   10321: result <= 12'b011010101111;
   10322: result <= 12'b011010101111;
   10323: result <= 12'b011010101111;
   10324: result <= 12'b011010101111;
   10325: result <= 12'b011010110000;
   10326: result <= 12'b011010110000;
   10327: result <= 12'b011010110000;
   10328: result <= 12'b011010110000;
   10329: result <= 12'b011010110000;
   10330: result <= 12'b011010110000;
   10331: result <= 12'b011010110000;
   10332: result <= 12'b011010110000;
   10333: result <= 12'b011010110000;
   10334: result <= 12'b011010110001;
   10335: result <= 12'b011010110001;
   10336: result <= 12'b011010110001;
   10337: result <= 12'b011010110001;
   10338: result <= 12'b011010110001;
   10339: result <= 12'b011010110001;
   10340: result <= 12'b011010110001;
   10341: result <= 12'b011010110001;
   10342: result <= 12'b011010110001;
   10343: result <= 12'b011010110010;
   10344: result <= 12'b011010110010;
   10345: result <= 12'b011010110010;
   10346: result <= 12'b011010110010;
   10347: result <= 12'b011010110010;
   10348: result <= 12'b011010110010;
   10349: result <= 12'b011010110010;
   10350: result <= 12'b011010110010;
   10351: result <= 12'b011010110010;
   10352: result <= 12'b011010110010;
   10353: result <= 12'b011010110011;
   10354: result <= 12'b011010110011;
   10355: result <= 12'b011010110011;
   10356: result <= 12'b011010110011;
   10357: result <= 12'b011010110011;
   10358: result <= 12'b011010110011;
   10359: result <= 12'b011010110011;
   10360: result <= 12'b011010110011;
   10361: result <= 12'b011010110011;
   10362: result <= 12'b011010110100;
   10363: result <= 12'b011010110100;
   10364: result <= 12'b011010110100;
   10365: result <= 12'b011010110100;
   10366: result <= 12'b011010110100;
   10367: result <= 12'b011010110100;
   10368: result <= 12'b011010110100;
   10369: result <= 12'b011010110100;
   10370: result <= 12'b011010110100;
   10371: result <= 12'b011010110101;
   10372: result <= 12'b011010110101;
   10373: result <= 12'b011010110101;
   10374: result <= 12'b011010110101;
   10375: result <= 12'b011010110101;
   10376: result <= 12'b011010110101;
   10377: result <= 12'b011010110101;
   10378: result <= 12'b011010110101;
   10379: result <= 12'b011010110101;
   10380: result <= 12'b011010110101;
   10381: result <= 12'b011010110110;
   10382: result <= 12'b011010110110;
   10383: result <= 12'b011010110110;
   10384: result <= 12'b011010110110;
   10385: result <= 12'b011010110110;
   10386: result <= 12'b011010110110;
   10387: result <= 12'b011010110110;
   10388: result <= 12'b011010110110;
   10389: result <= 12'b011010110110;
   10390: result <= 12'b011010110111;
   10391: result <= 12'b011010110111;
   10392: result <= 12'b011010110111;
   10393: result <= 12'b011010110111;
   10394: result <= 12'b011010110111;
   10395: result <= 12'b011010110111;
   10396: result <= 12'b011010110111;
   10397: result <= 12'b011010110111;
   10398: result <= 12'b011010110111;
   10399: result <= 12'b011010110111;
   10400: result <= 12'b011010111000;
   10401: result <= 12'b011010111000;
   10402: result <= 12'b011010111000;
   10403: result <= 12'b011010111000;
   10404: result <= 12'b011010111000;
   10405: result <= 12'b011010111000;
   10406: result <= 12'b011010111000;
   10407: result <= 12'b011010111000;
   10408: result <= 12'b011010111000;
   10409: result <= 12'b011010111001;
   10410: result <= 12'b011010111001;
   10411: result <= 12'b011010111001;
   10412: result <= 12'b011010111001;
   10413: result <= 12'b011010111001;
   10414: result <= 12'b011010111001;
   10415: result <= 12'b011010111001;
   10416: result <= 12'b011010111001;
   10417: result <= 12'b011010111001;
   10418: result <= 12'b011010111010;
   10419: result <= 12'b011010111010;
   10420: result <= 12'b011010111010;
   10421: result <= 12'b011010111010;
   10422: result <= 12'b011010111010;
   10423: result <= 12'b011010111010;
   10424: result <= 12'b011010111010;
   10425: result <= 12'b011010111010;
   10426: result <= 12'b011010111010;
   10427: result <= 12'b011010111010;
   10428: result <= 12'b011010111011;
   10429: result <= 12'b011010111011;
   10430: result <= 12'b011010111011;
   10431: result <= 12'b011010111011;
   10432: result <= 12'b011010111011;
   10433: result <= 12'b011010111011;
   10434: result <= 12'b011010111011;
   10435: result <= 12'b011010111011;
   10436: result <= 12'b011010111011;
   10437: result <= 12'b011010111100;
   10438: result <= 12'b011010111100;
   10439: result <= 12'b011010111100;
   10440: result <= 12'b011010111100;
   10441: result <= 12'b011010111100;
   10442: result <= 12'b011010111100;
   10443: result <= 12'b011010111100;
   10444: result <= 12'b011010111100;
   10445: result <= 12'b011010111100;
   10446: result <= 12'b011010111100;
   10447: result <= 12'b011010111101;
   10448: result <= 12'b011010111101;
   10449: result <= 12'b011010111101;
   10450: result <= 12'b011010111101;
   10451: result <= 12'b011010111101;
   10452: result <= 12'b011010111101;
   10453: result <= 12'b011010111101;
   10454: result <= 12'b011010111101;
   10455: result <= 12'b011010111101;
   10456: result <= 12'b011010111110;
   10457: result <= 12'b011010111110;
   10458: result <= 12'b011010111110;
   10459: result <= 12'b011010111110;
   10460: result <= 12'b011010111110;
   10461: result <= 12'b011010111110;
   10462: result <= 12'b011010111110;
   10463: result <= 12'b011010111110;
   10464: result <= 12'b011010111110;
   10465: result <= 12'b011010111110;
   10466: result <= 12'b011010111111;
   10467: result <= 12'b011010111111;
   10468: result <= 12'b011010111111;
   10469: result <= 12'b011010111111;
   10470: result <= 12'b011010111111;
   10471: result <= 12'b011010111111;
   10472: result <= 12'b011010111111;
   10473: result <= 12'b011010111111;
   10474: result <= 12'b011010111111;
   10475: result <= 12'b011011000000;
   10476: result <= 12'b011011000000;
   10477: result <= 12'b011011000000;
   10478: result <= 12'b011011000000;
   10479: result <= 12'b011011000000;
   10480: result <= 12'b011011000000;
   10481: result <= 12'b011011000000;
   10482: result <= 12'b011011000000;
   10483: result <= 12'b011011000000;
   10484: result <= 12'b011011000000;
   10485: result <= 12'b011011000001;
   10486: result <= 12'b011011000001;
   10487: result <= 12'b011011000001;
   10488: result <= 12'b011011000001;
   10489: result <= 12'b011011000001;
   10490: result <= 12'b011011000001;
   10491: result <= 12'b011011000001;
   10492: result <= 12'b011011000001;
   10493: result <= 12'b011011000001;
   10494: result <= 12'b011011000010;
   10495: result <= 12'b011011000010;
   10496: result <= 12'b011011000010;
   10497: result <= 12'b011011000010;
   10498: result <= 12'b011011000010;
   10499: result <= 12'b011011000010;
   10500: result <= 12'b011011000010;
   10501: result <= 12'b011011000010;
   10502: result <= 12'b011011000010;
   10503: result <= 12'b011011000010;
   10504: result <= 12'b011011000011;
   10505: result <= 12'b011011000011;
   10506: result <= 12'b011011000011;
   10507: result <= 12'b011011000011;
   10508: result <= 12'b011011000011;
   10509: result <= 12'b011011000011;
   10510: result <= 12'b011011000011;
   10511: result <= 12'b011011000011;
   10512: result <= 12'b011011000011;
   10513: result <= 12'b011011000100;
   10514: result <= 12'b011011000100;
   10515: result <= 12'b011011000100;
   10516: result <= 12'b011011000100;
   10517: result <= 12'b011011000100;
   10518: result <= 12'b011011000100;
   10519: result <= 12'b011011000100;
   10520: result <= 12'b011011000100;
   10521: result <= 12'b011011000100;
   10522: result <= 12'b011011000100;
   10523: result <= 12'b011011000101;
   10524: result <= 12'b011011000101;
   10525: result <= 12'b011011000101;
   10526: result <= 12'b011011000101;
   10527: result <= 12'b011011000101;
   10528: result <= 12'b011011000101;
   10529: result <= 12'b011011000101;
   10530: result <= 12'b011011000101;
   10531: result <= 12'b011011000101;
   10532: result <= 12'b011011000110;
   10533: result <= 12'b011011000110;
   10534: result <= 12'b011011000110;
   10535: result <= 12'b011011000110;
   10536: result <= 12'b011011000110;
   10537: result <= 12'b011011000110;
   10538: result <= 12'b011011000110;
   10539: result <= 12'b011011000110;
   10540: result <= 12'b011011000110;
   10541: result <= 12'b011011000110;
   10542: result <= 12'b011011000111;
   10543: result <= 12'b011011000111;
   10544: result <= 12'b011011000111;
   10545: result <= 12'b011011000111;
   10546: result <= 12'b011011000111;
   10547: result <= 12'b011011000111;
   10548: result <= 12'b011011000111;
   10549: result <= 12'b011011000111;
   10550: result <= 12'b011011000111;
   10551: result <= 12'b011011001000;
   10552: result <= 12'b011011001000;
   10553: result <= 12'b011011001000;
   10554: result <= 12'b011011001000;
   10555: result <= 12'b011011001000;
   10556: result <= 12'b011011001000;
   10557: result <= 12'b011011001000;
   10558: result <= 12'b011011001000;
   10559: result <= 12'b011011001000;
   10560: result <= 12'b011011001000;
   10561: result <= 12'b011011001001;
   10562: result <= 12'b011011001001;
   10563: result <= 12'b011011001001;
   10564: result <= 12'b011011001001;
   10565: result <= 12'b011011001001;
   10566: result <= 12'b011011001001;
   10567: result <= 12'b011011001001;
   10568: result <= 12'b011011001001;
   10569: result <= 12'b011011001001;
   10570: result <= 12'b011011001001;
   10571: result <= 12'b011011001010;
   10572: result <= 12'b011011001010;
   10573: result <= 12'b011011001010;
   10574: result <= 12'b011011001010;
   10575: result <= 12'b011011001010;
   10576: result <= 12'b011011001010;
   10577: result <= 12'b011011001010;
   10578: result <= 12'b011011001010;
   10579: result <= 12'b011011001010;
   10580: result <= 12'b011011001011;
   10581: result <= 12'b011011001011;
   10582: result <= 12'b011011001011;
   10583: result <= 12'b011011001011;
   10584: result <= 12'b011011001011;
   10585: result <= 12'b011011001011;
   10586: result <= 12'b011011001011;
   10587: result <= 12'b011011001011;
   10588: result <= 12'b011011001011;
   10589: result <= 12'b011011001011;
   10590: result <= 12'b011011001100;
   10591: result <= 12'b011011001100;
   10592: result <= 12'b011011001100;
   10593: result <= 12'b011011001100;
   10594: result <= 12'b011011001100;
   10595: result <= 12'b011011001100;
   10596: result <= 12'b011011001100;
   10597: result <= 12'b011011001100;
   10598: result <= 12'b011011001100;
   10599: result <= 12'b011011001100;
   10600: result <= 12'b011011001101;
   10601: result <= 12'b011011001101;
   10602: result <= 12'b011011001101;
   10603: result <= 12'b011011001101;
   10604: result <= 12'b011011001101;
   10605: result <= 12'b011011001101;
   10606: result <= 12'b011011001101;
   10607: result <= 12'b011011001101;
   10608: result <= 12'b011011001101;
   10609: result <= 12'b011011001110;
   10610: result <= 12'b011011001110;
   10611: result <= 12'b011011001110;
   10612: result <= 12'b011011001110;
   10613: result <= 12'b011011001110;
   10614: result <= 12'b011011001110;
   10615: result <= 12'b011011001110;
   10616: result <= 12'b011011001110;
   10617: result <= 12'b011011001110;
   10618: result <= 12'b011011001110;
   10619: result <= 12'b011011001111;
   10620: result <= 12'b011011001111;
   10621: result <= 12'b011011001111;
   10622: result <= 12'b011011001111;
   10623: result <= 12'b011011001111;
   10624: result <= 12'b011011001111;
   10625: result <= 12'b011011001111;
   10626: result <= 12'b011011001111;
   10627: result <= 12'b011011001111;
   10628: result <= 12'b011011001111;
   10629: result <= 12'b011011010000;
   10630: result <= 12'b011011010000;
   10631: result <= 12'b011011010000;
   10632: result <= 12'b011011010000;
   10633: result <= 12'b011011010000;
   10634: result <= 12'b011011010000;
   10635: result <= 12'b011011010000;
   10636: result <= 12'b011011010000;
   10637: result <= 12'b011011010000;
   10638: result <= 12'b011011010001;
   10639: result <= 12'b011011010001;
   10640: result <= 12'b011011010001;
   10641: result <= 12'b011011010001;
   10642: result <= 12'b011011010001;
   10643: result <= 12'b011011010001;
   10644: result <= 12'b011011010001;
   10645: result <= 12'b011011010001;
   10646: result <= 12'b011011010001;
   10647: result <= 12'b011011010001;
   10648: result <= 12'b011011010010;
   10649: result <= 12'b011011010010;
   10650: result <= 12'b011011010010;
   10651: result <= 12'b011011010010;
   10652: result <= 12'b011011010010;
   10653: result <= 12'b011011010010;
   10654: result <= 12'b011011010010;
   10655: result <= 12'b011011010010;
   10656: result <= 12'b011011010010;
   10657: result <= 12'b011011010010;
   10658: result <= 12'b011011010011;
   10659: result <= 12'b011011010011;
   10660: result <= 12'b011011010011;
   10661: result <= 12'b011011010011;
   10662: result <= 12'b011011010011;
   10663: result <= 12'b011011010011;
   10664: result <= 12'b011011010011;
   10665: result <= 12'b011011010011;
   10666: result <= 12'b011011010011;
   10667: result <= 12'b011011010011;
   10668: result <= 12'b011011010100;
   10669: result <= 12'b011011010100;
   10670: result <= 12'b011011010100;
   10671: result <= 12'b011011010100;
   10672: result <= 12'b011011010100;
   10673: result <= 12'b011011010100;
   10674: result <= 12'b011011010100;
   10675: result <= 12'b011011010100;
   10676: result <= 12'b011011010100;
   10677: result <= 12'b011011010101;
   10678: result <= 12'b011011010101;
   10679: result <= 12'b011011010101;
   10680: result <= 12'b011011010101;
   10681: result <= 12'b011011010101;
   10682: result <= 12'b011011010101;
   10683: result <= 12'b011011010101;
   10684: result <= 12'b011011010101;
   10685: result <= 12'b011011010101;
   10686: result <= 12'b011011010101;
   10687: result <= 12'b011011010110;
   10688: result <= 12'b011011010110;
   10689: result <= 12'b011011010110;
   10690: result <= 12'b011011010110;
   10691: result <= 12'b011011010110;
   10692: result <= 12'b011011010110;
   10693: result <= 12'b011011010110;
   10694: result <= 12'b011011010110;
   10695: result <= 12'b011011010110;
   10696: result <= 12'b011011010110;
   10697: result <= 12'b011011010111;
   10698: result <= 12'b011011010111;
   10699: result <= 12'b011011010111;
   10700: result <= 12'b011011010111;
   10701: result <= 12'b011011010111;
   10702: result <= 12'b011011010111;
   10703: result <= 12'b011011010111;
   10704: result <= 12'b011011010111;
   10705: result <= 12'b011011010111;
   10706: result <= 12'b011011010111;
   10707: result <= 12'b011011011000;
   10708: result <= 12'b011011011000;
   10709: result <= 12'b011011011000;
   10710: result <= 12'b011011011000;
   10711: result <= 12'b011011011000;
   10712: result <= 12'b011011011000;
   10713: result <= 12'b011011011000;
   10714: result <= 12'b011011011000;
   10715: result <= 12'b011011011000;
   10716: result <= 12'b011011011000;
   10717: result <= 12'b011011011001;
   10718: result <= 12'b011011011001;
   10719: result <= 12'b011011011001;
   10720: result <= 12'b011011011001;
   10721: result <= 12'b011011011001;
   10722: result <= 12'b011011011001;
   10723: result <= 12'b011011011001;
   10724: result <= 12'b011011011001;
   10725: result <= 12'b011011011001;
   10726: result <= 12'b011011011001;
   10727: result <= 12'b011011011010;
   10728: result <= 12'b011011011010;
   10729: result <= 12'b011011011010;
   10730: result <= 12'b011011011010;
   10731: result <= 12'b011011011010;
   10732: result <= 12'b011011011010;
   10733: result <= 12'b011011011010;
   10734: result <= 12'b011011011010;
   10735: result <= 12'b011011011010;
   10736: result <= 12'b011011011011;
   10737: result <= 12'b011011011011;
   10738: result <= 12'b011011011011;
   10739: result <= 12'b011011011011;
   10740: result <= 12'b011011011011;
   10741: result <= 12'b011011011011;
   10742: result <= 12'b011011011011;
   10743: result <= 12'b011011011011;
   10744: result <= 12'b011011011011;
   10745: result <= 12'b011011011011;
   10746: result <= 12'b011011011100;
   10747: result <= 12'b011011011100;
   10748: result <= 12'b011011011100;
   10749: result <= 12'b011011011100;
   10750: result <= 12'b011011011100;
   10751: result <= 12'b011011011100;
   10752: result <= 12'b011011011100;
   10753: result <= 12'b011011011100;
   10754: result <= 12'b011011011100;
   10755: result <= 12'b011011011100;
   10756: result <= 12'b011011011101;
   10757: result <= 12'b011011011101;
   10758: result <= 12'b011011011101;
   10759: result <= 12'b011011011101;
   10760: result <= 12'b011011011101;
   10761: result <= 12'b011011011101;
   10762: result <= 12'b011011011101;
   10763: result <= 12'b011011011101;
   10764: result <= 12'b011011011101;
   10765: result <= 12'b011011011101;
   10766: result <= 12'b011011011110;
   10767: result <= 12'b011011011110;
   10768: result <= 12'b011011011110;
   10769: result <= 12'b011011011110;
   10770: result <= 12'b011011011110;
   10771: result <= 12'b011011011110;
   10772: result <= 12'b011011011110;
   10773: result <= 12'b011011011110;
   10774: result <= 12'b011011011110;
   10775: result <= 12'b011011011110;
   10776: result <= 12'b011011011111;
   10777: result <= 12'b011011011111;
   10778: result <= 12'b011011011111;
   10779: result <= 12'b011011011111;
   10780: result <= 12'b011011011111;
   10781: result <= 12'b011011011111;
   10782: result <= 12'b011011011111;
   10783: result <= 12'b011011011111;
   10784: result <= 12'b011011011111;
   10785: result <= 12'b011011011111;
   10786: result <= 12'b011011100000;
   10787: result <= 12'b011011100000;
   10788: result <= 12'b011011100000;
   10789: result <= 12'b011011100000;
   10790: result <= 12'b011011100000;
   10791: result <= 12'b011011100000;
   10792: result <= 12'b011011100000;
   10793: result <= 12'b011011100000;
   10794: result <= 12'b011011100000;
   10795: result <= 12'b011011100000;
   10796: result <= 12'b011011100001;
   10797: result <= 12'b011011100001;
   10798: result <= 12'b011011100001;
   10799: result <= 12'b011011100001;
   10800: result <= 12'b011011100001;
   10801: result <= 12'b011011100001;
   10802: result <= 12'b011011100001;
   10803: result <= 12'b011011100001;
   10804: result <= 12'b011011100001;
   10805: result <= 12'b011011100001;
   10806: result <= 12'b011011100010;
   10807: result <= 12'b011011100010;
   10808: result <= 12'b011011100010;
   10809: result <= 12'b011011100010;
   10810: result <= 12'b011011100010;
   10811: result <= 12'b011011100010;
   10812: result <= 12'b011011100010;
   10813: result <= 12'b011011100010;
   10814: result <= 12'b011011100010;
   10815: result <= 12'b011011100010;
   10816: result <= 12'b011011100011;
   10817: result <= 12'b011011100011;
   10818: result <= 12'b011011100011;
   10819: result <= 12'b011011100011;
   10820: result <= 12'b011011100011;
   10821: result <= 12'b011011100011;
   10822: result <= 12'b011011100011;
   10823: result <= 12'b011011100011;
   10824: result <= 12'b011011100011;
   10825: result <= 12'b011011100011;
   10826: result <= 12'b011011100100;
   10827: result <= 12'b011011100100;
   10828: result <= 12'b011011100100;
   10829: result <= 12'b011011100100;
   10830: result <= 12'b011011100100;
   10831: result <= 12'b011011100100;
   10832: result <= 12'b011011100100;
   10833: result <= 12'b011011100100;
   10834: result <= 12'b011011100100;
   10835: result <= 12'b011011100100;
   10836: result <= 12'b011011100101;
   10837: result <= 12'b011011100101;
   10838: result <= 12'b011011100101;
   10839: result <= 12'b011011100101;
   10840: result <= 12'b011011100101;
   10841: result <= 12'b011011100101;
   10842: result <= 12'b011011100101;
   10843: result <= 12'b011011100101;
   10844: result <= 12'b011011100101;
   10845: result <= 12'b011011100101;
   10846: result <= 12'b011011100110;
   10847: result <= 12'b011011100110;
   10848: result <= 12'b011011100110;
   10849: result <= 12'b011011100110;
   10850: result <= 12'b011011100110;
   10851: result <= 12'b011011100110;
   10852: result <= 12'b011011100110;
   10853: result <= 12'b011011100110;
   10854: result <= 12'b011011100110;
   10855: result <= 12'b011011100110;
   10856: result <= 12'b011011100111;
   10857: result <= 12'b011011100111;
   10858: result <= 12'b011011100111;
   10859: result <= 12'b011011100111;
   10860: result <= 12'b011011100111;
   10861: result <= 12'b011011100111;
   10862: result <= 12'b011011100111;
   10863: result <= 12'b011011100111;
   10864: result <= 12'b011011100111;
   10865: result <= 12'b011011100111;
   10866: result <= 12'b011011101000;
   10867: result <= 12'b011011101000;
   10868: result <= 12'b011011101000;
   10869: result <= 12'b011011101000;
   10870: result <= 12'b011011101000;
   10871: result <= 12'b011011101000;
   10872: result <= 12'b011011101000;
   10873: result <= 12'b011011101000;
   10874: result <= 12'b011011101000;
   10875: result <= 12'b011011101000;
   10876: result <= 12'b011011101001;
   10877: result <= 12'b011011101001;
   10878: result <= 12'b011011101001;
   10879: result <= 12'b011011101001;
   10880: result <= 12'b011011101001;
   10881: result <= 12'b011011101001;
   10882: result <= 12'b011011101001;
   10883: result <= 12'b011011101001;
   10884: result <= 12'b011011101001;
   10885: result <= 12'b011011101001;
   10886: result <= 12'b011011101010;
   10887: result <= 12'b011011101010;
   10888: result <= 12'b011011101010;
   10889: result <= 12'b011011101010;
   10890: result <= 12'b011011101010;
   10891: result <= 12'b011011101010;
   10892: result <= 12'b011011101010;
   10893: result <= 12'b011011101010;
   10894: result <= 12'b011011101010;
   10895: result <= 12'b011011101010;
   10896: result <= 12'b011011101010;
   10897: result <= 12'b011011101011;
   10898: result <= 12'b011011101011;
   10899: result <= 12'b011011101011;
   10900: result <= 12'b011011101011;
   10901: result <= 12'b011011101011;
   10902: result <= 12'b011011101011;
   10903: result <= 12'b011011101011;
   10904: result <= 12'b011011101011;
   10905: result <= 12'b011011101011;
   10906: result <= 12'b011011101011;
   10907: result <= 12'b011011101100;
   10908: result <= 12'b011011101100;
   10909: result <= 12'b011011101100;
   10910: result <= 12'b011011101100;
   10911: result <= 12'b011011101100;
   10912: result <= 12'b011011101100;
   10913: result <= 12'b011011101100;
   10914: result <= 12'b011011101100;
   10915: result <= 12'b011011101100;
   10916: result <= 12'b011011101100;
   10917: result <= 12'b011011101101;
   10918: result <= 12'b011011101101;
   10919: result <= 12'b011011101101;
   10920: result <= 12'b011011101101;
   10921: result <= 12'b011011101101;
   10922: result <= 12'b011011101101;
   10923: result <= 12'b011011101101;
   10924: result <= 12'b011011101101;
   10925: result <= 12'b011011101101;
   10926: result <= 12'b011011101101;
   10927: result <= 12'b011011101110;
   10928: result <= 12'b011011101110;
   10929: result <= 12'b011011101110;
   10930: result <= 12'b011011101110;
   10931: result <= 12'b011011101110;
   10932: result <= 12'b011011101110;
   10933: result <= 12'b011011101110;
   10934: result <= 12'b011011101110;
   10935: result <= 12'b011011101110;
   10936: result <= 12'b011011101110;
   10937: result <= 12'b011011101111;
   10938: result <= 12'b011011101111;
   10939: result <= 12'b011011101111;
   10940: result <= 12'b011011101111;
   10941: result <= 12'b011011101111;
   10942: result <= 12'b011011101111;
   10943: result <= 12'b011011101111;
   10944: result <= 12'b011011101111;
   10945: result <= 12'b011011101111;
   10946: result <= 12'b011011101111;
   10947: result <= 12'b011011110000;
   10948: result <= 12'b011011110000;
   10949: result <= 12'b011011110000;
   10950: result <= 12'b011011110000;
   10951: result <= 12'b011011110000;
   10952: result <= 12'b011011110000;
   10953: result <= 12'b011011110000;
   10954: result <= 12'b011011110000;
   10955: result <= 12'b011011110000;
   10956: result <= 12'b011011110000;
   10957: result <= 12'b011011110000;
   10958: result <= 12'b011011110001;
   10959: result <= 12'b011011110001;
   10960: result <= 12'b011011110001;
   10961: result <= 12'b011011110001;
   10962: result <= 12'b011011110001;
   10963: result <= 12'b011011110001;
   10964: result <= 12'b011011110001;
   10965: result <= 12'b011011110001;
   10966: result <= 12'b011011110001;
   10967: result <= 12'b011011110001;
   10968: result <= 12'b011011110010;
   10969: result <= 12'b011011110010;
   10970: result <= 12'b011011110010;
   10971: result <= 12'b011011110010;
   10972: result <= 12'b011011110010;
   10973: result <= 12'b011011110010;
   10974: result <= 12'b011011110010;
   10975: result <= 12'b011011110010;
   10976: result <= 12'b011011110010;
   10977: result <= 12'b011011110010;
   10978: result <= 12'b011011110011;
   10979: result <= 12'b011011110011;
   10980: result <= 12'b011011110011;
   10981: result <= 12'b011011110011;
   10982: result <= 12'b011011110011;
   10983: result <= 12'b011011110011;
   10984: result <= 12'b011011110011;
   10985: result <= 12'b011011110011;
   10986: result <= 12'b011011110011;
   10987: result <= 12'b011011110011;
   10988: result <= 12'b011011110011;
   10989: result <= 12'b011011110100;
   10990: result <= 12'b011011110100;
   10991: result <= 12'b011011110100;
   10992: result <= 12'b011011110100;
   10993: result <= 12'b011011110100;
   10994: result <= 12'b011011110100;
   10995: result <= 12'b011011110100;
   10996: result <= 12'b011011110100;
   10997: result <= 12'b011011110100;
   10998: result <= 12'b011011110100;
   10999: result <= 12'b011011110101;
   11000: result <= 12'b011011110101;
   11001: result <= 12'b011011110101;
   11002: result <= 12'b011011110101;
   11003: result <= 12'b011011110101;
   11004: result <= 12'b011011110101;
   11005: result <= 12'b011011110101;
   11006: result <= 12'b011011110101;
   11007: result <= 12'b011011110101;
   11008: result <= 12'b011011110101;
   11009: result <= 12'b011011110110;
   11010: result <= 12'b011011110110;
   11011: result <= 12'b011011110110;
   11012: result <= 12'b011011110110;
   11013: result <= 12'b011011110110;
   11014: result <= 12'b011011110110;
   11015: result <= 12'b011011110110;
   11016: result <= 12'b011011110110;
   11017: result <= 12'b011011110110;
   11018: result <= 12'b011011110110;
   11019: result <= 12'b011011110111;
   11020: result <= 12'b011011110111;
   11021: result <= 12'b011011110111;
   11022: result <= 12'b011011110111;
   11023: result <= 12'b011011110111;
   11024: result <= 12'b011011110111;
   11025: result <= 12'b011011110111;
   11026: result <= 12'b011011110111;
   11027: result <= 12'b011011110111;
   11028: result <= 12'b011011110111;
   11029: result <= 12'b011011110111;
   11030: result <= 12'b011011111000;
   11031: result <= 12'b011011111000;
   11032: result <= 12'b011011111000;
   11033: result <= 12'b011011111000;
   11034: result <= 12'b011011111000;
   11035: result <= 12'b011011111000;
   11036: result <= 12'b011011111000;
   11037: result <= 12'b011011111000;
   11038: result <= 12'b011011111000;
   11039: result <= 12'b011011111000;
   11040: result <= 12'b011011111001;
   11041: result <= 12'b011011111001;
   11042: result <= 12'b011011111001;
   11043: result <= 12'b011011111001;
   11044: result <= 12'b011011111001;
   11045: result <= 12'b011011111001;
   11046: result <= 12'b011011111001;
   11047: result <= 12'b011011111001;
   11048: result <= 12'b011011111001;
   11049: result <= 12'b011011111001;
   11050: result <= 12'b011011111001;
   11051: result <= 12'b011011111010;
   11052: result <= 12'b011011111010;
   11053: result <= 12'b011011111010;
   11054: result <= 12'b011011111010;
   11055: result <= 12'b011011111010;
   11056: result <= 12'b011011111010;
   11057: result <= 12'b011011111010;
   11058: result <= 12'b011011111010;
   11059: result <= 12'b011011111010;
   11060: result <= 12'b011011111010;
   11061: result <= 12'b011011111011;
   11062: result <= 12'b011011111011;
   11063: result <= 12'b011011111011;
   11064: result <= 12'b011011111011;
   11065: result <= 12'b011011111011;
   11066: result <= 12'b011011111011;
   11067: result <= 12'b011011111011;
   11068: result <= 12'b011011111011;
   11069: result <= 12'b011011111011;
   11070: result <= 12'b011011111011;
   11071: result <= 12'b011011111100;
   11072: result <= 12'b011011111100;
   11073: result <= 12'b011011111100;
   11074: result <= 12'b011011111100;
   11075: result <= 12'b011011111100;
   11076: result <= 12'b011011111100;
   11077: result <= 12'b011011111100;
   11078: result <= 12'b011011111100;
   11079: result <= 12'b011011111100;
   11080: result <= 12'b011011111100;
   11081: result <= 12'b011011111100;
   11082: result <= 12'b011011111101;
   11083: result <= 12'b011011111101;
   11084: result <= 12'b011011111101;
   11085: result <= 12'b011011111101;
   11086: result <= 12'b011011111101;
   11087: result <= 12'b011011111101;
   11088: result <= 12'b011011111101;
   11089: result <= 12'b011011111101;
   11090: result <= 12'b011011111101;
   11091: result <= 12'b011011111101;
   11092: result <= 12'b011011111110;
   11093: result <= 12'b011011111110;
   11094: result <= 12'b011011111110;
   11095: result <= 12'b011011111110;
   11096: result <= 12'b011011111110;
   11097: result <= 12'b011011111110;
   11098: result <= 12'b011011111110;
   11099: result <= 12'b011011111110;
   11100: result <= 12'b011011111110;
   11101: result <= 12'b011011111110;
   11102: result <= 12'b011011111110;
   11103: result <= 12'b011011111111;
   11104: result <= 12'b011011111111;
   11105: result <= 12'b011011111111;
   11106: result <= 12'b011011111111;
   11107: result <= 12'b011011111111;
   11108: result <= 12'b011011111111;
   11109: result <= 12'b011011111111;
   11110: result <= 12'b011011111111;
   11111: result <= 12'b011011111111;
   11112: result <= 12'b011011111111;
   11113: result <= 12'b011100000000;
   11114: result <= 12'b011100000000;
   11115: result <= 12'b011100000000;
   11116: result <= 12'b011100000000;
   11117: result <= 12'b011100000000;
   11118: result <= 12'b011100000000;
   11119: result <= 12'b011100000000;
   11120: result <= 12'b011100000000;
   11121: result <= 12'b011100000000;
   11122: result <= 12'b011100000000;
   11123: result <= 12'b011100000000;
   11124: result <= 12'b011100000001;
   11125: result <= 12'b011100000001;
   11126: result <= 12'b011100000001;
   11127: result <= 12'b011100000001;
   11128: result <= 12'b011100000001;
   11129: result <= 12'b011100000001;
   11130: result <= 12'b011100000001;
   11131: result <= 12'b011100000001;
   11132: result <= 12'b011100000001;
   11133: result <= 12'b011100000001;
   11134: result <= 12'b011100000010;
   11135: result <= 12'b011100000010;
   11136: result <= 12'b011100000010;
   11137: result <= 12'b011100000010;
   11138: result <= 12'b011100000010;
   11139: result <= 12'b011100000010;
   11140: result <= 12'b011100000010;
   11141: result <= 12'b011100000010;
   11142: result <= 12'b011100000010;
   11143: result <= 12'b011100000010;
   11144: result <= 12'b011100000010;
   11145: result <= 12'b011100000011;
   11146: result <= 12'b011100000011;
   11147: result <= 12'b011100000011;
   11148: result <= 12'b011100000011;
   11149: result <= 12'b011100000011;
   11150: result <= 12'b011100000011;
   11151: result <= 12'b011100000011;
   11152: result <= 12'b011100000011;
   11153: result <= 12'b011100000011;
   11154: result <= 12'b011100000011;
   11155: result <= 12'b011100000011;
   11156: result <= 12'b011100000100;
   11157: result <= 12'b011100000100;
   11158: result <= 12'b011100000100;
   11159: result <= 12'b011100000100;
   11160: result <= 12'b011100000100;
   11161: result <= 12'b011100000100;
   11162: result <= 12'b011100000100;
   11163: result <= 12'b011100000100;
   11164: result <= 12'b011100000100;
   11165: result <= 12'b011100000100;
   11166: result <= 12'b011100000101;
   11167: result <= 12'b011100000101;
   11168: result <= 12'b011100000101;
   11169: result <= 12'b011100000101;
   11170: result <= 12'b011100000101;
   11171: result <= 12'b011100000101;
   11172: result <= 12'b011100000101;
   11173: result <= 12'b011100000101;
   11174: result <= 12'b011100000101;
   11175: result <= 12'b011100000101;
   11176: result <= 12'b011100000101;
   11177: result <= 12'b011100000110;
   11178: result <= 12'b011100000110;
   11179: result <= 12'b011100000110;
   11180: result <= 12'b011100000110;
   11181: result <= 12'b011100000110;
   11182: result <= 12'b011100000110;
   11183: result <= 12'b011100000110;
   11184: result <= 12'b011100000110;
   11185: result <= 12'b011100000110;
   11186: result <= 12'b011100000110;
   11187: result <= 12'b011100000110;
   11188: result <= 12'b011100000111;
   11189: result <= 12'b011100000111;
   11190: result <= 12'b011100000111;
   11191: result <= 12'b011100000111;
   11192: result <= 12'b011100000111;
   11193: result <= 12'b011100000111;
   11194: result <= 12'b011100000111;
   11195: result <= 12'b011100000111;
   11196: result <= 12'b011100000111;
   11197: result <= 12'b011100000111;
   11198: result <= 12'b011100001000;
   11199: result <= 12'b011100001000;
   11200: result <= 12'b011100001000;
   11201: result <= 12'b011100001000;
   11202: result <= 12'b011100001000;
   11203: result <= 12'b011100001000;
   11204: result <= 12'b011100001000;
   11205: result <= 12'b011100001000;
   11206: result <= 12'b011100001000;
   11207: result <= 12'b011100001000;
   11208: result <= 12'b011100001000;
   11209: result <= 12'b011100001001;
   11210: result <= 12'b011100001001;
   11211: result <= 12'b011100001001;
   11212: result <= 12'b011100001001;
   11213: result <= 12'b011100001001;
   11214: result <= 12'b011100001001;
   11215: result <= 12'b011100001001;
   11216: result <= 12'b011100001001;
   11217: result <= 12'b011100001001;
   11218: result <= 12'b011100001001;
   11219: result <= 12'b011100001001;
   11220: result <= 12'b011100001010;
   11221: result <= 12'b011100001010;
   11222: result <= 12'b011100001010;
   11223: result <= 12'b011100001010;
   11224: result <= 12'b011100001010;
   11225: result <= 12'b011100001010;
   11226: result <= 12'b011100001010;
   11227: result <= 12'b011100001010;
   11228: result <= 12'b011100001010;
   11229: result <= 12'b011100001010;
   11230: result <= 12'b011100001011;
   11231: result <= 12'b011100001011;
   11232: result <= 12'b011100001011;
   11233: result <= 12'b011100001011;
   11234: result <= 12'b011100001011;
   11235: result <= 12'b011100001011;
   11236: result <= 12'b011100001011;
   11237: result <= 12'b011100001011;
   11238: result <= 12'b011100001011;
   11239: result <= 12'b011100001011;
   11240: result <= 12'b011100001011;
   11241: result <= 12'b011100001100;
   11242: result <= 12'b011100001100;
   11243: result <= 12'b011100001100;
   11244: result <= 12'b011100001100;
   11245: result <= 12'b011100001100;
   11246: result <= 12'b011100001100;
   11247: result <= 12'b011100001100;
   11248: result <= 12'b011100001100;
   11249: result <= 12'b011100001100;
   11250: result <= 12'b011100001100;
   11251: result <= 12'b011100001100;
   11252: result <= 12'b011100001101;
   11253: result <= 12'b011100001101;
   11254: result <= 12'b011100001101;
   11255: result <= 12'b011100001101;
   11256: result <= 12'b011100001101;
   11257: result <= 12'b011100001101;
   11258: result <= 12'b011100001101;
   11259: result <= 12'b011100001101;
   11260: result <= 12'b011100001101;
   11261: result <= 12'b011100001101;
   11262: result <= 12'b011100001101;
   11263: result <= 12'b011100001110;
   11264: result <= 12'b011100001110;
   11265: result <= 12'b011100001110;
   11266: result <= 12'b011100001110;
   11267: result <= 12'b011100001110;
   11268: result <= 12'b011100001110;
   11269: result <= 12'b011100001110;
   11270: result <= 12'b011100001110;
   11271: result <= 12'b011100001110;
   11272: result <= 12'b011100001110;
   11273: result <= 12'b011100001111;
   11274: result <= 12'b011100001111;
   11275: result <= 12'b011100001111;
   11276: result <= 12'b011100001111;
   11277: result <= 12'b011100001111;
   11278: result <= 12'b011100001111;
   11279: result <= 12'b011100001111;
   11280: result <= 12'b011100001111;
   11281: result <= 12'b011100001111;
   11282: result <= 12'b011100001111;
   11283: result <= 12'b011100001111;
   11284: result <= 12'b011100010000;
   11285: result <= 12'b011100010000;
   11286: result <= 12'b011100010000;
   11287: result <= 12'b011100010000;
   11288: result <= 12'b011100010000;
   11289: result <= 12'b011100010000;
   11290: result <= 12'b011100010000;
   11291: result <= 12'b011100010000;
   11292: result <= 12'b011100010000;
   11293: result <= 12'b011100010000;
   11294: result <= 12'b011100010000;
   11295: result <= 12'b011100010001;
   11296: result <= 12'b011100010001;
   11297: result <= 12'b011100010001;
   11298: result <= 12'b011100010001;
   11299: result <= 12'b011100010001;
   11300: result <= 12'b011100010001;
   11301: result <= 12'b011100010001;
   11302: result <= 12'b011100010001;
   11303: result <= 12'b011100010001;
   11304: result <= 12'b011100010001;
   11305: result <= 12'b011100010001;
   11306: result <= 12'b011100010010;
   11307: result <= 12'b011100010010;
   11308: result <= 12'b011100010010;
   11309: result <= 12'b011100010010;
   11310: result <= 12'b011100010010;
   11311: result <= 12'b011100010010;
   11312: result <= 12'b011100010010;
   11313: result <= 12'b011100010010;
   11314: result <= 12'b011100010010;
   11315: result <= 12'b011100010010;
   11316: result <= 12'b011100010010;
   11317: result <= 12'b011100010011;
   11318: result <= 12'b011100010011;
   11319: result <= 12'b011100010011;
   11320: result <= 12'b011100010011;
   11321: result <= 12'b011100010011;
   11322: result <= 12'b011100010011;
   11323: result <= 12'b011100010011;
   11324: result <= 12'b011100010011;
   11325: result <= 12'b011100010011;
   11326: result <= 12'b011100010011;
   11327: result <= 12'b011100010011;
   11328: result <= 12'b011100010100;
   11329: result <= 12'b011100010100;
   11330: result <= 12'b011100010100;
   11331: result <= 12'b011100010100;
   11332: result <= 12'b011100010100;
   11333: result <= 12'b011100010100;
   11334: result <= 12'b011100010100;
   11335: result <= 12'b011100010100;
   11336: result <= 12'b011100010100;
   11337: result <= 12'b011100010100;
   11338: result <= 12'b011100010100;
   11339: result <= 12'b011100010101;
   11340: result <= 12'b011100010101;
   11341: result <= 12'b011100010101;
   11342: result <= 12'b011100010101;
   11343: result <= 12'b011100010101;
   11344: result <= 12'b011100010101;
   11345: result <= 12'b011100010101;
   11346: result <= 12'b011100010101;
   11347: result <= 12'b011100010101;
   11348: result <= 12'b011100010101;
   11349: result <= 12'b011100010101;
   11350: result <= 12'b011100010110;
   11351: result <= 12'b011100010110;
   11352: result <= 12'b011100010110;
   11353: result <= 12'b011100010110;
   11354: result <= 12'b011100010110;
   11355: result <= 12'b011100010110;
   11356: result <= 12'b011100010110;
   11357: result <= 12'b011100010110;
   11358: result <= 12'b011100010110;
   11359: result <= 12'b011100010110;
   11360: result <= 12'b011100010110;
   11361: result <= 12'b011100010111;
   11362: result <= 12'b011100010111;
   11363: result <= 12'b011100010111;
   11364: result <= 12'b011100010111;
   11365: result <= 12'b011100010111;
   11366: result <= 12'b011100010111;
   11367: result <= 12'b011100010111;
   11368: result <= 12'b011100010111;
   11369: result <= 12'b011100010111;
   11370: result <= 12'b011100010111;
   11371: result <= 12'b011100010111;
   11372: result <= 12'b011100011000;
   11373: result <= 12'b011100011000;
   11374: result <= 12'b011100011000;
   11375: result <= 12'b011100011000;
   11376: result <= 12'b011100011000;
   11377: result <= 12'b011100011000;
   11378: result <= 12'b011100011000;
   11379: result <= 12'b011100011000;
   11380: result <= 12'b011100011000;
   11381: result <= 12'b011100011000;
   11382: result <= 12'b011100011000;
   11383: result <= 12'b011100011001;
   11384: result <= 12'b011100011001;
   11385: result <= 12'b011100011001;
   11386: result <= 12'b011100011001;
   11387: result <= 12'b011100011001;
   11388: result <= 12'b011100011001;
   11389: result <= 12'b011100011001;
   11390: result <= 12'b011100011001;
   11391: result <= 12'b011100011001;
   11392: result <= 12'b011100011001;
   11393: result <= 12'b011100011001;
   11394: result <= 12'b011100011010;
   11395: result <= 12'b011100011010;
   11396: result <= 12'b011100011010;
   11397: result <= 12'b011100011010;
   11398: result <= 12'b011100011010;
   11399: result <= 12'b011100011010;
   11400: result <= 12'b011100011010;
   11401: result <= 12'b011100011010;
   11402: result <= 12'b011100011010;
   11403: result <= 12'b011100011010;
   11404: result <= 12'b011100011010;
   11405: result <= 12'b011100011011;
   11406: result <= 12'b011100011011;
   11407: result <= 12'b011100011011;
   11408: result <= 12'b011100011011;
   11409: result <= 12'b011100011011;
   11410: result <= 12'b011100011011;
   11411: result <= 12'b011100011011;
   11412: result <= 12'b011100011011;
   11413: result <= 12'b011100011011;
   11414: result <= 12'b011100011011;
   11415: result <= 12'b011100011011;
   11416: result <= 12'b011100011100;
   11417: result <= 12'b011100011100;
   11418: result <= 12'b011100011100;
   11419: result <= 12'b011100011100;
   11420: result <= 12'b011100011100;
   11421: result <= 12'b011100011100;
   11422: result <= 12'b011100011100;
   11423: result <= 12'b011100011100;
   11424: result <= 12'b011100011100;
   11425: result <= 12'b011100011100;
   11426: result <= 12'b011100011100;
   11427: result <= 12'b011100011101;
   11428: result <= 12'b011100011101;
   11429: result <= 12'b011100011101;
   11430: result <= 12'b011100011101;
   11431: result <= 12'b011100011101;
   11432: result <= 12'b011100011101;
   11433: result <= 12'b011100011101;
   11434: result <= 12'b011100011101;
   11435: result <= 12'b011100011101;
   11436: result <= 12'b011100011101;
   11437: result <= 12'b011100011101;
   11438: result <= 12'b011100011110;
   11439: result <= 12'b011100011110;
   11440: result <= 12'b011100011110;
   11441: result <= 12'b011100011110;
   11442: result <= 12'b011100011110;
   11443: result <= 12'b011100011110;
   11444: result <= 12'b011100011110;
   11445: result <= 12'b011100011110;
   11446: result <= 12'b011100011110;
   11447: result <= 12'b011100011110;
   11448: result <= 12'b011100011110;
   11449: result <= 12'b011100011111;
   11450: result <= 12'b011100011111;
   11451: result <= 12'b011100011111;
   11452: result <= 12'b011100011111;
   11453: result <= 12'b011100011111;
   11454: result <= 12'b011100011111;
   11455: result <= 12'b011100011111;
   11456: result <= 12'b011100011111;
   11457: result <= 12'b011100011111;
   11458: result <= 12'b011100011111;
   11459: result <= 12'b011100011111;
   11460: result <= 12'b011100011111;
   11461: result <= 12'b011100100000;
   11462: result <= 12'b011100100000;
   11463: result <= 12'b011100100000;
   11464: result <= 12'b011100100000;
   11465: result <= 12'b011100100000;
   11466: result <= 12'b011100100000;
   11467: result <= 12'b011100100000;
   11468: result <= 12'b011100100000;
   11469: result <= 12'b011100100000;
   11470: result <= 12'b011100100000;
   11471: result <= 12'b011100100000;
   11472: result <= 12'b011100100001;
   11473: result <= 12'b011100100001;
   11474: result <= 12'b011100100001;
   11475: result <= 12'b011100100001;
   11476: result <= 12'b011100100001;
   11477: result <= 12'b011100100001;
   11478: result <= 12'b011100100001;
   11479: result <= 12'b011100100001;
   11480: result <= 12'b011100100001;
   11481: result <= 12'b011100100001;
   11482: result <= 12'b011100100001;
   11483: result <= 12'b011100100010;
   11484: result <= 12'b011100100010;
   11485: result <= 12'b011100100010;
   11486: result <= 12'b011100100010;
   11487: result <= 12'b011100100010;
   11488: result <= 12'b011100100010;
   11489: result <= 12'b011100100010;
   11490: result <= 12'b011100100010;
   11491: result <= 12'b011100100010;
   11492: result <= 12'b011100100010;
   11493: result <= 12'b011100100010;
   11494: result <= 12'b011100100011;
   11495: result <= 12'b011100100011;
   11496: result <= 12'b011100100011;
   11497: result <= 12'b011100100011;
   11498: result <= 12'b011100100011;
   11499: result <= 12'b011100100011;
   11500: result <= 12'b011100100011;
   11501: result <= 12'b011100100011;
   11502: result <= 12'b011100100011;
   11503: result <= 12'b011100100011;
   11504: result <= 12'b011100100011;
   11505: result <= 12'b011100100011;
   11506: result <= 12'b011100100100;
   11507: result <= 12'b011100100100;
   11508: result <= 12'b011100100100;
   11509: result <= 12'b011100100100;
   11510: result <= 12'b011100100100;
   11511: result <= 12'b011100100100;
   11512: result <= 12'b011100100100;
   11513: result <= 12'b011100100100;
   11514: result <= 12'b011100100100;
   11515: result <= 12'b011100100100;
   11516: result <= 12'b011100100100;
   11517: result <= 12'b011100100101;
   11518: result <= 12'b011100100101;
   11519: result <= 12'b011100100101;
   11520: result <= 12'b011100100101;
   11521: result <= 12'b011100100101;
   11522: result <= 12'b011100100101;
   11523: result <= 12'b011100100101;
   11524: result <= 12'b011100100101;
   11525: result <= 12'b011100100101;
   11526: result <= 12'b011100100101;
   11527: result <= 12'b011100100101;
   11528: result <= 12'b011100100110;
   11529: result <= 12'b011100100110;
   11530: result <= 12'b011100100110;
   11531: result <= 12'b011100100110;
   11532: result <= 12'b011100100110;
   11533: result <= 12'b011100100110;
   11534: result <= 12'b011100100110;
   11535: result <= 12'b011100100110;
   11536: result <= 12'b011100100110;
   11537: result <= 12'b011100100110;
   11538: result <= 12'b011100100110;
   11539: result <= 12'b011100100110;
   11540: result <= 12'b011100100111;
   11541: result <= 12'b011100100111;
   11542: result <= 12'b011100100111;
   11543: result <= 12'b011100100111;
   11544: result <= 12'b011100100111;
   11545: result <= 12'b011100100111;
   11546: result <= 12'b011100100111;
   11547: result <= 12'b011100100111;
   11548: result <= 12'b011100100111;
   11549: result <= 12'b011100100111;
   11550: result <= 12'b011100100111;
   11551: result <= 12'b011100101000;
   11552: result <= 12'b011100101000;
   11553: result <= 12'b011100101000;
   11554: result <= 12'b011100101000;
   11555: result <= 12'b011100101000;
   11556: result <= 12'b011100101000;
   11557: result <= 12'b011100101000;
   11558: result <= 12'b011100101000;
   11559: result <= 12'b011100101000;
   11560: result <= 12'b011100101000;
   11561: result <= 12'b011100101000;
   11562: result <= 12'b011100101001;
   11563: result <= 12'b011100101001;
   11564: result <= 12'b011100101001;
   11565: result <= 12'b011100101001;
   11566: result <= 12'b011100101001;
   11567: result <= 12'b011100101001;
   11568: result <= 12'b011100101001;
   11569: result <= 12'b011100101001;
   11570: result <= 12'b011100101001;
   11571: result <= 12'b011100101001;
   11572: result <= 12'b011100101001;
   11573: result <= 12'b011100101001;
   11574: result <= 12'b011100101010;
   11575: result <= 12'b011100101010;
   11576: result <= 12'b011100101010;
   11577: result <= 12'b011100101010;
   11578: result <= 12'b011100101010;
   11579: result <= 12'b011100101010;
   11580: result <= 12'b011100101010;
   11581: result <= 12'b011100101010;
   11582: result <= 12'b011100101010;
   11583: result <= 12'b011100101010;
   11584: result <= 12'b011100101010;
   11585: result <= 12'b011100101011;
   11586: result <= 12'b011100101011;
   11587: result <= 12'b011100101011;
   11588: result <= 12'b011100101011;
   11589: result <= 12'b011100101011;
   11590: result <= 12'b011100101011;
   11591: result <= 12'b011100101011;
   11592: result <= 12'b011100101011;
   11593: result <= 12'b011100101011;
   11594: result <= 12'b011100101011;
   11595: result <= 12'b011100101011;
   11596: result <= 12'b011100101011;
   11597: result <= 12'b011100101100;
   11598: result <= 12'b011100101100;
   11599: result <= 12'b011100101100;
   11600: result <= 12'b011100101100;
   11601: result <= 12'b011100101100;
   11602: result <= 12'b011100101100;
   11603: result <= 12'b011100101100;
   11604: result <= 12'b011100101100;
   11605: result <= 12'b011100101100;
   11606: result <= 12'b011100101100;
   11607: result <= 12'b011100101100;
   11608: result <= 12'b011100101101;
   11609: result <= 12'b011100101101;
   11610: result <= 12'b011100101101;
   11611: result <= 12'b011100101101;
   11612: result <= 12'b011100101101;
   11613: result <= 12'b011100101101;
   11614: result <= 12'b011100101101;
   11615: result <= 12'b011100101101;
   11616: result <= 12'b011100101101;
   11617: result <= 12'b011100101101;
   11618: result <= 12'b011100101101;
   11619: result <= 12'b011100101101;
   11620: result <= 12'b011100101110;
   11621: result <= 12'b011100101110;
   11622: result <= 12'b011100101110;
   11623: result <= 12'b011100101110;
   11624: result <= 12'b011100101110;
   11625: result <= 12'b011100101110;
   11626: result <= 12'b011100101110;
   11627: result <= 12'b011100101110;
   11628: result <= 12'b011100101110;
   11629: result <= 12'b011100101110;
   11630: result <= 12'b011100101110;
   11631: result <= 12'b011100101111;
   11632: result <= 12'b011100101111;
   11633: result <= 12'b011100101111;
   11634: result <= 12'b011100101111;
   11635: result <= 12'b011100101111;
   11636: result <= 12'b011100101111;
   11637: result <= 12'b011100101111;
   11638: result <= 12'b011100101111;
   11639: result <= 12'b011100101111;
   11640: result <= 12'b011100101111;
   11641: result <= 12'b011100101111;
   11642: result <= 12'b011100101111;
   11643: result <= 12'b011100110000;
   11644: result <= 12'b011100110000;
   11645: result <= 12'b011100110000;
   11646: result <= 12'b011100110000;
   11647: result <= 12'b011100110000;
   11648: result <= 12'b011100110000;
   11649: result <= 12'b011100110000;
   11650: result <= 12'b011100110000;
   11651: result <= 12'b011100110000;
   11652: result <= 12'b011100110000;
   11653: result <= 12'b011100110000;
   11654: result <= 12'b011100110001;
   11655: result <= 12'b011100110001;
   11656: result <= 12'b011100110001;
   11657: result <= 12'b011100110001;
   11658: result <= 12'b011100110001;
   11659: result <= 12'b011100110001;
   11660: result <= 12'b011100110001;
   11661: result <= 12'b011100110001;
   11662: result <= 12'b011100110001;
   11663: result <= 12'b011100110001;
   11664: result <= 12'b011100110001;
   11665: result <= 12'b011100110001;
   11666: result <= 12'b011100110010;
   11667: result <= 12'b011100110010;
   11668: result <= 12'b011100110010;
   11669: result <= 12'b011100110010;
   11670: result <= 12'b011100110010;
   11671: result <= 12'b011100110010;
   11672: result <= 12'b011100110010;
   11673: result <= 12'b011100110010;
   11674: result <= 12'b011100110010;
   11675: result <= 12'b011100110010;
   11676: result <= 12'b011100110010;
   11677: result <= 12'b011100110010;
   11678: result <= 12'b011100110011;
   11679: result <= 12'b011100110011;
   11680: result <= 12'b011100110011;
   11681: result <= 12'b011100110011;
   11682: result <= 12'b011100110011;
   11683: result <= 12'b011100110011;
   11684: result <= 12'b011100110011;
   11685: result <= 12'b011100110011;
   11686: result <= 12'b011100110011;
   11687: result <= 12'b011100110011;
   11688: result <= 12'b011100110011;
   11689: result <= 12'b011100110100;
   11690: result <= 12'b011100110100;
   11691: result <= 12'b011100110100;
   11692: result <= 12'b011100110100;
   11693: result <= 12'b011100110100;
   11694: result <= 12'b011100110100;
   11695: result <= 12'b011100110100;
   11696: result <= 12'b011100110100;
   11697: result <= 12'b011100110100;
   11698: result <= 12'b011100110100;
   11699: result <= 12'b011100110100;
   11700: result <= 12'b011100110100;
   11701: result <= 12'b011100110101;
   11702: result <= 12'b011100110101;
   11703: result <= 12'b011100110101;
   11704: result <= 12'b011100110101;
   11705: result <= 12'b011100110101;
   11706: result <= 12'b011100110101;
   11707: result <= 12'b011100110101;
   11708: result <= 12'b011100110101;
   11709: result <= 12'b011100110101;
   11710: result <= 12'b011100110101;
   11711: result <= 12'b011100110101;
   11712: result <= 12'b011100110101;
   11713: result <= 12'b011100110110;
   11714: result <= 12'b011100110110;
   11715: result <= 12'b011100110110;
   11716: result <= 12'b011100110110;
   11717: result <= 12'b011100110110;
   11718: result <= 12'b011100110110;
   11719: result <= 12'b011100110110;
   11720: result <= 12'b011100110110;
   11721: result <= 12'b011100110110;
   11722: result <= 12'b011100110110;
   11723: result <= 12'b011100110110;
   11724: result <= 12'b011100110110;
   11725: result <= 12'b011100110111;
   11726: result <= 12'b011100110111;
   11727: result <= 12'b011100110111;
   11728: result <= 12'b011100110111;
   11729: result <= 12'b011100110111;
   11730: result <= 12'b011100110111;
   11731: result <= 12'b011100110111;
   11732: result <= 12'b011100110111;
   11733: result <= 12'b011100110111;
   11734: result <= 12'b011100110111;
   11735: result <= 12'b011100110111;
   11736: result <= 12'b011100110111;
   11737: result <= 12'b011100111000;
   11738: result <= 12'b011100111000;
   11739: result <= 12'b011100111000;
   11740: result <= 12'b011100111000;
   11741: result <= 12'b011100111000;
   11742: result <= 12'b011100111000;
   11743: result <= 12'b011100111000;
   11744: result <= 12'b011100111000;
   11745: result <= 12'b011100111000;
   11746: result <= 12'b011100111000;
   11747: result <= 12'b011100111000;
   11748: result <= 12'b011100111001;
   11749: result <= 12'b011100111001;
   11750: result <= 12'b011100111001;
   11751: result <= 12'b011100111001;
   11752: result <= 12'b011100111001;
   11753: result <= 12'b011100111001;
   11754: result <= 12'b011100111001;
   11755: result <= 12'b011100111001;
   11756: result <= 12'b011100111001;
   11757: result <= 12'b011100111001;
   11758: result <= 12'b011100111001;
   11759: result <= 12'b011100111001;
   11760: result <= 12'b011100111010;
   11761: result <= 12'b011100111010;
   11762: result <= 12'b011100111010;
   11763: result <= 12'b011100111010;
   11764: result <= 12'b011100111010;
   11765: result <= 12'b011100111010;
   11766: result <= 12'b011100111010;
   11767: result <= 12'b011100111010;
   11768: result <= 12'b011100111010;
   11769: result <= 12'b011100111010;
   11770: result <= 12'b011100111010;
   11771: result <= 12'b011100111010;
   11772: result <= 12'b011100111011;
   11773: result <= 12'b011100111011;
   11774: result <= 12'b011100111011;
   11775: result <= 12'b011100111011;
   11776: result <= 12'b011100111011;
   11777: result <= 12'b011100111011;
   11778: result <= 12'b011100111011;
   11779: result <= 12'b011100111011;
   11780: result <= 12'b011100111011;
   11781: result <= 12'b011100111011;
   11782: result <= 12'b011100111011;
   11783: result <= 12'b011100111011;
   11784: result <= 12'b011100111100;
   11785: result <= 12'b011100111100;
   11786: result <= 12'b011100111100;
   11787: result <= 12'b011100111100;
   11788: result <= 12'b011100111100;
   11789: result <= 12'b011100111100;
   11790: result <= 12'b011100111100;
   11791: result <= 12'b011100111100;
   11792: result <= 12'b011100111100;
   11793: result <= 12'b011100111100;
   11794: result <= 12'b011100111100;
   11795: result <= 12'b011100111100;
   11796: result <= 12'b011100111101;
   11797: result <= 12'b011100111101;
   11798: result <= 12'b011100111101;
   11799: result <= 12'b011100111101;
   11800: result <= 12'b011100111101;
   11801: result <= 12'b011100111101;
   11802: result <= 12'b011100111101;
   11803: result <= 12'b011100111101;
   11804: result <= 12'b011100111101;
   11805: result <= 12'b011100111101;
   11806: result <= 12'b011100111101;
   11807: result <= 12'b011100111101;
   11808: result <= 12'b011100111110;
   11809: result <= 12'b011100111110;
   11810: result <= 12'b011100111110;
   11811: result <= 12'b011100111110;
   11812: result <= 12'b011100111110;
   11813: result <= 12'b011100111110;
   11814: result <= 12'b011100111110;
   11815: result <= 12'b011100111110;
   11816: result <= 12'b011100111110;
   11817: result <= 12'b011100111110;
   11818: result <= 12'b011100111110;
   11819: result <= 12'b011100111110;
   11820: result <= 12'b011100111111;
   11821: result <= 12'b011100111111;
   11822: result <= 12'b011100111111;
   11823: result <= 12'b011100111111;
   11824: result <= 12'b011100111111;
   11825: result <= 12'b011100111111;
   11826: result <= 12'b011100111111;
   11827: result <= 12'b011100111111;
   11828: result <= 12'b011100111111;
   11829: result <= 12'b011100111111;
   11830: result <= 12'b011100111111;
   11831: result <= 12'b011100111111;
   11832: result <= 12'b011101000000;
   11833: result <= 12'b011101000000;
   11834: result <= 12'b011101000000;
   11835: result <= 12'b011101000000;
   11836: result <= 12'b011101000000;
   11837: result <= 12'b011101000000;
   11838: result <= 12'b011101000000;
   11839: result <= 12'b011101000000;
   11840: result <= 12'b011101000000;
   11841: result <= 12'b011101000000;
   11842: result <= 12'b011101000000;
   11843: result <= 12'b011101000000;
   11844: result <= 12'b011101000001;
   11845: result <= 12'b011101000001;
   11846: result <= 12'b011101000001;
   11847: result <= 12'b011101000001;
   11848: result <= 12'b011101000001;
   11849: result <= 12'b011101000001;
   11850: result <= 12'b011101000001;
   11851: result <= 12'b011101000001;
   11852: result <= 12'b011101000001;
   11853: result <= 12'b011101000001;
   11854: result <= 12'b011101000001;
   11855: result <= 12'b011101000001;
   11856: result <= 12'b011101000010;
   11857: result <= 12'b011101000010;
   11858: result <= 12'b011101000010;
   11859: result <= 12'b011101000010;
   11860: result <= 12'b011101000010;
   11861: result <= 12'b011101000010;
   11862: result <= 12'b011101000010;
   11863: result <= 12'b011101000010;
   11864: result <= 12'b011101000010;
   11865: result <= 12'b011101000010;
   11866: result <= 12'b011101000010;
   11867: result <= 12'b011101000010;
   11868: result <= 12'b011101000011;
   11869: result <= 12'b011101000011;
   11870: result <= 12'b011101000011;
   11871: result <= 12'b011101000011;
   11872: result <= 12'b011101000011;
   11873: result <= 12'b011101000011;
   11874: result <= 12'b011101000011;
   11875: result <= 12'b011101000011;
   11876: result <= 12'b011101000011;
   11877: result <= 12'b011101000011;
   11878: result <= 12'b011101000011;
   11879: result <= 12'b011101000011;
   11880: result <= 12'b011101000100;
   11881: result <= 12'b011101000100;
   11882: result <= 12'b011101000100;
   11883: result <= 12'b011101000100;
   11884: result <= 12'b011101000100;
   11885: result <= 12'b011101000100;
   11886: result <= 12'b011101000100;
   11887: result <= 12'b011101000100;
   11888: result <= 12'b011101000100;
   11889: result <= 12'b011101000100;
   11890: result <= 12'b011101000100;
   11891: result <= 12'b011101000100;
   11892: result <= 12'b011101000100;
   11893: result <= 12'b011101000101;
   11894: result <= 12'b011101000101;
   11895: result <= 12'b011101000101;
   11896: result <= 12'b011101000101;
   11897: result <= 12'b011101000101;
   11898: result <= 12'b011101000101;
   11899: result <= 12'b011101000101;
   11900: result <= 12'b011101000101;
   11901: result <= 12'b011101000101;
   11902: result <= 12'b011101000101;
   11903: result <= 12'b011101000101;
   11904: result <= 12'b011101000101;
   11905: result <= 12'b011101000110;
   11906: result <= 12'b011101000110;
   11907: result <= 12'b011101000110;
   11908: result <= 12'b011101000110;
   11909: result <= 12'b011101000110;
   11910: result <= 12'b011101000110;
   11911: result <= 12'b011101000110;
   11912: result <= 12'b011101000110;
   11913: result <= 12'b011101000110;
   11914: result <= 12'b011101000110;
   11915: result <= 12'b011101000110;
   11916: result <= 12'b011101000110;
   11917: result <= 12'b011101000111;
   11918: result <= 12'b011101000111;
   11919: result <= 12'b011101000111;
   11920: result <= 12'b011101000111;
   11921: result <= 12'b011101000111;
   11922: result <= 12'b011101000111;
   11923: result <= 12'b011101000111;
   11924: result <= 12'b011101000111;
   11925: result <= 12'b011101000111;
   11926: result <= 12'b011101000111;
   11927: result <= 12'b011101000111;
   11928: result <= 12'b011101000111;
   11929: result <= 12'b011101001000;
   11930: result <= 12'b011101001000;
   11931: result <= 12'b011101001000;
   11932: result <= 12'b011101001000;
   11933: result <= 12'b011101001000;
   11934: result <= 12'b011101001000;
   11935: result <= 12'b011101001000;
   11936: result <= 12'b011101001000;
   11937: result <= 12'b011101001000;
   11938: result <= 12'b011101001000;
   11939: result <= 12'b011101001000;
   11940: result <= 12'b011101001000;
   11941: result <= 12'b011101001000;
   11942: result <= 12'b011101001001;
   11943: result <= 12'b011101001001;
   11944: result <= 12'b011101001001;
   11945: result <= 12'b011101001001;
   11946: result <= 12'b011101001001;
   11947: result <= 12'b011101001001;
   11948: result <= 12'b011101001001;
   11949: result <= 12'b011101001001;
   11950: result <= 12'b011101001001;
   11951: result <= 12'b011101001001;
   11952: result <= 12'b011101001001;
   11953: result <= 12'b011101001001;
   11954: result <= 12'b011101001010;
   11955: result <= 12'b011101001010;
   11956: result <= 12'b011101001010;
   11957: result <= 12'b011101001010;
   11958: result <= 12'b011101001010;
   11959: result <= 12'b011101001010;
   11960: result <= 12'b011101001010;
   11961: result <= 12'b011101001010;
   11962: result <= 12'b011101001010;
   11963: result <= 12'b011101001010;
   11964: result <= 12'b011101001010;
   11965: result <= 12'b011101001010;
   11966: result <= 12'b011101001011;
   11967: result <= 12'b011101001011;
   11968: result <= 12'b011101001011;
   11969: result <= 12'b011101001011;
   11970: result <= 12'b011101001011;
   11971: result <= 12'b011101001011;
   11972: result <= 12'b011101001011;
   11973: result <= 12'b011101001011;
   11974: result <= 12'b011101001011;
   11975: result <= 12'b011101001011;
   11976: result <= 12'b011101001011;
   11977: result <= 12'b011101001011;
   11978: result <= 12'b011101001011;
   11979: result <= 12'b011101001100;
   11980: result <= 12'b011101001100;
   11981: result <= 12'b011101001100;
   11982: result <= 12'b011101001100;
   11983: result <= 12'b011101001100;
   11984: result <= 12'b011101001100;
   11985: result <= 12'b011101001100;
   11986: result <= 12'b011101001100;
   11987: result <= 12'b011101001100;
   11988: result <= 12'b011101001100;
   11989: result <= 12'b011101001100;
   11990: result <= 12'b011101001100;
   11991: result <= 12'b011101001101;
   11992: result <= 12'b011101001101;
   11993: result <= 12'b011101001101;
   11994: result <= 12'b011101001101;
   11995: result <= 12'b011101001101;
   11996: result <= 12'b011101001101;
   11997: result <= 12'b011101001101;
   11998: result <= 12'b011101001101;
   11999: result <= 12'b011101001101;
   12000: result <= 12'b011101001101;
   12001: result <= 12'b011101001101;
   12002: result <= 12'b011101001101;
   12003: result <= 12'b011101001101;
   12004: result <= 12'b011101001110;
   12005: result <= 12'b011101001110;
   12006: result <= 12'b011101001110;
   12007: result <= 12'b011101001110;
   12008: result <= 12'b011101001110;
   12009: result <= 12'b011101001110;
   12010: result <= 12'b011101001110;
   12011: result <= 12'b011101001110;
   12012: result <= 12'b011101001110;
   12013: result <= 12'b011101001110;
   12014: result <= 12'b011101001110;
   12015: result <= 12'b011101001110;
   12016: result <= 12'b011101001111;
   12017: result <= 12'b011101001111;
   12018: result <= 12'b011101001111;
   12019: result <= 12'b011101001111;
   12020: result <= 12'b011101001111;
   12021: result <= 12'b011101001111;
   12022: result <= 12'b011101001111;
   12023: result <= 12'b011101001111;
   12024: result <= 12'b011101001111;
   12025: result <= 12'b011101001111;
   12026: result <= 12'b011101001111;
   12027: result <= 12'b011101001111;
   12028: result <= 12'b011101001111;
   12029: result <= 12'b011101010000;
   12030: result <= 12'b011101010000;
   12031: result <= 12'b011101010000;
   12032: result <= 12'b011101010000;
   12033: result <= 12'b011101010000;
   12034: result <= 12'b011101010000;
   12035: result <= 12'b011101010000;
   12036: result <= 12'b011101010000;
   12037: result <= 12'b011101010000;
   12038: result <= 12'b011101010000;
   12039: result <= 12'b011101010000;
   12040: result <= 12'b011101010000;
   12041: result <= 12'b011101010001;
   12042: result <= 12'b011101010001;
   12043: result <= 12'b011101010001;
   12044: result <= 12'b011101010001;
   12045: result <= 12'b011101010001;
   12046: result <= 12'b011101010001;
   12047: result <= 12'b011101010001;
   12048: result <= 12'b011101010001;
   12049: result <= 12'b011101010001;
   12050: result <= 12'b011101010001;
   12051: result <= 12'b011101010001;
   12052: result <= 12'b011101010001;
   12053: result <= 12'b011101010001;
   12054: result <= 12'b011101010010;
   12055: result <= 12'b011101010010;
   12056: result <= 12'b011101010010;
   12057: result <= 12'b011101010010;
   12058: result <= 12'b011101010010;
   12059: result <= 12'b011101010010;
   12060: result <= 12'b011101010010;
   12061: result <= 12'b011101010010;
   12062: result <= 12'b011101010010;
   12063: result <= 12'b011101010010;
   12064: result <= 12'b011101010010;
   12065: result <= 12'b011101010010;
   12066: result <= 12'b011101010010;
   12067: result <= 12'b011101010011;
   12068: result <= 12'b011101010011;
   12069: result <= 12'b011101010011;
   12070: result <= 12'b011101010011;
   12071: result <= 12'b011101010011;
   12072: result <= 12'b011101010011;
   12073: result <= 12'b011101010011;
   12074: result <= 12'b011101010011;
   12075: result <= 12'b011101010011;
   12076: result <= 12'b011101010011;
   12077: result <= 12'b011101010011;
   12078: result <= 12'b011101010011;
   12079: result <= 12'b011101010100;
   12080: result <= 12'b011101010100;
   12081: result <= 12'b011101010100;
   12082: result <= 12'b011101010100;
   12083: result <= 12'b011101010100;
   12084: result <= 12'b011101010100;
   12085: result <= 12'b011101010100;
   12086: result <= 12'b011101010100;
   12087: result <= 12'b011101010100;
   12088: result <= 12'b011101010100;
   12089: result <= 12'b011101010100;
   12090: result <= 12'b011101010100;
   12091: result <= 12'b011101010100;
   12092: result <= 12'b011101010101;
   12093: result <= 12'b011101010101;
   12094: result <= 12'b011101010101;
   12095: result <= 12'b011101010101;
   12096: result <= 12'b011101010101;
   12097: result <= 12'b011101010101;
   12098: result <= 12'b011101010101;
   12099: result <= 12'b011101010101;
   12100: result <= 12'b011101010101;
   12101: result <= 12'b011101010101;
   12102: result <= 12'b011101010101;
   12103: result <= 12'b011101010101;
   12104: result <= 12'b011101010101;
   12105: result <= 12'b011101010110;
   12106: result <= 12'b011101010110;
   12107: result <= 12'b011101010110;
   12108: result <= 12'b011101010110;
   12109: result <= 12'b011101010110;
   12110: result <= 12'b011101010110;
   12111: result <= 12'b011101010110;
   12112: result <= 12'b011101010110;
   12113: result <= 12'b011101010110;
   12114: result <= 12'b011101010110;
   12115: result <= 12'b011101010110;
   12116: result <= 12'b011101010110;
   12117: result <= 12'b011101010111;
   12118: result <= 12'b011101010111;
   12119: result <= 12'b011101010111;
   12120: result <= 12'b011101010111;
   12121: result <= 12'b011101010111;
   12122: result <= 12'b011101010111;
   12123: result <= 12'b011101010111;
   12124: result <= 12'b011101010111;
   12125: result <= 12'b011101010111;
   12126: result <= 12'b011101010111;
   12127: result <= 12'b011101010111;
   12128: result <= 12'b011101010111;
   12129: result <= 12'b011101010111;
   12130: result <= 12'b011101011000;
   12131: result <= 12'b011101011000;
   12132: result <= 12'b011101011000;
   12133: result <= 12'b011101011000;
   12134: result <= 12'b011101011000;
   12135: result <= 12'b011101011000;
   12136: result <= 12'b011101011000;
   12137: result <= 12'b011101011000;
   12138: result <= 12'b011101011000;
   12139: result <= 12'b011101011000;
   12140: result <= 12'b011101011000;
   12141: result <= 12'b011101011000;
   12142: result <= 12'b011101011000;
   12143: result <= 12'b011101011001;
   12144: result <= 12'b011101011001;
   12145: result <= 12'b011101011001;
   12146: result <= 12'b011101011001;
   12147: result <= 12'b011101011001;
   12148: result <= 12'b011101011001;
   12149: result <= 12'b011101011001;
   12150: result <= 12'b011101011001;
   12151: result <= 12'b011101011001;
   12152: result <= 12'b011101011001;
   12153: result <= 12'b011101011001;
   12154: result <= 12'b011101011001;
   12155: result <= 12'b011101011001;
   12156: result <= 12'b011101011010;
   12157: result <= 12'b011101011010;
   12158: result <= 12'b011101011010;
   12159: result <= 12'b011101011010;
   12160: result <= 12'b011101011010;
   12161: result <= 12'b011101011010;
   12162: result <= 12'b011101011010;
   12163: result <= 12'b011101011010;
   12164: result <= 12'b011101011010;
   12165: result <= 12'b011101011010;
   12166: result <= 12'b011101011010;
   12167: result <= 12'b011101011010;
   12168: result <= 12'b011101011010;
   12169: result <= 12'b011101011011;
   12170: result <= 12'b011101011011;
   12171: result <= 12'b011101011011;
   12172: result <= 12'b011101011011;
   12173: result <= 12'b011101011011;
   12174: result <= 12'b011101011011;
   12175: result <= 12'b011101011011;
   12176: result <= 12'b011101011011;
   12177: result <= 12'b011101011011;
   12178: result <= 12'b011101011011;
   12179: result <= 12'b011101011011;
   12180: result <= 12'b011101011011;
   12181: result <= 12'b011101011011;
   12182: result <= 12'b011101011100;
   12183: result <= 12'b011101011100;
   12184: result <= 12'b011101011100;
   12185: result <= 12'b011101011100;
   12186: result <= 12'b011101011100;
   12187: result <= 12'b011101011100;
   12188: result <= 12'b011101011100;
   12189: result <= 12'b011101011100;
   12190: result <= 12'b011101011100;
   12191: result <= 12'b011101011100;
   12192: result <= 12'b011101011100;
   12193: result <= 12'b011101011100;
   12194: result <= 12'b011101011100;
   12195: result <= 12'b011101011101;
   12196: result <= 12'b011101011101;
   12197: result <= 12'b011101011101;
   12198: result <= 12'b011101011101;
   12199: result <= 12'b011101011101;
   12200: result <= 12'b011101011101;
   12201: result <= 12'b011101011101;
   12202: result <= 12'b011101011101;
   12203: result <= 12'b011101011101;
   12204: result <= 12'b011101011101;
   12205: result <= 12'b011101011101;
   12206: result <= 12'b011101011101;
   12207: result <= 12'b011101011101;
   12208: result <= 12'b011101011110;
   12209: result <= 12'b011101011110;
   12210: result <= 12'b011101011110;
   12211: result <= 12'b011101011110;
   12212: result <= 12'b011101011110;
   12213: result <= 12'b011101011110;
   12214: result <= 12'b011101011110;
   12215: result <= 12'b011101011110;
   12216: result <= 12'b011101011110;
   12217: result <= 12'b011101011110;
   12218: result <= 12'b011101011110;
   12219: result <= 12'b011101011110;
   12220: result <= 12'b011101011110;
   12221: result <= 12'b011101011111;
   12222: result <= 12'b011101011111;
   12223: result <= 12'b011101011111;
   12224: result <= 12'b011101011111;
   12225: result <= 12'b011101011111;
   12226: result <= 12'b011101011111;
   12227: result <= 12'b011101011111;
   12228: result <= 12'b011101011111;
   12229: result <= 12'b011101011111;
   12230: result <= 12'b011101011111;
   12231: result <= 12'b011101011111;
   12232: result <= 12'b011101011111;
   12233: result <= 12'b011101011111;
   12234: result <= 12'b011101100000;
   12235: result <= 12'b011101100000;
   12236: result <= 12'b011101100000;
   12237: result <= 12'b011101100000;
   12238: result <= 12'b011101100000;
   12239: result <= 12'b011101100000;
   12240: result <= 12'b011101100000;
   12241: result <= 12'b011101100000;
   12242: result <= 12'b011101100000;
   12243: result <= 12'b011101100000;
   12244: result <= 12'b011101100000;
   12245: result <= 12'b011101100000;
   12246: result <= 12'b011101100000;
   12247: result <= 12'b011101100001;
   12248: result <= 12'b011101100001;
   12249: result <= 12'b011101100001;
   12250: result <= 12'b011101100001;
   12251: result <= 12'b011101100001;
   12252: result <= 12'b011101100001;
   12253: result <= 12'b011101100001;
   12254: result <= 12'b011101100001;
   12255: result <= 12'b011101100001;
   12256: result <= 12'b011101100001;
   12257: result <= 12'b011101100001;
   12258: result <= 12'b011101100001;
   12259: result <= 12'b011101100001;
   12260: result <= 12'b011101100001;
   12261: result <= 12'b011101100010;
   12262: result <= 12'b011101100010;
   12263: result <= 12'b011101100010;
   12264: result <= 12'b011101100010;
   12265: result <= 12'b011101100010;
   12266: result <= 12'b011101100010;
   12267: result <= 12'b011101100010;
   12268: result <= 12'b011101100010;
   12269: result <= 12'b011101100010;
   12270: result <= 12'b011101100010;
   12271: result <= 12'b011101100010;
   12272: result <= 12'b011101100010;
   12273: result <= 12'b011101100010;
   12274: result <= 12'b011101100011;
   12275: result <= 12'b011101100011;
   12276: result <= 12'b011101100011;
   12277: result <= 12'b011101100011;
   12278: result <= 12'b011101100011;
   12279: result <= 12'b011101100011;
   12280: result <= 12'b011101100011;
   12281: result <= 12'b011101100011;
   12282: result <= 12'b011101100011;
   12283: result <= 12'b011101100011;
   12284: result <= 12'b011101100011;
   12285: result <= 12'b011101100011;
   12286: result <= 12'b011101100011;
   12287: result <= 12'b011101100100;
   12288: result <= 12'b011101100100;
   12289: result <= 12'b011101100100;
   12290: result <= 12'b011101100100;
   12291: result <= 12'b011101100100;
   12292: result <= 12'b011101100100;
   12293: result <= 12'b011101100100;
   12294: result <= 12'b011101100100;
   12295: result <= 12'b011101100100;
   12296: result <= 12'b011101100100;
   12297: result <= 12'b011101100100;
   12298: result <= 12'b011101100100;
   12299: result <= 12'b011101100100;
   12300: result <= 12'b011101100101;
   12301: result <= 12'b011101100101;
   12302: result <= 12'b011101100101;
   12303: result <= 12'b011101100101;
   12304: result <= 12'b011101100101;
   12305: result <= 12'b011101100101;
   12306: result <= 12'b011101100101;
   12307: result <= 12'b011101100101;
   12308: result <= 12'b011101100101;
   12309: result <= 12'b011101100101;
   12310: result <= 12'b011101100101;
   12311: result <= 12'b011101100101;
   12312: result <= 12'b011101100101;
   12313: result <= 12'b011101100101;
   12314: result <= 12'b011101100110;
   12315: result <= 12'b011101100110;
   12316: result <= 12'b011101100110;
   12317: result <= 12'b011101100110;
   12318: result <= 12'b011101100110;
   12319: result <= 12'b011101100110;
   12320: result <= 12'b011101100110;
   12321: result <= 12'b011101100110;
   12322: result <= 12'b011101100110;
   12323: result <= 12'b011101100110;
   12324: result <= 12'b011101100110;
   12325: result <= 12'b011101100110;
   12326: result <= 12'b011101100110;
   12327: result <= 12'b011101100111;
   12328: result <= 12'b011101100111;
   12329: result <= 12'b011101100111;
   12330: result <= 12'b011101100111;
   12331: result <= 12'b011101100111;
   12332: result <= 12'b011101100111;
   12333: result <= 12'b011101100111;
   12334: result <= 12'b011101100111;
   12335: result <= 12'b011101100111;
   12336: result <= 12'b011101100111;
   12337: result <= 12'b011101100111;
   12338: result <= 12'b011101100111;
   12339: result <= 12'b011101100111;
   12340: result <= 12'b011101100111;
   12341: result <= 12'b011101101000;
   12342: result <= 12'b011101101000;
   12343: result <= 12'b011101101000;
   12344: result <= 12'b011101101000;
   12345: result <= 12'b011101101000;
   12346: result <= 12'b011101101000;
   12347: result <= 12'b011101101000;
   12348: result <= 12'b011101101000;
   12349: result <= 12'b011101101000;
   12350: result <= 12'b011101101000;
   12351: result <= 12'b011101101000;
   12352: result <= 12'b011101101000;
   12353: result <= 12'b011101101000;
   12354: result <= 12'b011101101001;
   12355: result <= 12'b011101101001;
   12356: result <= 12'b011101101001;
   12357: result <= 12'b011101101001;
   12358: result <= 12'b011101101001;
   12359: result <= 12'b011101101001;
   12360: result <= 12'b011101101001;
   12361: result <= 12'b011101101001;
   12362: result <= 12'b011101101001;
   12363: result <= 12'b011101101001;
   12364: result <= 12'b011101101001;
   12365: result <= 12'b011101101001;
   12366: result <= 12'b011101101001;
   12367: result <= 12'b011101101001;
   12368: result <= 12'b011101101010;
   12369: result <= 12'b011101101010;
   12370: result <= 12'b011101101010;
   12371: result <= 12'b011101101010;
   12372: result <= 12'b011101101010;
   12373: result <= 12'b011101101010;
   12374: result <= 12'b011101101010;
   12375: result <= 12'b011101101010;
   12376: result <= 12'b011101101010;
   12377: result <= 12'b011101101010;
   12378: result <= 12'b011101101010;
   12379: result <= 12'b011101101010;
   12380: result <= 12'b011101101010;
   12381: result <= 12'b011101101011;
   12382: result <= 12'b011101101011;
   12383: result <= 12'b011101101011;
   12384: result <= 12'b011101101011;
   12385: result <= 12'b011101101011;
   12386: result <= 12'b011101101011;
   12387: result <= 12'b011101101011;
   12388: result <= 12'b011101101011;
   12389: result <= 12'b011101101011;
   12390: result <= 12'b011101101011;
   12391: result <= 12'b011101101011;
   12392: result <= 12'b011101101011;
   12393: result <= 12'b011101101011;
   12394: result <= 12'b011101101011;
   12395: result <= 12'b011101101100;
   12396: result <= 12'b011101101100;
   12397: result <= 12'b011101101100;
   12398: result <= 12'b011101101100;
   12399: result <= 12'b011101101100;
   12400: result <= 12'b011101101100;
   12401: result <= 12'b011101101100;
   12402: result <= 12'b011101101100;
   12403: result <= 12'b011101101100;
   12404: result <= 12'b011101101100;
   12405: result <= 12'b011101101100;
   12406: result <= 12'b011101101100;
   12407: result <= 12'b011101101100;
   12408: result <= 12'b011101101100;
   12409: result <= 12'b011101101101;
   12410: result <= 12'b011101101101;
   12411: result <= 12'b011101101101;
   12412: result <= 12'b011101101101;
   12413: result <= 12'b011101101101;
   12414: result <= 12'b011101101101;
   12415: result <= 12'b011101101101;
   12416: result <= 12'b011101101101;
   12417: result <= 12'b011101101101;
   12418: result <= 12'b011101101101;
   12419: result <= 12'b011101101101;
   12420: result <= 12'b011101101101;
   12421: result <= 12'b011101101101;
   12422: result <= 12'b011101101110;
   12423: result <= 12'b011101101110;
   12424: result <= 12'b011101101110;
   12425: result <= 12'b011101101110;
   12426: result <= 12'b011101101110;
   12427: result <= 12'b011101101110;
   12428: result <= 12'b011101101110;
   12429: result <= 12'b011101101110;
   12430: result <= 12'b011101101110;
   12431: result <= 12'b011101101110;
   12432: result <= 12'b011101101110;
   12433: result <= 12'b011101101110;
   12434: result <= 12'b011101101110;
   12435: result <= 12'b011101101110;
   12436: result <= 12'b011101101111;
   12437: result <= 12'b011101101111;
   12438: result <= 12'b011101101111;
   12439: result <= 12'b011101101111;
   12440: result <= 12'b011101101111;
   12441: result <= 12'b011101101111;
   12442: result <= 12'b011101101111;
   12443: result <= 12'b011101101111;
   12444: result <= 12'b011101101111;
   12445: result <= 12'b011101101111;
   12446: result <= 12'b011101101111;
   12447: result <= 12'b011101101111;
   12448: result <= 12'b011101101111;
   12449: result <= 12'b011101101111;
   12450: result <= 12'b011101110000;
   12451: result <= 12'b011101110000;
   12452: result <= 12'b011101110000;
   12453: result <= 12'b011101110000;
   12454: result <= 12'b011101110000;
   12455: result <= 12'b011101110000;
   12456: result <= 12'b011101110000;
   12457: result <= 12'b011101110000;
   12458: result <= 12'b011101110000;
   12459: result <= 12'b011101110000;
   12460: result <= 12'b011101110000;
   12461: result <= 12'b011101110000;
   12462: result <= 12'b011101110000;
   12463: result <= 12'b011101110000;
   12464: result <= 12'b011101110001;
   12465: result <= 12'b011101110001;
   12466: result <= 12'b011101110001;
   12467: result <= 12'b011101110001;
   12468: result <= 12'b011101110001;
   12469: result <= 12'b011101110001;
   12470: result <= 12'b011101110001;
   12471: result <= 12'b011101110001;
   12472: result <= 12'b011101110001;
   12473: result <= 12'b011101110001;
   12474: result <= 12'b011101110001;
   12475: result <= 12'b011101110001;
   12476: result <= 12'b011101110001;
   12477: result <= 12'b011101110001;
   12478: result <= 12'b011101110010;
   12479: result <= 12'b011101110010;
   12480: result <= 12'b011101110010;
   12481: result <= 12'b011101110010;
   12482: result <= 12'b011101110010;
   12483: result <= 12'b011101110010;
   12484: result <= 12'b011101110010;
   12485: result <= 12'b011101110010;
   12486: result <= 12'b011101110010;
   12487: result <= 12'b011101110010;
   12488: result <= 12'b011101110010;
   12489: result <= 12'b011101110010;
   12490: result <= 12'b011101110010;
   12491: result <= 12'b011101110010;
   12492: result <= 12'b011101110011;
   12493: result <= 12'b011101110011;
   12494: result <= 12'b011101110011;
   12495: result <= 12'b011101110011;
   12496: result <= 12'b011101110011;
   12497: result <= 12'b011101110011;
   12498: result <= 12'b011101110011;
   12499: result <= 12'b011101110011;
   12500: result <= 12'b011101110011;
   12501: result <= 12'b011101110011;
   12502: result <= 12'b011101110011;
   12503: result <= 12'b011101110011;
   12504: result <= 12'b011101110011;
   12505: result <= 12'b011101110011;
   12506: result <= 12'b011101110100;
   12507: result <= 12'b011101110100;
   12508: result <= 12'b011101110100;
   12509: result <= 12'b011101110100;
   12510: result <= 12'b011101110100;
   12511: result <= 12'b011101110100;
   12512: result <= 12'b011101110100;
   12513: result <= 12'b011101110100;
   12514: result <= 12'b011101110100;
   12515: result <= 12'b011101110100;
   12516: result <= 12'b011101110100;
   12517: result <= 12'b011101110100;
   12518: result <= 12'b011101110100;
   12519: result <= 12'b011101110100;
   12520: result <= 12'b011101110101;
   12521: result <= 12'b011101110101;
   12522: result <= 12'b011101110101;
   12523: result <= 12'b011101110101;
   12524: result <= 12'b011101110101;
   12525: result <= 12'b011101110101;
   12526: result <= 12'b011101110101;
   12527: result <= 12'b011101110101;
   12528: result <= 12'b011101110101;
   12529: result <= 12'b011101110101;
   12530: result <= 12'b011101110101;
   12531: result <= 12'b011101110101;
   12532: result <= 12'b011101110101;
   12533: result <= 12'b011101110101;
   12534: result <= 12'b011101110110;
   12535: result <= 12'b011101110110;
   12536: result <= 12'b011101110110;
   12537: result <= 12'b011101110110;
   12538: result <= 12'b011101110110;
   12539: result <= 12'b011101110110;
   12540: result <= 12'b011101110110;
   12541: result <= 12'b011101110110;
   12542: result <= 12'b011101110110;
   12543: result <= 12'b011101110110;
   12544: result <= 12'b011101110110;
   12545: result <= 12'b011101110110;
   12546: result <= 12'b011101110110;
   12547: result <= 12'b011101110110;
   12548: result <= 12'b011101110111;
   12549: result <= 12'b011101110111;
   12550: result <= 12'b011101110111;
   12551: result <= 12'b011101110111;
   12552: result <= 12'b011101110111;
   12553: result <= 12'b011101110111;
   12554: result <= 12'b011101110111;
   12555: result <= 12'b011101110111;
   12556: result <= 12'b011101110111;
   12557: result <= 12'b011101110111;
   12558: result <= 12'b011101110111;
   12559: result <= 12'b011101110111;
   12560: result <= 12'b011101110111;
   12561: result <= 12'b011101110111;
   12562: result <= 12'b011101111000;
   12563: result <= 12'b011101111000;
   12564: result <= 12'b011101111000;
   12565: result <= 12'b011101111000;
   12566: result <= 12'b011101111000;
   12567: result <= 12'b011101111000;
   12568: result <= 12'b011101111000;
   12569: result <= 12'b011101111000;
   12570: result <= 12'b011101111000;
   12571: result <= 12'b011101111000;
   12572: result <= 12'b011101111000;
   12573: result <= 12'b011101111000;
   12574: result <= 12'b011101111000;
   12575: result <= 12'b011101111000;
   12576: result <= 12'b011101111001;
   12577: result <= 12'b011101111001;
   12578: result <= 12'b011101111001;
   12579: result <= 12'b011101111001;
   12580: result <= 12'b011101111001;
   12581: result <= 12'b011101111001;
   12582: result <= 12'b011101111001;
   12583: result <= 12'b011101111001;
   12584: result <= 12'b011101111001;
   12585: result <= 12'b011101111001;
   12586: result <= 12'b011101111001;
   12587: result <= 12'b011101111001;
   12588: result <= 12'b011101111001;
   12589: result <= 12'b011101111001;
   12590: result <= 12'b011101111010;
   12591: result <= 12'b011101111010;
   12592: result <= 12'b011101111010;
   12593: result <= 12'b011101111010;
   12594: result <= 12'b011101111010;
   12595: result <= 12'b011101111010;
   12596: result <= 12'b011101111010;
   12597: result <= 12'b011101111010;
   12598: result <= 12'b011101111010;
   12599: result <= 12'b011101111010;
   12600: result <= 12'b011101111010;
   12601: result <= 12'b011101111010;
   12602: result <= 12'b011101111010;
   12603: result <= 12'b011101111010;
   12604: result <= 12'b011101111010;
   12605: result <= 12'b011101111011;
   12606: result <= 12'b011101111011;
   12607: result <= 12'b011101111011;
   12608: result <= 12'b011101111011;
   12609: result <= 12'b011101111011;
   12610: result <= 12'b011101111011;
   12611: result <= 12'b011101111011;
   12612: result <= 12'b011101111011;
   12613: result <= 12'b011101111011;
   12614: result <= 12'b011101111011;
   12615: result <= 12'b011101111011;
   12616: result <= 12'b011101111011;
   12617: result <= 12'b011101111011;
   12618: result <= 12'b011101111011;
   12619: result <= 12'b011101111100;
   12620: result <= 12'b011101111100;
   12621: result <= 12'b011101111100;
   12622: result <= 12'b011101111100;
   12623: result <= 12'b011101111100;
   12624: result <= 12'b011101111100;
   12625: result <= 12'b011101111100;
   12626: result <= 12'b011101111100;
   12627: result <= 12'b011101111100;
   12628: result <= 12'b011101111100;
   12629: result <= 12'b011101111100;
   12630: result <= 12'b011101111100;
   12631: result <= 12'b011101111100;
   12632: result <= 12'b011101111100;
   12633: result <= 12'b011101111100;
   12634: result <= 12'b011101111101;
   12635: result <= 12'b011101111101;
   12636: result <= 12'b011101111101;
   12637: result <= 12'b011101111101;
   12638: result <= 12'b011101111101;
   12639: result <= 12'b011101111101;
   12640: result <= 12'b011101111101;
   12641: result <= 12'b011101111101;
   12642: result <= 12'b011101111101;
   12643: result <= 12'b011101111101;
   12644: result <= 12'b011101111101;
   12645: result <= 12'b011101111101;
   12646: result <= 12'b011101111101;
   12647: result <= 12'b011101111101;
   12648: result <= 12'b011101111110;
   12649: result <= 12'b011101111110;
   12650: result <= 12'b011101111110;
   12651: result <= 12'b011101111110;
   12652: result <= 12'b011101111110;
   12653: result <= 12'b011101111110;
   12654: result <= 12'b011101111110;
   12655: result <= 12'b011101111110;
   12656: result <= 12'b011101111110;
   12657: result <= 12'b011101111110;
   12658: result <= 12'b011101111110;
   12659: result <= 12'b011101111110;
   12660: result <= 12'b011101111110;
   12661: result <= 12'b011101111110;
   12662: result <= 12'b011101111110;
   12663: result <= 12'b011101111111;
   12664: result <= 12'b011101111111;
   12665: result <= 12'b011101111111;
   12666: result <= 12'b011101111111;
   12667: result <= 12'b011101111111;
   12668: result <= 12'b011101111111;
   12669: result <= 12'b011101111111;
   12670: result <= 12'b011101111111;
   12671: result <= 12'b011101111111;
   12672: result <= 12'b011101111111;
   12673: result <= 12'b011101111111;
   12674: result <= 12'b011101111111;
   12675: result <= 12'b011101111111;
   12676: result <= 12'b011101111111;
   12677: result <= 12'b011110000000;
   12678: result <= 12'b011110000000;
   12679: result <= 12'b011110000000;
   12680: result <= 12'b011110000000;
   12681: result <= 12'b011110000000;
   12682: result <= 12'b011110000000;
   12683: result <= 12'b011110000000;
   12684: result <= 12'b011110000000;
   12685: result <= 12'b011110000000;
   12686: result <= 12'b011110000000;
   12687: result <= 12'b011110000000;
   12688: result <= 12'b011110000000;
   12689: result <= 12'b011110000000;
   12690: result <= 12'b011110000000;
   12691: result <= 12'b011110000000;
   12692: result <= 12'b011110000001;
   12693: result <= 12'b011110000001;
   12694: result <= 12'b011110000001;
   12695: result <= 12'b011110000001;
   12696: result <= 12'b011110000001;
   12697: result <= 12'b011110000001;
   12698: result <= 12'b011110000001;
   12699: result <= 12'b011110000001;
   12700: result <= 12'b011110000001;
   12701: result <= 12'b011110000001;
   12702: result <= 12'b011110000001;
   12703: result <= 12'b011110000001;
   12704: result <= 12'b011110000001;
   12705: result <= 12'b011110000001;
   12706: result <= 12'b011110000001;
   12707: result <= 12'b011110000010;
   12708: result <= 12'b011110000010;
   12709: result <= 12'b011110000010;
   12710: result <= 12'b011110000010;
   12711: result <= 12'b011110000010;
   12712: result <= 12'b011110000010;
   12713: result <= 12'b011110000010;
   12714: result <= 12'b011110000010;
   12715: result <= 12'b011110000010;
   12716: result <= 12'b011110000010;
   12717: result <= 12'b011110000010;
   12718: result <= 12'b011110000010;
   12719: result <= 12'b011110000010;
   12720: result <= 12'b011110000010;
   12721: result <= 12'b011110000011;
   12722: result <= 12'b011110000011;
   12723: result <= 12'b011110000011;
   12724: result <= 12'b011110000011;
   12725: result <= 12'b011110000011;
   12726: result <= 12'b011110000011;
   12727: result <= 12'b011110000011;
   12728: result <= 12'b011110000011;
   12729: result <= 12'b011110000011;
   12730: result <= 12'b011110000011;
   12731: result <= 12'b011110000011;
   12732: result <= 12'b011110000011;
   12733: result <= 12'b011110000011;
   12734: result <= 12'b011110000011;
   12735: result <= 12'b011110000011;
   12736: result <= 12'b011110000100;
   12737: result <= 12'b011110000100;
   12738: result <= 12'b011110000100;
   12739: result <= 12'b011110000100;
   12740: result <= 12'b011110000100;
   12741: result <= 12'b011110000100;
   12742: result <= 12'b011110000100;
   12743: result <= 12'b011110000100;
   12744: result <= 12'b011110000100;
   12745: result <= 12'b011110000100;
   12746: result <= 12'b011110000100;
   12747: result <= 12'b011110000100;
   12748: result <= 12'b011110000100;
   12749: result <= 12'b011110000100;
   12750: result <= 12'b011110000100;
   12751: result <= 12'b011110000101;
   12752: result <= 12'b011110000101;
   12753: result <= 12'b011110000101;
   12754: result <= 12'b011110000101;
   12755: result <= 12'b011110000101;
   12756: result <= 12'b011110000101;
   12757: result <= 12'b011110000101;
   12758: result <= 12'b011110000101;
   12759: result <= 12'b011110000101;
   12760: result <= 12'b011110000101;
   12761: result <= 12'b011110000101;
   12762: result <= 12'b011110000101;
   12763: result <= 12'b011110000101;
   12764: result <= 12'b011110000101;
   12765: result <= 12'b011110000101;
   12766: result <= 12'b011110000110;
   12767: result <= 12'b011110000110;
   12768: result <= 12'b011110000110;
   12769: result <= 12'b011110000110;
   12770: result <= 12'b011110000110;
   12771: result <= 12'b011110000110;
   12772: result <= 12'b011110000110;
   12773: result <= 12'b011110000110;
   12774: result <= 12'b011110000110;
   12775: result <= 12'b011110000110;
   12776: result <= 12'b011110000110;
   12777: result <= 12'b011110000110;
   12778: result <= 12'b011110000110;
   12779: result <= 12'b011110000110;
   12780: result <= 12'b011110000110;
   12781: result <= 12'b011110000111;
   12782: result <= 12'b011110000111;
   12783: result <= 12'b011110000111;
   12784: result <= 12'b011110000111;
   12785: result <= 12'b011110000111;
   12786: result <= 12'b011110000111;
   12787: result <= 12'b011110000111;
   12788: result <= 12'b011110000111;
   12789: result <= 12'b011110000111;
   12790: result <= 12'b011110000111;
   12791: result <= 12'b011110000111;
   12792: result <= 12'b011110000111;
   12793: result <= 12'b011110000111;
   12794: result <= 12'b011110000111;
   12795: result <= 12'b011110000111;
   12796: result <= 12'b011110001000;
   12797: result <= 12'b011110001000;
   12798: result <= 12'b011110001000;
   12799: result <= 12'b011110001000;
   12800: result <= 12'b011110001000;
   12801: result <= 12'b011110001000;
   12802: result <= 12'b011110001000;
   12803: result <= 12'b011110001000;
   12804: result <= 12'b011110001000;
   12805: result <= 12'b011110001000;
   12806: result <= 12'b011110001000;
   12807: result <= 12'b011110001000;
   12808: result <= 12'b011110001000;
   12809: result <= 12'b011110001000;
   12810: result <= 12'b011110001000;
   12811: result <= 12'b011110001001;
   12812: result <= 12'b011110001001;
   12813: result <= 12'b011110001001;
   12814: result <= 12'b011110001001;
   12815: result <= 12'b011110001001;
   12816: result <= 12'b011110001001;
   12817: result <= 12'b011110001001;
   12818: result <= 12'b011110001001;
   12819: result <= 12'b011110001001;
   12820: result <= 12'b011110001001;
   12821: result <= 12'b011110001001;
   12822: result <= 12'b011110001001;
   12823: result <= 12'b011110001001;
   12824: result <= 12'b011110001001;
   12825: result <= 12'b011110001001;
   12826: result <= 12'b011110001001;
   12827: result <= 12'b011110001010;
   12828: result <= 12'b011110001010;
   12829: result <= 12'b011110001010;
   12830: result <= 12'b011110001010;
   12831: result <= 12'b011110001010;
   12832: result <= 12'b011110001010;
   12833: result <= 12'b011110001010;
   12834: result <= 12'b011110001010;
   12835: result <= 12'b011110001010;
   12836: result <= 12'b011110001010;
   12837: result <= 12'b011110001010;
   12838: result <= 12'b011110001010;
   12839: result <= 12'b011110001010;
   12840: result <= 12'b011110001010;
   12841: result <= 12'b011110001010;
   12842: result <= 12'b011110001011;
   12843: result <= 12'b011110001011;
   12844: result <= 12'b011110001011;
   12845: result <= 12'b011110001011;
   12846: result <= 12'b011110001011;
   12847: result <= 12'b011110001011;
   12848: result <= 12'b011110001011;
   12849: result <= 12'b011110001011;
   12850: result <= 12'b011110001011;
   12851: result <= 12'b011110001011;
   12852: result <= 12'b011110001011;
   12853: result <= 12'b011110001011;
   12854: result <= 12'b011110001011;
   12855: result <= 12'b011110001011;
   12856: result <= 12'b011110001011;
   12857: result <= 12'b011110001100;
   12858: result <= 12'b011110001100;
   12859: result <= 12'b011110001100;
   12860: result <= 12'b011110001100;
   12861: result <= 12'b011110001100;
   12862: result <= 12'b011110001100;
   12863: result <= 12'b011110001100;
   12864: result <= 12'b011110001100;
   12865: result <= 12'b011110001100;
   12866: result <= 12'b011110001100;
   12867: result <= 12'b011110001100;
   12868: result <= 12'b011110001100;
   12869: result <= 12'b011110001100;
   12870: result <= 12'b011110001100;
   12871: result <= 12'b011110001100;
   12872: result <= 12'b011110001100;
   12873: result <= 12'b011110001101;
   12874: result <= 12'b011110001101;
   12875: result <= 12'b011110001101;
   12876: result <= 12'b011110001101;
   12877: result <= 12'b011110001101;
   12878: result <= 12'b011110001101;
   12879: result <= 12'b011110001101;
   12880: result <= 12'b011110001101;
   12881: result <= 12'b011110001101;
   12882: result <= 12'b011110001101;
   12883: result <= 12'b011110001101;
   12884: result <= 12'b011110001101;
   12885: result <= 12'b011110001101;
   12886: result <= 12'b011110001101;
   12887: result <= 12'b011110001101;
   12888: result <= 12'b011110001110;
   12889: result <= 12'b011110001110;
   12890: result <= 12'b011110001110;
   12891: result <= 12'b011110001110;
   12892: result <= 12'b011110001110;
   12893: result <= 12'b011110001110;
   12894: result <= 12'b011110001110;
   12895: result <= 12'b011110001110;
   12896: result <= 12'b011110001110;
   12897: result <= 12'b011110001110;
   12898: result <= 12'b011110001110;
   12899: result <= 12'b011110001110;
   12900: result <= 12'b011110001110;
   12901: result <= 12'b011110001110;
   12902: result <= 12'b011110001110;
   12903: result <= 12'b011110001111;
   12904: result <= 12'b011110001111;
   12905: result <= 12'b011110001111;
   12906: result <= 12'b011110001111;
   12907: result <= 12'b011110001111;
   12908: result <= 12'b011110001111;
   12909: result <= 12'b011110001111;
   12910: result <= 12'b011110001111;
   12911: result <= 12'b011110001111;
   12912: result <= 12'b011110001111;
   12913: result <= 12'b011110001111;
   12914: result <= 12'b011110001111;
   12915: result <= 12'b011110001111;
   12916: result <= 12'b011110001111;
   12917: result <= 12'b011110001111;
   12918: result <= 12'b011110001111;
   12919: result <= 12'b011110010000;
   12920: result <= 12'b011110010000;
   12921: result <= 12'b011110010000;
   12922: result <= 12'b011110010000;
   12923: result <= 12'b011110010000;
   12924: result <= 12'b011110010000;
   12925: result <= 12'b011110010000;
   12926: result <= 12'b011110010000;
   12927: result <= 12'b011110010000;
   12928: result <= 12'b011110010000;
   12929: result <= 12'b011110010000;
   12930: result <= 12'b011110010000;
   12931: result <= 12'b011110010000;
   12932: result <= 12'b011110010000;
   12933: result <= 12'b011110010000;
   12934: result <= 12'b011110010000;
   12935: result <= 12'b011110010001;
   12936: result <= 12'b011110010001;
   12937: result <= 12'b011110010001;
   12938: result <= 12'b011110010001;
   12939: result <= 12'b011110010001;
   12940: result <= 12'b011110010001;
   12941: result <= 12'b011110010001;
   12942: result <= 12'b011110010001;
   12943: result <= 12'b011110010001;
   12944: result <= 12'b011110010001;
   12945: result <= 12'b011110010001;
   12946: result <= 12'b011110010001;
   12947: result <= 12'b011110010001;
   12948: result <= 12'b011110010001;
   12949: result <= 12'b011110010001;
   12950: result <= 12'b011110010010;
   12951: result <= 12'b011110010010;
   12952: result <= 12'b011110010010;
   12953: result <= 12'b011110010010;
   12954: result <= 12'b011110010010;
   12955: result <= 12'b011110010010;
   12956: result <= 12'b011110010010;
   12957: result <= 12'b011110010010;
   12958: result <= 12'b011110010010;
   12959: result <= 12'b011110010010;
   12960: result <= 12'b011110010010;
   12961: result <= 12'b011110010010;
   12962: result <= 12'b011110010010;
   12963: result <= 12'b011110010010;
   12964: result <= 12'b011110010010;
   12965: result <= 12'b011110010010;
   12966: result <= 12'b011110010011;
   12967: result <= 12'b011110010011;
   12968: result <= 12'b011110010011;
   12969: result <= 12'b011110010011;
   12970: result <= 12'b011110010011;
   12971: result <= 12'b011110010011;
   12972: result <= 12'b011110010011;
   12973: result <= 12'b011110010011;
   12974: result <= 12'b011110010011;
   12975: result <= 12'b011110010011;
   12976: result <= 12'b011110010011;
   12977: result <= 12'b011110010011;
   12978: result <= 12'b011110010011;
   12979: result <= 12'b011110010011;
   12980: result <= 12'b011110010011;
   12981: result <= 12'b011110010011;
   12982: result <= 12'b011110010100;
   12983: result <= 12'b011110010100;
   12984: result <= 12'b011110010100;
   12985: result <= 12'b011110010100;
   12986: result <= 12'b011110010100;
   12987: result <= 12'b011110010100;
   12988: result <= 12'b011110010100;
   12989: result <= 12'b011110010100;
   12990: result <= 12'b011110010100;
   12991: result <= 12'b011110010100;
   12992: result <= 12'b011110010100;
   12993: result <= 12'b011110010100;
   12994: result <= 12'b011110010100;
   12995: result <= 12'b011110010100;
   12996: result <= 12'b011110010100;
   12997: result <= 12'b011110010100;
   12998: result <= 12'b011110010101;
   12999: result <= 12'b011110010101;
   13000: result <= 12'b011110010101;
   13001: result <= 12'b011110010101;
   13002: result <= 12'b011110010101;
   13003: result <= 12'b011110010101;
   13004: result <= 12'b011110010101;
   13005: result <= 12'b011110010101;
   13006: result <= 12'b011110010101;
   13007: result <= 12'b011110010101;
   13008: result <= 12'b011110010101;
   13009: result <= 12'b011110010101;
   13010: result <= 12'b011110010101;
   13011: result <= 12'b011110010101;
   13012: result <= 12'b011110010101;
   13013: result <= 12'b011110010101;
   13014: result <= 12'b011110010110;
   13015: result <= 12'b011110010110;
   13016: result <= 12'b011110010110;
   13017: result <= 12'b011110010110;
   13018: result <= 12'b011110010110;
   13019: result <= 12'b011110010110;
   13020: result <= 12'b011110010110;
   13021: result <= 12'b011110010110;
   13022: result <= 12'b011110010110;
   13023: result <= 12'b011110010110;
   13024: result <= 12'b011110010110;
   13025: result <= 12'b011110010110;
   13026: result <= 12'b011110010110;
   13027: result <= 12'b011110010110;
   13028: result <= 12'b011110010110;
   13029: result <= 12'b011110010110;
   13030: result <= 12'b011110010111;
   13031: result <= 12'b011110010111;
   13032: result <= 12'b011110010111;
   13033: result <= 12'b011110010111;
   13034: result <= 12'b011110010111;
   13035: result <= 12'b011110010111;
   13036: result <= 12'b011110010111;
   13037: result <= 12'b011110010111;
   13038: result <= 12'b011110010111;
   13039: result <= 12'b011110010111;
   13040: result <= 12'b011110010111;
   13041: result <= 12'b011110010111;
   13042: result <= 12'b011110010111;
   13043: result <= 12'b011110010111;
   13044: result <= 12'b011110010111;
   13045: result <= 12'b011110010111;
   13046: result <= 12'b011110011000;
   13047: result <= 12'b011110011000;
   13048: result <= 12'b011110011000;
   13049: result <= 12'b011110011000;
   13050: result <= 12'b011110011000;
   13051: result <= 12'b011110011000;
   13052: result <= 12'b011110011000;
   13053: result <= 12'b011110011000;
   13054: result <= 12'b011110011000;
   13055: result <= 12'b011110011000;
   13056: result <= 12'b011110011000;
   13057: result <= 12'b011110011000;
   13058: result <= 12'b011110011000;
   13059: result <= 12'b011110011000;
   13060: result <= 12'b011110011000;
   13061: result <= 12'b011110011000;
   13062: result <= 12'b011110011001;
   13063: result <= 12'b011110011001;
   13064: result <= 12'b011110011001;
   13065: result <= 12'b011110011001;
   13066: result <= 12'b011110011001;
   13067: result <= 12'b011110011001;
   13068: result <= 12'b011110011001;
   13069: result <= 12'b011110011001;
   13070: result <= 12'b011110011001;
   13071: result <= 12'b011110011001;
   13072: result <= 12'b011110011001;
   13073: result <= 12'b011110011001;
   13074: result <= 12'b011110011001;
   13075: result <= 12'b011110011001;
   13076: result <= 12'b011110011001;
   13077: result <= 12'b011110011001;
   13078: result <= 12'b011110011001;
   13079: result <= 12'b011110011010;
   13080: result <= 12'b011110011010;
   13081: result <= 12'b011110011010;
   13082: result <= 12'b011110011010;
   13083: result <= 12'b011110011010;
   13084: result <= 12'b011110011010;
   13085: result <= 12'b011110011010;
   13086: result <= 12'b011110011010;
   13087: result <= 12'b011110011010;
   13088: result <= 12'b011110011010;
   13089: result <= 12'b011110011010;
   13090: result <= 12'b011110011010;
   13091: result <= 12'b011110011010;
   13092: result <= 12'b011110011010;
   13093: result <= 12'b011110011010;
   13094: result <= 12'b011110011010;
   13095: result <= 12'b011110011011;
   13096: result <= 12'b011110011011;
   13097: result <= 12'b011110011011;
   13098: result <= 12'b011110011011;
   13099: result <= 12'b011110011011;
   13100: result <= 12'b011110011011;
   13101: result <= 12'b011110011011;
   13102: result <= 12'b011110011011;
   13103: result <= 12'b011110011011;
   13104: result <= 12'b011110011011;
   13105: result <= 12'b011110011011;
   13106: result <= 12'b011110011011;
   13107: result <= 12'b011110011011;
   13108: result <= 12'b011110011011;
   13109: result <= 12'b011110011011;
   13110: result <= 12'b011110011011;
   13111: result <= 12'b011110011011;
   13112: result <= 12'b011110011100;
   13113: result <= 12'b011110011100;
   13114: result <= 12'b011110011100;
   13115: result <= 12'b011110011100;
   13116: result <= 12'b011110011100;
   13117: result <= 12'b011110011100;
   13118: result <= 12'b011110011100;
   13119: result <= 12'b011110011100;
   13120: result <= 12'b011110011100;
   13121: result <= 12'b011110011100;
   13122: result <= 12'b011110011100;
   13123: result <= 12'b011110011100;
   13124: result <= 12'b011110011100;
   13125: result <= 12'b011110011100;
   13126: result <= 12'b011110011100;
   13127: result <= 12'b011110011100;
   13128: result <= 12'b011110011101;
   13129: result <= 12'b011110011101;
   13130: result <= 12'b011110011101;
   13131: result <= 12'b011110011101;
   13132: result <= 12'b011110011101;
   13133: result <= 12'b011110011101;
   13134: result <= 12'b011110011101;
   13135: result <= 12'b011110011101;
   13136: result <= 12'b011110011101;
   13137: result <= 12'b011110011101;
   13138: result <= 12'b011110011101;
   13139: result <= 12'b011110011101;
   13140: result <= 12'b011110011101;
   13141: result <= 12'b011110011101;
   13142: result <= 12'b011110011101;
   13143: result <= 12'b011110011101;
   13144: result <= 12'b011110011101;
   13145: result <= 12'b011110011110;
   13146: result <= 12'b011110011110;
   13147: result <= 12'b011110011110;
   13148: result <= 12'b011110011110;
   13149: result <= 12'b011110011110;
   13150: result <= 12'b011110011110;
   13151: result <= 12'b011110011110;
   13152: result <= 12'b011110011110;
   13153: result <= 12'b011110011110;
   13154: result <= 12'b011110011110;
   13155: result <= 12'b011110011110;
   13156: result <= 12'b011110011110;
   13157: result <= 12'b011110011110;
   13158: result <= 12'b011110011110;
   13159: result <= 12'b011110011110;
   13160: result <= 12'b011110011110;
   13161: result <= 12'b011110011111;
   13162: result <= 12'b011110011111;
   13163: result <= 12'b011110011111;
   13164: result <= 12'b011110011111;
   13165: result <= 12'b011110011111;
   13166: result <= 12'b011110011111;
   13167: result <= 12'b011110011111;
   13168: result <= 12'b011110011111;
   13169: result <= 12'b011110011111;
   13170: result <= 12'b011110011111;
   13171: result <= 12'b011110011111;
   13172: result <= 12'b011110011111;
   13173: result <= 12'b011110011111;
   13174: result <= 12'b011110011111;
   13175: result <= 12'b011110011111;
   13176: result <= 12'b011110011111;
   13177: result <= 12'b011110011111;
   13178: result <= 12'b011110100000;
   13179: result <= 12'b011110100000;
   13180: result <= 12'b011110100000;
   13181: result <= 12'b011110100000;
   13182: result <= 12'b011110100000;
   13183: result <= 12'b011110100000;
   13184: result <= 12'b011110100000;
   13185: result <= 12'b011110100000;
   13186: result <= 12'b011110100000;
   13187: result <= 12'b011110100000;
   13188: result <= 12'b011110100000;
   13189: result <= 12'b011110100000;
   13190: result <= 12'b011110100000;
   13191: result <= 12'b011110100000;
   13192: result <= 12'b011110100000;
   13193: result <= 12'b011110100000;
   13194: result <= 12'b011110100000;
   13195: result <= 12'b011110100001;
   13196: result <= 12'b011110100001;
   13197: result <= 12'b011110100001;
   13198: result <= 12'b011110100001;
   13199: result <= 12'b011110100001;
   13200: result <= 12'b011110100001;
   13201: result <= 12'b011110100001;
   13202: result <= 12'b011110100001;
   13203: result <= 12'b011110100001;
   13204: result <= 12'b011110100001;
   13205: result <= 12'b011110100001;
   13206: result <= 12'b011110100001;
   13207: result <= 12'b011110100001;
   13208: result <= 12'b011110100001;
   13209: result <= 12'b011110100001;
   13210: result <= 12'b011110100001;
   13211: result <= 12'b011110100001;
   13212: result <= 12'b011110100010;
   13213: result <= 12'b011110100010;
   13214: result <= 12'b011110100010;
   13215: result <= 12'b011110100010;
   13216: result <= 12'b011110100010;
   13217: result <= 12'b011110100010;
   13218: result <= 12'b011110100010;
   13219: result <= 12'b011110100010;
   13220: result <= 12'b011110100010;
   13221: result <= 12'b011110100010;
   13222: result <= 12'b011110100010;
   13223: result <= 12'b011110100010;
   13224: result <= 12'b011110100010;
   13225: result <= 12'b011110100010;
   13226: result <= 12'b011110100010;
   13227: result <= 12'b011110100010;
   13228: result <= 12'b011110100010;
   13229: result <= 12'b011110100011;
   13230: result <= 12'b011110100011;
   13231: result <= 12'b011110100011;
   13232: result <= 12'b011110100011;
   13233: result <= 12'b011110100011;
   13234: result <= 12'b011110100011;
   13235: result <= 12'b011110100011;
   13236: result <= 12'b011110100011;
   13237: result <= 12'b011110100011;
   13238: result <= 12'b011110100011;
   13239: result <= 12'b011110100011;
   13240: result <= 12'b011110100011;
   13241: result <= 12'b011110100011;
   13242: result <= 12'b011110100011;
   13243: result <= 12'b011110100011;
   13244: result <= 12'b011110100011;
   13245: result <= 12'b011110100011;
   13246: result <= 12'b011110100100;
   13247: result <= 12'b011110100100;
   13248: result <= 12'b011110100100;
   13249: result <= 12'b011110100100;
   13250: result <= 12'b011110100100;
   13251: result <= 12'b011110100100;
   13252: result <= 12'b011110100100;
   13253: result <= 12'b011110100100;
   13254: result <= 12'b011110100100;
   13255: result <= 12'b011110100100;
   13256: result <= 12'b011110100100;
   13257: result <= 12'b011110100100;
   13258: result <= 12'b011110100100;
   13259: result <= 12'b011110100100;
   13260: result <= 12'b011110100100;
   13261: result <= 12'b011110100100;
   13262: result <= 12'b011110100100;
   13263: result <= 12'b011110100100;
   13264: result <= 12'b011110100101;
   13265: result <= 12'b011110100101;
   13266: result <= 12'b011110100101;
   13267: result <= 12'b011110100101;
   13268: result <= 12'b011110100101;
   13269: result <= 12'b011110100101;
   13270: result <= 12'b011110100101;
   13271: result <= 12'b011110100101;
   13272: result <= 12'b011110100101;
   13273: result <= 12'b011110100101;
   13274: result <= 12'b011110100101;
   13275: result <= 12'b011110100101;
   13276: result <= 12'b011110100101;
   13277: result <= 12'b011110100101;
   13278: result <= 12'b011110100101;
   13279: result <= 12'b011110100101;
   13280: result <= 12'b011110100101;
   13281: result <= 12'b011110100110;
   13282: result <= 12'b011110100110;
   13283: result <= 12'b011110100110;
   13284: result <= 12'b011110100110;
   13285: result <= 12'b011110100110;
   13286: result <= 12'b011110100110;
   13287: result <= 12'b011110100110;
   13288: result <= 12'b011110100110;
   13289: result <= 12'b011110100110;
   13290: result <= 12'b011110100110;
   13291: result <= 12'b011110100110;
   13292: result <= 12'b011110100110;
   13293: result <= 12'b011110100110;
   13294: result <= 12'b011110100110;
   13295: result <= 12'b011110100110;
   13296: result <= 12'b011110100110;
   13297: result <= 12'b011110100110;
   13298: result <= 12'b011110100111;
   13299: result <= 12'b011110100111;
   13300: result <= 12'b011110100111;
   13301: result <= 12'b011110100111;
   13302: result <= 12'b011110100111;
   13303: result <= 12'b011110100111;
   13304: result <= 12'b011110100111;
   13305: result <= 12'b011110100111;
   13306: result <= 12'b011110100111;
   13307: result <= 12'b011110100111;
   13308: result <= 12'b011110100111;
   13309: result <= 12'b011110100111;
   13310: result <= 12'b011110100111;
   13311: result <= 12'b011110100111;
   13312: result <= 12'b011110100111;
   13313: result <= 12'b011110100111;
   13314: result <= 12'b011110100111;
   13315: result <= 12'b011110100111;
   13316: result <= 12'b011110101000;
   13317: result <= 12'b011110101000;
   13318: result <= 12'b011110101000;
   13319: result <= 12'b011110101000;
   13320: result <= 12'b011110101000;
   13321: result <= 12'b011110101000;
   13322: result <= 12'b011110101000;
   13323: result <= 12'b011110101000;
   13324: result <= 12'b011110101000;
   13325: result <= 12'b011110101000;
   13326: result <= 12'b011110101000;
   13327: result <= 12'b011110101000;
   13328: result <= 12'b011110101000;
   13329: result <= 12'b011110101000;
   13330: result <= 12'b011110101000;
   13331: result <= 12'b011110101000;
   13332: result <= 12'b011110101000;
   13333: result <= 12'b011110101001;
   13334: result <= 12'b011110101001;
   13335: result <= 12'b011110101001;
   13336: result <= 12'b011110101001;
   13337: result <= 12'b011110101001;
   13338: result <= 12'b011110101001;
   13339: result <= 12'b011110101001;
   13340: result <= 12'b011110101001;
   13341: result <= 12'b011110101001;
   13342: result <= 12'b011110101001;
   13343: result <= 12'b011110101001;
   13344: result <= 12'b011110101001;
   13345: result <= 12'b011110101001;
   13346: result <= 12'b011110101001;
   13347: result <= 12'b011110101001;
   13348: result <= 12'b011110101001;
   13349: result <= 12'b011110101001;
   13350: result <= 12'b011110101001;
   13351: result <= 12'b011110101010;
   13352: result <= 12'b011110101010;
   13353: result <= 12'b011110101010;
   13354: result <= 12'b011110101010;
   13355: result <= 12'b011110101010;
   13356: result <= 12'b011110101010;
   13357: result <= 12'b011110101010;
   13358: result <= 12'b011110101010;
   13359: result <= 12'b011110101010;
   13360: result <= 12'b011110101010;
   13361: result <= 12'b011110101010;
   13362: result <= 12'b011110101010;
   13363: result <= 12'b011110101010;
   13364: result <= 12'b011110101010;
   13365: result <= 12'b011110101010;
   13366: result <= 12'b011110101010;
   13367: result <= 12'b011110101010;
   13368: result <= 12'b011110101010;
   13369: result <= 12'b011110101011;
   13370: result <= 12'b011110101011;
   13371: result <= 12'b011110101011;
   13372: result <= 12'b011110101011;
   13373: result <= 12'b011110101011;
   13374: result <= 12'b011110101011;
   13375: result <= 12'b011110101011;
   13376: result <= 12'b011110101011;
   13377: result <= 12'b011110101011;
   13378: result <= 12'b011110101011;
   13379: result <= 12'b011110101011;
   13380: result <= 12'b011110101011;
   13381: result <= 12'b011110101011;
   13382: result <= 12'b011110101011;
   13383: result <= 12'b011110101011;
   13384: result <= 12'b011110101011;
   13385: result <= 12'b011110101011;
   13386: result <= 12'b011110101011;
   13387: result <= 12'b011110101100;
   13388: result <= 12'b011110101100;
   13389: result <= 12'b011110101100;
   13390: result <= 12'b011110101100;
   13391: result <= 12'b011110101100;
   13392: result <= 12'b011110101100;
   13393: result <= 12'b011110101100;
   13394: result <= 12'b011110101100;
   13395: result <= 12'b011110101100;
   13396: result <= 12'b011110101100;
   13397: result <= 12'b011110101100;
   13398: result <= 12'b011110101100;
   13399: result <= 12'b011110101100;
   13400: result <= 12'b011110101100;
   13401: result <= 12'b011110101100;
   13402: result <= 12'b011110101100;
   13403: result <= 12'b011110101100;
   13404: result <= 12'b011110101100;
   13405: result <= 12'b011110101101;
   13406: result <= 12'b011110101101;
   13407: result <= 12'b011110101101;
   13408: result <= 12'b011110101101;
   13409: result <= 12'b011110101101;
   13410: result <= 12'b011110101101;
   13411: result <= 12'b011110101101;
   13412: result <= 12'b011110101101;
   13413: result <= 12'b011110101101;
   13414: result <= 12'b011110101101;
   13415: result <= 12'b011110101101;
   13416: result <= 12'b011110101101;
   13417: result <= 12'b011110101101;
   13418: result <= 12'b011110101101;
   13419: result <= 12'b011110101101;
   13420: result <= 12'b011110101101;
   13421: result <= 12'b011110101101;
   13422: result <= 12'b011110101101;
   13423: result <= 12'b011110101110;
   13424: result <= 12'b011110101110;
   13425: result <= 12'b011110101110;
   13426: result <= 12'b011110101110;
   13427: result <= 12'b011110101110;
   13428: result <= 12'b011110101110;
   13429: result <= 12'b011110101110;
   13430: result <= 12'b011110101110;
   13431: result <= 12'b011110101110;
   13432: result <= 12'b011110101110;
   13433: result <= 12'b011110101110;
   13434: result <= 12'b011110101110;
   13435: result <= 12'b011110101110;
   13436: result <= 12'b011110101110;
   13437: result <= 12'b011110101110;
   13438: result <= 12'b011110101110;
   13439: result <= 12'b011110101110;
   13440: result <= 12'b011110101110;
   13441: result <= 12'b011110101111;
   13442: result <= 12'b011110101111;
   13443: result <= 12'b011110101111;
   13444: result <= 12'b011110101111;
   13445: result <= 12'b011110101111;
   13446: result <= 12'b011110101111;
   13447: result <= 12'b011110101111;
   13448: result <= 12'b011110101111;
   13449: result <= 12'b011110101111;
   13450: result <= 12'b011110101111;
   13451: result <= 12'b011110101111;
   13452: result <= 12'b011110101111;
   13453: result <= 12'b011110101111;
   13454: result <= 12'b011110101111;
   13455: result <= 12'b011110101111;
   13456: result <= 12'b011110101111;
   13457: result <= 12'b011110101111;
   13458: result <= 12'b011110101111;
   13459: result <= 12'b011110101111;
   13460: result <= 12'b011110110000;
   13461: result <= 12'b011110110000;
   13462: result <= 12'b011110110000;
   13463: result <= 12'b011110110000;
   13464: result <= 12'b011110110000;
   13465: result <= 12'b011110110000;
   13466: result <= 12'b011110110000;
   13467: result <= 12'b011110110000;
   13468: result <= 12'b011110110000;
   13469: result <= 12'b011110110000;
   13470: result <= 12'b011110110000;
   13471: result <= 12'b011110110000;
   13472: result <= 12'b011110110000;
   13473: result <= 12'b011110110000;
   13474: result <= 12'b011110110000;
   13475: result <= 12'b011110110000;
   13476: result <= 12'b011110110000;
   13477: result <= 12'b011110110000;
   13478: result <= 12'b011110110001;
   13479: result <= 12'b011110110001;
   13480: result <= 12'b011110110001;
   13481: result <= 12'b011110110001;
   13482: result <= 12'b011110110001;
   13483: result <= 12'b011110110001;
   13484: result <= 12'b011110110001;
   13485: result <= 12'b011110110001;
   13486: result <= 12'b011110110001;
   13487: result <= 12'b011110110001;
   13488: result <= 12'b011110110001;
   13489: result <= 12'b011110110001;
   13490: result <= 12'b011110110001;
   13491: result <= 12'b011110110001;
   13492: result <= 12'b011110110001;
   13493: result <= 12'b011110110001;
   13494: result <= 12'b011110110001;
   13495: result <= 12'b011110110001;
   13496: result <= 12'b011110110001;
   13497: result <= 12'b011110110010;
   13498: result <= 12'b011110110010;
   13499: result <= 12'b011110110010;
   13500: result <= 12'b011110110010;
   13501: result <= 12'b011110110010;
   13502: result <= 12'b011110110010;
   13503: result <= 12'b011110110010;
   13504: result <= 12'b011110110010;
   13505: result <= 12'b011110110010;
   13506: result <= 12'b011110110010;
   13507: result <= 12'b011110110010;
   13508: result <= 12'b011110110010;
   13509: result <= 12'b011110110010;
   13510: result <= 12'b011110110010;
   13511: result <= 12'b011110110010;
   13512: result <= 12'b011110110010;
   13513: result <= 12'b011110110010;
   13514: result <= 12'b011110110010;
   13515: result <= 12'b011110110011;
   13516: result <= 12'b011110110011;
   13517: result <= 12'b011110110011;
   13518: result <= 12'b011110110011;
   13519: result <= 12'b011110110011;
   13520: result <= 12'b011110110011;
   13521: result <= 12'b011110110011;
   13522: result <= 12'b011110110011;
   13523: result <= 12'b011110110011;
   13524: result <= 12'b011110110011;
   13525: result <= 12'b011110110011;
   13526: result <= 12'b011110110011;
   13527: result <= 12'b011110110011;
   13528: result <= 12'b011110110011;
   13529: result <= 12'b011110110011;
   13530: result <= 12'b011110110011;
   13531: result <= 12'b011110110011;
   13532: result <= 12'b011110110011;
   13533: result <= 12'b011110110011;
   13534: result <= 12'b011110110100;
   13535: result <= 12'b011110110100;
   13536: result <= 12'b011110110100;
   13537: result <= 12'b011110110100;
   13538: result <= 12'b011110110100;
   13539: result <= 12'b011110110100;
   13540: result <= 12'b011110110100;
   13541: result <= 12'b011110110100;
   13542: result <= 12'b011110110100;
   13543: result <= 12'b011110110100;
   13544: result <= 12'b011110110100;
   13545: result <= 12'b011110110100;
   13546: result <= 12'b011110110100;
   13547: result <= 12'b011110110100;
   13548: result <= 12'b011110110100;
   13549: result <= 12'b011110110100;
   13550: result <= 12'b011110110100;
   13551: result <= 12'b011110110100;
   13552: result <= 12'b011110110100;
   13553: result <= 12'b011110110101;
   13554: result <= 12'b011110110101;
   13555: result <= 12'b011110110101;
   13556: result <= 12'b011110110101;
   13557: result <= 12'b011110110101;
   13558: result <= 12'b011110110101;
   13559: result <= 12'b011110110101;
   13560: result <= 12'b011110110101;
   13561: result <= 12'b011110110101;
   13562: result <= 12'b011110110101;
   13563: result <= 12'b011110110101;
   13564: result <= 12'b011110110101;
   13565: result <= 12'b011110110101;
   13566: result <= 12'b011110110101;
   13567: result <= 12'b011110110101;
   13568: result <= 12'b011110110101;
   13569: result <= 12'b011110110101;
   13570: result <= 12'b011110110101;
   13571: result <= 12'b011110110101;
   13572: result <= 12'b011110110110;
   13573: result <= 12'b011110110110;
   13574: result <= 12'b011110110110;
   13575: result <= 12'b011110110110;
   13576: result <= 12'b011110110110;
   13577: result <= 12'b011110110110;
   13578: result <= 12'b011110110110;
   13579: result <= 12'b011110110110;
   13580: result <= 12'b011110110110;
   13581: result <= 12'b011110110110;
   13582: result <= 12'b011110110110;
   13583: result <= 12'b011110110110;
   13584: result <= 12'b011110110110;
   13585: result <= 12'b011110110110;
   13586: result <= 12'b011110110110;
   13587: result <= 12'b011110110110;
   13588: result <= 12'b011110110110;
   13589: result <= 12'b011110110110;
   13590: result <= 12'b011110110110;
   13591: result <= 12'b011110110111;
   13592: result <= 12'b011110110111;
   13593: result <= 12'b011110110111;
   13594: result <= 12'b011110110111;
   13595: result <= 12'b011110110111;
   13596: result <= 12'b011110110111;
   13597: result <= 12'b011110110111;
   13598: result <= 12'b011110110111;
   13599: result <= 12'b011110110111;
   13600: result <= 12'b011110110111;
   13601: result <= 12'b011110110111;
   13602: result <= 12'b011110110111;
   13603: result <= 12'b011110110111;
   13604: result <= 12'b011110110111;
   13605: result <= 12'b011110110111;
   13606: result <= 12'b011110110111;
   13607: result <= 12'b011110110111;
   13608: result <= 12'b011110110111;
   13609: result <= 12'b011110110111;
   13610: result <= 12'b011110110111;
   13611: result <= 12'b011110111000;
   13612: result <= 12'b011110111000;
   13613: result <= 12'b011110111000;
   13614: result <= 12'b011110111000;
   13615: result <= 12'b011110111000;
   13616: result <= 12'b011110111000;
   13617: result <= 12'b011110111000;
   13618: result <= 12'b011110111000;
   13619: result <= 12'b011110111000;
   13620: result <= 12'b011110111000;
   13621: result <= 12'b011110111000;
   13622: result <= 12'b011110111000;
   13623: result <= 12'b011110111000;
   13624: result <= 12'b011110111000;
   13625: result <= 12'b011110111000;
   13626: result <= 12'b011110111000;
   13627: result <= 12'b011110111000;
   13628: result <= 12'b011110111000;
   13629: result <= 12'b011110111000;
   13630: result <= 12'b011110111001;
   13631: result <= 12'b011110111001;
   13632: result <= 12'b011110111001;
   13633: result <= 12'b011110111001;
   13634: result <= 12'b011110111001;
   13635: result <= 12'b011110111001;
   13636: result <= 12'b011110111001;
   13637: result <= 12'b011110111001;
   13638: result <= 12'b011110111001;
   13639: result <= 12'b011110111001;
   13640: result <= 12'b011110111001;
   13641: result <= 12'b011110111001;
   13642: result <= 12'b011110111001;
   13643: result <= 12'b011110111001;
   13644: result <= 12'b011110111001;
   13645: result <= 12'b011110111001;
   13646: result <= 12'b011110111001;
   13647: result <= 12'b011110111001;
   13648: result <= 12'b011110111001;
   13649: result <= 12'b011110111001;
   13650: result <= 12'b011110111010;
   13651: result <= 12'b011110111010;
   13652: result <= 12'b011110111010;
   13653: result <= 12'b011110111010;
   13654: result <= 12'b011110111010;
   13655: result <= 12'b011110111010;
   13656: result <= 12'b011110111010;
   13657: result <= 12'b011110111010;
   13658: result <= 12'b011110111010;
   13659: result <= 12'b011110111010;
   13660: result <= 12'b011110111010;
   13661: result <= 12'b011110111010;
   13662: result <= 12'b011110111010;
   13663: result <= 12'b011110111010;
   13664: result <= 12'b011110111010;
   13665: result <= 12'b011110111010;
   13666: result <= 12'b011110111010;
   13667: result <= 12'b011110111010;
   13668: result <= 12'b011110111010;
   13669: result <= 12'b011110111011;
   13670: result <= 12'b011110111011;
   13671: result <= 12'b011110111011;
   13672: result <= 12'b011110111011;
   13673: result <= 12'b011110111011;
   13674: result <= 12'b011110111011;
   13675: result <= 12'b011110111011;
   13676: result <= 12'b011110111011;
   13677: result <= 12'b011110111011;
   13678: result <= 12'b011110111011;
   13679: result <= 12'b011110111011;
   13680: result <= 12'b011110111011;
   13681: result <= 12'b011110111011;
   13682: result <= 12'b011110111011;
   13683: result <= 12'b011110111011;
   13684: result <= 12'b011110111011;
   13685: result <= 12'b011110111011;
   13686: result <= 12'b011110111011;
   13687: result <= 12'b011110111011;
   13688: result <= 12'b011110111011;
   13689: result <= 12'b011110111100;
   13690: result <= 12'b011110111100;
   13691: result <= 12'b011110111100;
   13692: result <= 12'b011110111100;
   13693: result <= 12'b011110111100;
   13694: result <= 12'b011110111100;
   13695: result <= 12'b011110111100;
   13696: result <= 12'b011110111100;
   13697: result <= 12'b011110111100;
   13698: result <= 12'b011110111100;
   13699: result <= 12'b011110111100;
   13700: result <= 12'b011110111100;
   13701: result <= 12'b011110111100;
   13702: result <= 12'b011110111100;
   13703: result <= 12'b011110111100;
   13704: result <= 12'b011110111100;
   13705: result <= 12'b011110111100;
   13706: result <= 12'b011110111100;
   13707: result <= 12'b011110111100;
   13708: result <= 12'b011110111100;
   13709: result <= 12'b011110111101;
   13710: result <= 12'b011110111101;
   13711: result <= 12'b011110111101;
   13712: result <= 12'b011110111101;
   13713: result <= 12'b011110111101;
   13714: result <= 12'b011110111101;
   13715: result <= 12'b011110111101;
   13716: result <= 12'b011110111101;
   13717: result <= 12'b011110111101;
   13718: result <= 12'b011110111101;
   13719: result <= 12'b011110111101;
   13720: result <= 12'b011110111101;
   13721: result <= 12'b011110111101;
   13722: result <= 12'b011110111101;
   13723: result <= 12'b011110111101;
   13724: result <= 12'b011110111101;
   13725: result <= 12'b011110111101;
   13726: result <= 12'b011110111101;
   13727: result <= 12'b011110111101;
   13728: result <= 12'b011110111101;
   13729: result <= 12'b011110111110;
   13730: result <= 12'b011110111110;
   13731: result <= 12'b011110111110;
   13732: result <= 12'b011110111110;
   13733: result <= 12'b011110111110;
   13734: result <= 12'b011110111110;
   13735: result <= 12'b011110111110;
   13736: result <= 12'b011110111110;
   13737: result <= 12'b011110111110;
   13738: result <= 12'b011110111110;
   13739: result <= 12'b011110111110;
   13740: result <= 12'b011110111110;
   13741: result <= 12'b011110111110;
   13742: result <= 12'b011110111110;
   13743: result <= 12'b011110111110;
   13744: result <= 12'b011110111110;
   13745: result <= 12'b011110111110;
   13746: result <= 12'b011110111110;
   13747: result <= 12'b011110111110;
   13748: result <= 12'b011110111110;
   13749: result <= 12'b011110111110;
   13750: result <= 12'b011110111111;
   13751: result <= 12'b011110111111;
   13752: result <= 12'b011110111111;
   13753: result <= 12'b011110111111;
   13754: result <= 12'b011110111111;
   13755: result <= 12'b011110111111;
   13756: result <= 12'b011110111111;
   13757: result <= 12'b011110111111;
   13758: result <= 12'b011110111111;
   13759: result <= 12'b011110111111;
   13760: result <= 12'b011110111111;
   13761: result <= 12'b011110111111;
   13762: result <= 12'b011110111111;
   13763: result <= 12'b011110111111;
   13764: result <= 12'b011110111111;
   13765: result <= 12'b011110111111;
   13766: result <= 12'b011110111111;
   13767: result <= 12'b011110111111;
   13768: result <= 12'b011110111111;
   13769: result <= 12'b011110111111;
   13770: result <= 12'b011111000000;
   13771: result <= 12'b011111000000;
   13772: result <= 12'b011111000000;
   13773: result <= 12'b011111000000;
   13774: result <= 12'b011111000000;
   13775: result <= 12'b011111000000;
   13776: result <= 12'b011111000000;
   13777: result <= 12'b011111000000;
   13778: result <= 12'b011111000000;
   13779: result <= 12'b011111000000;
   13780: result <= 12'b011111000000;
   13781: result <= 12'b011111000000;
   13782: result <= 12'b011111000000;
   13783: result <= 12'b011111000000;
   13784: result <= 12'b011111000000;
   13785: result <= 12'b011111000000;
   13786: result <= 12'b011111000000;
   13787: result <= 12'b011111000000;
   13788: result <= 12'b011111000000;
   13789: result <= 12'b011111000000;
   13790: result <= 12'b011111000000;
   13791: result <= 12'b011111000001;
   13792: result <= 12'b011111000001;
   13793: result <= 12'b011111000001;
   13794: result <= 12'b011111000001;
   13795: result <= 12'b011111000001;
   13796: result <= 12'b011111000001;
   13797: result <= 12'b011111000001;
   13798: result <= 12'b011111000001;
   13799: result <= 12'b011111000001;
   13800: result <= 12'b011111000001;
   13801: result <= 12'b011111000001;
   13802: result <= 12'b011111000001;
   13803: result <= 12'b011111000001;
   13804: result <= 12'b011111000001;
   13805: result <= 12'b011111000001;
   13806: result <= 12'b011111000001;
   13807: result <= 12'b011111000001;
   13808: result <= 12'b011111000001;
   13809: result <= 12'b011111000001;
   13810: result <= 12'b011111000001;
   13811: result <= 12'b011111000010;
   13812: result <= 12'b011111000010;
   13813: result <= 12'b011111000010;
   13814: result <= 12'b011111000010;
   13815: result <= 12'b011111000010;
   13816: result <= 12'b011111000010;
   13817: result <= 12'b011111000010;
   13818: result <= 12'b011111000010;
   13819: result <= 12'b011111000010;
   13820: result <= 12'b011111000010;
   13821: result <= 12'b011111000010;
   13822: result <= 12'b011111000010;
   13823: result <= 12'b011111000010;
   13824: result <= 12'b011111000010;
   13825: result <= 12'b011111000010;
   13826: result <= 12'b011111000010;
   13827: result <= 12'b011111000010;
   13828: result <= 12'b011111000010;
   13829: result <= 12'b011111000010;
   13830: result <= 12'b011111000010;
   13831: result <= 12'b011111000010;
   13832: result <= 12'b011111000011;
   13833: result <= 12'b011111000011;
   13834: result <= 12'b011111000011;
   13835: result <= 12'b011111000011;
   13836: result <= 12'b011111000011;
   13837: result <= 12'b011111000011;
   13838: result <= 12'b011111000011;
   13839: result <= 12'b011111000011;
   13840: result <= 12'b011111000011;
   13841: result <= 12'b011111000011;
   13842: result <= 12'b011111000011;
   13843: result <= 12'b011111000011;
   13844: result <= 12'b011111000011;
   13845: result <= 12'b011111000011;
   13846: result <= 12'b011111000011;
   13847: result <= 12'b011111000011;
   13848: result <= 12'b011111000011;
   13849: result <= 12'b011111000011;
   13850: result <= 12'b011111000011;
   13851: result <= 12'b011111000011;
   13852: result <= 12'b011111000011;
   13853: result <= 12'b011111000011;
   13854: result <= 12'b011111000100;
   13855: result <= 12'b011111000100;
   13856: result <= 12'b011111000100;
   13857: result <= 12'b011111000100;
   13858: result <= 12'b011111000100;
   13859: result <= 12'b011111000100;
   13860: result <= 12'b011111000100;
   13861: result <= 12'b011111000100;
   13862: result <= 12'b011111000100;
   13863: result <= 12'b011111000100;
   13864: result <= 12'b011111000100;
   13865: result <= 12'b011111000100;
   13866: result <= 12'b011111000100;
   13867: result <= 12'b011111000100;
   13868: result <= 12'b011111000100;
   13869: result <= 12'b011111000100;
   13870: result <= 12'b011111000100;
   13871: result <= 12'b011111000100;
   13872: result <= 12'b011111000100;
   13873: result <= 12'b011111000100;
   13874: result <= 12'b011111000100;
   13875: result <= 12'b011111000101;
   13876: result <= 12'b011111000101;
   13877: result <= 12'b011111000101;
   13878: result <= 12'b011111000101;
   13879: result <= 12'b011111000101;
   13880: result <= 12'b011111000101;
   13881: result <= 12'b011111000101;
   13882: result <= 12'b011111000101;
   13883: result <= 12'b011111000101;
   13884: result <= 12'b011111000101;
   13885: result <= 12'b011111000101;
   13886: result <= 12'b011111000101;
   13887: result <= 12'b011111000101;
   13888: result <= 12'b011111000101;
   13889: result <= 12'b011111000101;
   13890: result <= 12'b011111000101;
   13891: result <= 12'b011111000101;
   13892: result <= 12'b011111000101;
   13893: result <= 12'b011111000101;
   13894: result <= 12'b011111000101;
   13895: result <= 12'b011111000101;
   13896: result <= 12'b011111000110;
   13897: result <= 12'b011111000110;
   13898: result <= 12'b011111000110;
   13899: result <= 12'b011111000110;
   13900: result <= 12'b011111000110;
   13901: result <= 12'b011111000110;
   13902: result <= 12'b011111000110;
   13903: result <= 12'b011111000110;
   13904: result <= 12'b011111000110;
   13905: result <= 12'b011111000110;
   13906: result <= 12'b011111000110;
   13907: result <= 12'b011111000110;
   13908: result <= 12'b011111000110;
   13909: result <= 12'b011111000110;
   13910: result <= 12'b011111000110;
   13911: result <= 12'b011111000110;
   13912: result <= 12'b011111000110;
   13913: result <= 12'b011111000110;
   13914: result <= 12'b011111000110;
   13915: result <= 12'b011111000110;
   13916: result <= 12'b011111000110;
   13917: result <= 12'b011111000110;
   13918: result <= 12'b011111000111;
   13919: result <= 12'b011111000111;
   13920: result <= 12'b011111000111;
   13921: result <= 12'b011111000111;
   13922: result <= 12'b011111000111;
   13923: result <= 12'b011111000111;
   13924: result <= 12'b011111000111;
   13925: result <= 12'b011111000111;
   13926: result <= 12'b011111000111;
   13927: result <= 12'b011111000111;
   13928: result <= 12'b011111000111;
   13929: result <= 12'b011111000111;
   13930: result <= 12'b011111000111;
   13931: result <= 12'b011111000111;
   13932: result <= 12'b011111000111;
   13933: result <= 12'b011111000111;
   13934: result <= 12'b011111000111;
   13935: result <= 12'b011111000111;
   13936: result <= 12'b011111000111;
   13937: result <= 12'b011111000111;
   13938: result <= 12'b011111000111;
   13939: result <= 12'b011111000111;
   13940: result <= 12'b011111001000;
   13941: result <= 12'b011111001000;
   13942: result <= 12'b011111001000;
   13943: result <= 12'b011111001000;
   13944: result <= 12'b011111001000;
   13945: result <= 12'b011111001000;
   13946: result <= 12'b011111001000;
   13947: result <= 12'b011111001000;
   13948: result <= 12'b011111001000;
   13949: result <= 12'b011111001000;
   13950: result <= 12'b011111001000;
   13951: result <= 12'b011111001000;
   13952: result <= 12'b011111001000;
   13953: result <= 12'b011111001000;
   13954: result <= 12'b011111001000;
   13955: result <= 12'b011111001000;
   13956: result <= 12'b011111001000;
   13957: result <= 12'b011111001000;
   13958: result <= 12'b011111001000;
   13959: result <= 12'b011111001000;
   13960: result <= 12'b011111001000;
   13961: result <= 12'b011111001000;
   13962: result <= 12'b011111001001;
   13963: result <= 12'b011111001001;
   13964: result <= 12'b011111001001;
   13965: result <= 12'b011111001001;
   13966: result <= 12'b011111001001;
   13967: result <= 12'b011111001001;
   13968: result <= 12'b011111001001;
   13969: result <= 12'b011111001001;
   13970: result <= 12'b011111001001;
   13971: result <= 12'b011111001001;
   13972: result <= 12'b011111001001;
   13973: result <= 12'b011111001001;
   13974: result <= 12'b011111001001;
   13975: result <= 12'b011111001001;
   13976: result <= 12'b011111001001;
   13977: result <= 12'b011111001001;
   13978: result <= 12'b011111001001;
   13979: result <= 12'b011111001001;
   13980: result <= 12'b011111001001;
   13981: result <= 12'b011111001001;
   13982: result <= 12'b011111001001;
   13983: result <= 12'b011111001001;
   13984: result <= 12'b011111001010;
   13985: result <= 12'b011111001010;
   13986: result <= 12'b011111001010;
   13987: result <= 12'b011111001010;
   13988: result <= 12'b011111001010;
   13989: result <= 12'b011111001010;
   13990: result <= 12'b011111001010;
   13991: result <= 12'b011111001010;
   13992: result <= 12'b011111001010;
   13993: result <= 12'b011111001010;
   13994: result <= 12'b011111001010;
   13995: result <= 12'b011111001010;
   13996: result <= 12'b011111001010;
   13997: result <= 12'b011111001010;
   13998: result <= 12'b011111001010;
   13999: result <= 12'b011111001010;
   14000: result <= 12'b011111001010;
   14001: result <= 12'b011111001010;
   14002: result <= 12'b011111001010;
   14003: result <= 12'b011111001010;
   14004: result <= 12'b011111001010;
   14005: result <= 12'b011111001010;
   14006: result <= 12'b011111001011;
   14007: result <= 12'b011111001011;
   14008: result <= 12'b011111001011;
   14009: result <= 12'b011111001011;
   14010: result <= 12'b011111001011;
   14011: result <= 12'b011111001011;
   14012: result <= 12'b011111001011;
   14013: result <= 12'b011111001011;
   14014: result <= 12'b011111001011;
   14015: result <= 12'b011111001011;
   14016: result <= 12'b011111001011;
   14017: result <= 12'b011111001011;
   14018: result <= 12'b011111001011;
   14019: result <= 12'b011111001011;
   14020: result <= 12'b011111001011;
   14021: result <= 12'b011111001011;
   14022: result <= 12'b011111001011;
   14023: result <= 12'b011111001011;
   14024: result <= 12'b011111001011;
   14025: result <= 12'b011111001011;
   14026: result <= 12'b011111001011;
   14027: result <= 12'b011111001011;
   14028: result <= 12'b011111001011;
   14029: result <= 12'b011111001100;
   14030: result <= 12'b011111001100;
   14031: result <= 12'b011111001100;
   14032: result <= 12'b011111001100;
   14033: result <= 12'b011111001100;
   14034: result <= 12'b011111001100;
   14035: result <= 12'b011111001100;
   14036: result <= 12'b011111001100;
   14037: result <= 12'b011111001100;
   14038: result <= 12'b011111001100;
   14039: result <= 12'b011111001100;
   14040: result <= 12'b011111001100;
   14041: result <= 12'b011111001100;
   14042: result <= 12'b011111001100;
   14043: result <= 12'b011111001100;
   14044: result <= 12'b011111001100;
   14045: result <= 12'b011111001100;
   14046: result <= 12'b011111001100;
   14047: result <= 12'b011111001100;
   14048: result <= 12'b011111001100;
   14049: result <= 12'b011111001100;
   14050: result <= 12'b011111001100;
   14051: result <= 12'b011111001100;
   14052: result <= 12'b011111001101;
   14053: result <= 12'b011111001101;
   14054: result <= 12'b011111001101;
   14055: result <= 12'b011111001101;
   14056: result <= 12'b011111001101;
   14057: result <= 12'b011111001101;
   14058: result <= 12'b011111001101;
   14059: result <= 12'b011111001101;
   14060: result <= 12'b011111001101;
   14061: result <= 12'b011111001101;
   14062: result <= 12'b011111001101;
   14063: result <= 12'b011111001101;
   14064: result <= 12'b011111001101;
   14065: result <= 12'b011111001101;
   14066: result <= 12'b011111001101;
   14067: result <= 12'b011111001101;
   14068: result <= 12'b011111001101;
   14069: result <= 12'b011111001101;
   14070: result <= 12'b011111001101;
   14071: result <= 12'b011111001101;
   14072: result <= 12'b011111001101;
   14073: result <= 12'b011111001101;
   14074: result <= 12'b011111001101;
   14075: result <= 12'b011111001110;
   14076: result <= 12'b011111001110;
   14077: result <= 12'b011111001110;
   14078: result <= 12'b011111001110;
   14079: result <= 12'b011111001110;
   14080: result <= 12'b011111001110;
   14081: result <= 12'b011111001110;
   14082: result <= 12'b011111001110;
   14083: result <= 12'b011111001110;
   14084: result <= 12'b011111001110;
   14085: result <= 12'b011111001110;
   14086: result <= 12'b011111001110;
   14087: result <= 12'b011111001110;
   14088: result <= 12'b011111001110;
   14089: result <= 12'b011111001110;
   14090: result <= 12'b011111001110;
   14091: result <= 12'b011111001110;
   14092: result <= 12'b011111001110;
   14093: result <= 12'b011111001110;
   14094: result <= 12'b011111001110;
   14095: result <= 12'b011111001110;
   14096: result <= 12'b011111001110;
   14097: result <= 12'b011111001110;
   14098: result <= 12'b011111001111;
   14099: result <= 12'b011111001111;
   14100: result <= 12'b011111001111;
   14101: result <= 12'b011111001111;
   14102: result <= 12'b011111001111;
   14103: result <= 12'b011111001111;
   14104: result <= 12'b011111001111;
   14105: result <= 12'b011111001111;
   14106: result <= 12'b011111001111;
   14107: result <= 12'b011111001111;
   14108: result <= 12'b011111001111;
   14109: result <= 12'b011111001111;
   14110: result <= 12'b011111001111;
   14111: result <= 12'b011111001111;
   14112: result <= 12'b011111001111;
   14113: result <= 12'b011111001111;
   14114: result <= 12'b011111001111;
   14115: result <= 12'b011111001111;
   14116: result <= 12'b011111001111;
   14117: result <= 12'b011111001111;
   14118: result <= 12'b011111001111;
   14119: result <= 12'b011111001111;
   14120: result <= 12'b011111001111;
   14121: result <= 12'b011111001111;
   14122: result <= 12'b011111010000;
   14123: result <= 12'b011111010000;
   14124: result <= 12'b011111010000;
   14125: result <= 12'b011111010000;
   14126: result <= 12'b011111010000;
   14127: result <= 12'b011111010000;
   14128: result <= 12'b011111010000;
   14129: result <= 12'b011111010000;
   14130: result <= 12'b011111010000;
   14131: result <= 12'b011111010000;
   14132: result <= 12'b011111010000;
   14133: result <= 12'b011111010000;
   14134: result <= 12'b011111010000;
   14135: result <= 12'b011111010000;
   14136: result <= 12'b011111010000;
   14137: result <= 12'b011111010000;
   14138: result <= 12'b011111010000;
   14139: result <= 12'b011111010000;
   14140: result <= 12'b011111010000;
   14141: result <= 12'b011111010000;
   14142: result <= 12'b011111010000;
   14143: result <= 12'b011111010000;
   14144: result <= 12'b011111010000;
   14145: result <= 12'b011111010000;
   14146: result <= 12'b011111010001;
   14147: result <= 12'b011111010001;
   14148: result <= 12'b011111010001;
   14149: result <= 12'b011111010001;
   14150: result <= 12'b011111010001;
   14151: result <= 12'b011111010001;
   14152: result <= 12'b011111010001;
   14153: result <= 12'b011111010001;
   14154: result <= 12'b011111010001;
   14155: result <= 12'b011111010001;
   14156: result <= 12'b011111010001;
   14157: result <= 12'b011111010001;
   14158: result <= 12'b011111010001;
   14159: result <= 12'b011111010001;
   14160: result <= 12'b011111010001;
   14161: result <= 12'b011111010001;
   14162: result <= 12'b011111010001;
   14163: result <= 12'b011111010001;
   14164: result <= 12'b011111010001;
   14165: result <= 12'b011111010001;
   14166: result <= 12'b011111010001;
   14167: result <= 12'b011111010001;
   14168: result <= 12'b011111010001;
   14169: result <= 12'b011111010001;
   14170: result <= 12'b011111010010;
   14171: result <= 12'b011111010010;
   14172: result <= 12'b011111010010;
   14173: result <= 12'b011111010010;
   14174: result <= 12'b011111010010;
   14175: result <= 12'b011111010010;
   14176: result <= 12'b011111010010;
   14177: result <= 12'b011111010010;
   14178: result <= 12'b011111010010;
   14179: result <= 12'b011111010010;
   14180: result <= 12'b011111010010;
   14181: result <= 12'b011111010010;
   14182: result <= 12'b011111010010;
   14183: result <= 12'b011111010010;
   14184: result <= 12'b011111010010;
   14185: result <= 12'b011111010010;
   14186: result <= 12'b011111010010;
   14187: result <= 12'b011111010010;
   14188: result <= 12'b011111010010;
   14189: result <= 12'b011111010010;
   14190: result <= 12'b011111010010;
   14191: result <= 12'b011111010010;
   14192: result <= 12'b011111010010;
   14193: result <= 12'b011111010010;
   14194: result <= 12'b011111010011;
   14195: result <= 12'b011111010011;
   14196: result <= 12'b011111010011;
   14197: result <= 12'b011111010011;
   14198: result <= 12'b011111010011;
   14199: result <= 12'b011111010011;
   14200: result <= 12'b011111010011;
   14201: result <= 12'b011111010011;
   14202: result <= 12'b011111010011;
   14203: result <= 12'b011111010011;
   14204: result <= 12'b011111010011;
   14205: result <= 12'b011111010011;
   14206: result <= 12'b011111010011;
   14207: result <= 12'b011111010011;
   14208: result <= 12'b011111010011;
   14209: result <= 12'b011111010011;
   14210: result <= 12'b011111010011;
   14211: result <= 12'b011111010011;
   14212: result <= 12'b011111010011;
   14213: result <= 12'b011111010011;
   14214: result <= 12'b011111010011;
   14215: result <= 12'b011111010011;
   14216: result <= 12'b011111010011;
   14217: result <= 12'b011111010011;
   14218: result <= 12'b011111010011;
   14219: result <= 12'b011111010100;
   14220: result <= 12'b011111010100;
   14221: result <= 12'b011111010100;
   14222: result <= 12'b011111010100;
   14223: result <= 12'b011111010100;
   14224: result <= 12'b011111010100;
   14225: result <= 12'b011111010100;
   14226: result <= 12'b011111010100;
   14227: result <= 12'b011111010100;
   14228: result <= 12'b011111010100;
   14229: result <= 12'b011111010100;
   14230: result <= 12'b011111010100;
   14231: result <= 12'b011111010100;
   14232: result <= 12'b011111010100;
   14233: result <= 12'b011111010100;
   14234: result <= 12'b011111010100;
   14235: result <= 12'b011111010100;
   14236: result <= 12'b011111010100;
   14237: result <= 12'b011111010100;
   14238: result <= 12'b011111010100;
   14239: result <= 12'b011111010100;
   14240: result <= 12'b011111010100;
   14241: result <= 12'b011111010100;
   14242: result <= 12'b011111010100;
   14243: result <= 12'b011111010101;
   14244: result <= 12'b011111010101;
   14245: result <= 12'b011111010101;
   14246: result <= 12'b011111010101;
   14247: result <= 12'b011111010101;
   14248: result <= 12'b011111010101;
   14249: result <= 12'b011111010101;
   14250: result <= 12'b011111010101;
   14251: result <= 12'b011111010101;
   14252: result <= 12'b011111010101;
   14253: result <= 12'b011111010101;
   14254: result <= 12'b011111010101;
   14255: result <= 12'b011111010101;
   14256: result <= 12'b011111010101;
   14257: result <= 12'b011111010101;
   14258: result <= 12'b011111010101;
   14259: result <= 12'b011111010101;
   14260: result <= 12'b011111010101;
   14261: result <= 12'b011111010101;
   14262: result <= 12'b011111010101;
   14263: result <= 12'b011111010101;
   14264: result <= 12'b011111010101;
   14265: result <= 12'b011111010101;
   14266: result <= 12'b011111010101;
   14267: result <= 12'b011111010101;
   14268: result <= 12'b011111010110;
   14269: result <= 12'b011111010110;
   14270: result <= 12'b011111010110;
   14271: result <= 12'b011111010110;
   14272: result <= 12'b011111010110;
   14273: result <= 12'b011111010110;
   14274: result <= 12'b011111010110;
   14275: result <= 12'b011111010110;
   14276: result <= 12'b011111010110;
   14277: result <= 12'b011111010110;
   14278: result <= 12'b011111010110;
   14279: result <= 12'b011111010110;
   14280: result <= 12'b011111010110;
   14281: result <= 12'b011111010110;
   14282: result <= 12'b011111010110;
   14283: result <= 12'b011111010110;
   14284: result <= 12'b011111010110;
   14285: result <= 12'b011111010110;
   14286: result <= 12'b011111010110;
   14287: result <= 12'b011111010110;
   14288: result <= 12'b011111010110;
   14289: result <= 12'b011111010110;
   14290: result <= 12'b011111010110;
   14291: result <= 12'b011111010110;
   14292: result <= 12'b011111010110;
   14293: result <= 12'b011111010110;
   14294: result <= 12'b011111010111;
   14295: result <= 12'b011111010111;
   14296: result <= 12'b011111010111;
   14297: result <= 12'b011111010111;
   14298: result <= 12'b011111010111;
   14299: result <= 12'b011111010111;
   14300: result <= 12'b011111010111;
   14301: result <= 12'b011111010111;
   14302: result <= 12'b011111010111;
   14303: result <= 12'b011111010111;
   14304: result <= 12'b011111010111;
   14305: result <= 12'b011111010111;
   14306: result <= 12'b011111010111;
   14307: result <= 12'b011111010111;
   14308: result <= 12'b011111010111;
   14309: result <= 12'b011111010111;
   14310: result <= 12'b011111010111;
   14311: result <= 12'b011111010111;
   14312: result <= 12'b011111010111;
   14313: result <= 12'b011111010111;
   14314: result <= 12'b011111010111;
   14315: result <= 12'b011111010111;
   14316: result <= 12'b011111010111;
   14317: result <= 12'b011111010111;
   14318: result <= 12'b011111010111;
   14319: result <= 12'b011111010111;
   14320: result <= 12'b011111011000;
   14321: result <= 12'b011111011000;
   14322: result <= 12'b011111011000;
   14323: result <= 12'b011111011000;
   14324: result <= 12'b011111011000;
   14325: result <= 12'b011111011000;
   14326: result <= 12'b011111011000;
   14327: result <= 12'b011111011000;
   14328: result <= 12'b011111011000;
   14329: result <= 12'b011111011000;
   14330: result <= 12'b011111011000;
   14331: result <= 12'b011111011000;
   14332: result <= 12'b011111011000;
   14333: result <= 12'b011111011000;
   14334: result <= 12'b011111011000;
   14335: result <= 12'b011111011000;
   14336: result <= 12'b011111011000;
   14337: result <= 12'b011111011000;
   14338: result <= 12'b011111011000;
   14339: result <= 12'b011111011000;
   14340: result <= 12'b011111011000;
   14341: result <= 12'b011111011000;
   14342: result <= 12'b011111011000;
   14343: result <= 12'b011111011000;
   14344: result <= 12'b011111011000;
   14345: result <= 12'b011111011000;
   14346: result <= 12'b011111011001;
   14347: result <= 12'b011111011001;
   14348: result <= 12'b011111011001;
   14349: result <= 12'b011111011001;
   14350: result <= 12'b011111011001;
   14351: result <= 12'b011111011001;
   14352: result <= 12'b011111011001;
   14353: result <= 12'b011111011001;
   14354: result <= 12'b011111011001;
   14355: result <= 12'b011111011001;
   14356: result <= 12'b011111011001;
   14357: result <= 12'b011111011001;
   14358: result <= 12'b011111011001;
   14359: result <= 12'b011111011001;
   14360: result <= 12'b011111011001;
   14361: result <= 12'b011111011001;
   14362: result <= 12'b011111011001;
   14363: result <= 12'b011111011001;
   14364: result <= 12'b011111011001;
   14365: result <= 12'b011111011001;
   14366: result <= 12'b011111011001;
   14367: result <= 12'b011111011001;
   14368: result <= 12'b011111011001;
   14369: result <= 12'b011111011001;
   14370: result <= 12'b011111011001;
   14371: result <= 12'b011111011001;
   14372: result <= 12'b011111011010;
   14373: result <= 12'b011111011010;
   14374: result <= 12'b011111011010;
   14375: result <= 12'b011111011010;
   14376: result <= 12'b011111011010;
   14377: result <= 12'b011111011010;
   14378: result <= 12'b011111011010;
   14379: result <= 12'b011111011010;
   14380: result <= 12'b011111011010;
   14381: result <= 12'b011111011010;
   14382: result <= 12'b011111011010;
   14383: result <= 12'b011111011010;
   14384: result <= 12'b011111011010;
   14385: result <= 12'b011111011010;
   14386: result <= 12'b011111011010;
   14387: result <= 12'b011111011010;
   14388: result <= 12'b011111011010;
   14389: result <= 12'b011111011010;
   14390: result <= 12'b011111011010;
   14391: result <= 12'b011111011010;
   14392: result <= 12'b011111011010;
   14393: result <= 12'b011111011010;
   14394: result <= 12'b011111011010;
   14395: result <= 12'b011111011010;
   14396: result <= 12'b011111011010;
   14397: result <= 12'b011111011010;
   14398: result <= 12'b011111011010;
   14399: result <= 12'b011111011011;
   14400: result <= 12'b011111011011;
   14401: result <= 12'b011111011011;
   14402: result <= 12'b011111011011;
   14403: result <= 12'b011111011011;
   14404: result <= 12'b011111011011;
   14405: result <= 12'b011111011011;
   14406: result <= 12'b011111011011;
   14407: result <= 12'b011111011011;
   14408: result <= 12'b011111011011;
   14409: result <= 12'b011111011011;
   14410: result <= 12'b011111011011;
   14411: result <= 12'b011111011011;
   14412: result <= 12'b011111011011;
   14413: result <= 12'b011111011011;
   14414: result <= 12'b011111011011;
   14415: result <= 12'b011111011011;
   14416: result <= 12'b011111011011;
   14417: result <= 12'b011111011011;
   14418: result <= 12'b011111011011;
   14419: result <= 12'b011111011011;
   14420: result <= 12'b011111011011;
   14421: result <= 12'b011111011011;
   14422: result <= 12'b011111011011;
   14423: result <= 12'b011111011011;
   14424: result <= 12'b011111011011;
   14425: result <= 12'b011111011011;
   14426: result <= 12'b011111011100;
   14427: result <= 12'b011111011100;
   14428: result <= 12'b011111011100;
   14429: result <= 12'b011111011100;
   14430: result <= 12'b011111011100;
   14431: result <= 12'b011111011100;
   14432: result <= 12'b011111011100;
   14433: result <= 12'b011111011100;
   14434: result <= 12'b011111011100;
   14435: result <= 12'b011111011100;
   14436: result <= 12'b011111011100;
   14437: result <= 12'b011111011100;
   14438: result <= 12'b011111011100;
   14439: result <= 12'b011111011100;
   14440: result <= 12'b011111011100;
   14441: result <= 12'b011111011100;
   14442: result <= 12'b011111011100;
   14443: result <= 12'b011111011100;
   14444: result <= 12'b011111011100;
   14445: result <= 12'b011111011100;
   14446: result <= 12'b011111011100;
   14447: result <= 12'b011111011100;
   14448: result <= 12'b011111011100;
   14449: result <= 12'b011111011100;
   14450: result <= 12'b011111011100;
   14451: result <= 12'b011111011100;
   14452: result <= 12'b011111011100;
   14453: result <= 12'b011111011101;
   14454: result <= 12'b011111011101;
   14455: result <= 12'b011111011101;
   14456: result <= 12'b011111011101;
   14457: result <= 12'b011111011101;
   14458: result <= 12'b011111011101;
   14459: result <= 12'b011111011101;
   14460: result <= 12'b011111011101;
   14461: result <= 12'b011111011101;
   14462: result <= 12'b011111011101;
   14463: result <= 12'b011111011101;
   14464: result <= 12'b011111011101;
   14465: result <= 12'b011111011101;
   14466: result <= 12'b011111011101;
   14467: result <= 12'b011111011101;
   14468: result <= 12'b011111011101;
   14469: result <= 12'b011111011101;
   14470: result <= 12'b011111011101;
   14471: result <= 12'b011111011101;
   14472: result <= 12'b011111011101;
   14473: result <= 12'b011111011101;
   14474: result <= 12'b011111011101;
   14475: result <= 12'b011111011101;
   14476: result <= 12'b011111011101;
   14477: result <= 12'b011111011101;
   14478: result <= 12'b011111011101;
   14479: result <= 12'b011111011101;
   14480: result <= 12'b011111011101;
   14481: result <= 12'b011111011110;
   14482: result <= 12'b011111011110;
   14483: result <= 12'b011111011110;
   14484: result <= 12'b011111011110;
   14485: result <= 12'b011111011110;
   14486: result <= 12'b011111011110;
   14487: result <= 12'b011111011110;
   14488: result <= 12'b011111011110;
   14489: result <= 12'b011111011110;
   14490: result <= 12'b011111011110;
   14491: result <= 12'b011111011110;
   14492: result <= 12'b011111011110;
   14493: result <= 12'b011111011110;
   14494: result <= 12'b011111011110;
   14495: result <= 12'b011111011110;
   14496: result <= 12'b011111011110;
   14497: result <= 12'b011111011110;
   14498: result <= 12'b011111011110;
   14499: result <= 12'b011111011110;
   14500: result <= 12'b011111011110;
   14501: result <= 12'b011111011110;
   14502: result <= 12'b011111011110;
   14503: result <= 12'b011111011110;
   14504: result <= 12'b011111011110;
   14505: result <= 12'b011111011110;
   14506: result <= 12'b011111011110;
   14507: result <= 12'b011111011110;
   14508: result <= 12'b011111011110;
   14509: result <= 12'b011111011110;
   14510: result <= 12'b011111011111;
   14511: result <= 12'b011111011111;
   14512: result <= 12'b011111011111;
   14513: result <= 12'b011111011111;
   14514: result <= 12'b011111011111;
   14515: result <= 12'b011111011111;
   14516: result <= 12'b011111011111;
   14517: result <= 12'b011111011111;
   14518: result <= 12'b011111011111;
   14519: result <= 12'b011111011111;
   14520: result <= 12'b011111011111;
   14521: result <= 12'b011111011111;
   14522: result <= 12'b011111011111;
   14523: result <= 12'b011111011111;
   14524: result <= 12'b011111011111;
   14525: result <= 12'b011111011111;
   14526: result <= 12'b011111011111;
   14527: result <= 12'b011111011111;
   14528: result <= 12'b011111011111;
   14529: result <= 12'b011111011111;
   14530: result <= 12'b011111011111;
   14531: result <= 12'b011111011111;
   14532: result <= 12'b011111011111;
   14533: result <= 12'b011111011111;
   14534: result <= 12'b011111011111;
   14535: result <= 12'b011111011111;
   14536: result <= 12'b011111011111;
   14537: result <= 12'b011111011111;
   14538: result <= 12'b011111100000;
   14539: result <= 12'b011111100000;
   14540: result <= 12'b011111100000;
   14541: result <= 12'b011111100000;
   14542: result <= 12'b011111100000;
   14543: result <= 12'b011111100000;
   14544: result <= 12'b011111100000;
   14545: result <= 12'b011111100000;
   14546: result <= 12'b011111100000;
   14547: result <= 12'b011111100000;
   14548: result <= 12'b011111100000;
   14549: result <= 12'b011111100000;
   14550: result <= 12'b011111100000;
   14551: result <= 12'b011111100000;
   14552: result <= 12'b011111100000;
   14553: result <= 12'b011111100000;
   14554: result <= 12'b011111100000;
   14555: result <= 12'b011111100000;
   14556: result <= 12'b011111100000;
   14557: result <= 12'b011111100000;
   14558: result <= 12'b011111100000;
   14559: result <= 12'b011111100000;
   14560: result <= 12'b011111100000;
   14561: result <= 12'b011111100000;
   14562: result <= 12'b011111100000;
   14563: result <= 12'b011111100000;
   14564: result <= 12'b011111100000;
   14565: result <= 12'b011111100000;
   14566: result <= 12'b011111100000;
   14567: result <= 12'b011111100001;
   14568: result <= 12'b011111100001;
   14569: result <= 12'b011111100001;
   14570: result <= 12'b011111100001;
   14571: result <= 12'b011111100001;
   14572: result <= 12'b011111100001;
   14573: result <= 12'b011111100001;
   14574: result <= 12'b011111100001;
   14575: result <= 12'b011111100001;
   14576: result <= 12'b011111100001;
   14577: result <= 12'b011111100001;
   14578: result <= 12'b011111100001;
   14579: result <= 12'b011111100001;
   14580: result <= 12'b011111100001;
   14581: result <= 12'b011111100001;
   14582: result <= 12'b011111100001;
   14583: result <= 12'b011111100001;
   14584: result <= 12'b011111100001;
   14585: result <= 12'b011111100001;
   14586: result <= 12'b011111100001;
   14587: result <= 12'b011111100001;
   14588: result <= 12'b011111100001;
   14589: result <= 12'b011111100001;
   14590: result <= 12'b011111100001;
   14591: result <= 12'b011111100001;
   14592: result <= 12'b011111100001;
   14593: result <= 12'b011111100001;
   14594: result <= 12'b011111100001;
   14595: result <= 12'b011111100001;
   14596: result <= 12'b011111100001;
   14597: result <= 12'b011111100010;
   14598: result <= 12'b011111100010;
   14599: result <= 12'b011111100010;
   14600: result <= 12'b011111100010;
   14601: result <= 12'b011111100010;
   14602: result <= 12'b011111100010;
   14603: result <= 12'b011111100010;
   14604: result <= 12'b011111100010;
   14605: result <= 12'b011111100010;
   14606: result <= 12'b011111100010;
   14607: result <= 12'b011111100010;
   14608: result <= 12'b011111100010;
   14609: result <= 12'b011111100010;
   14610: result <= 12'b011111100010;
   14611: result <= 12'b011111100010;
   14612: result <= 12'b011111100010;
   14613: result <= 12'b011111100010;
   14614: result <= 12'b011111100010;
   14615: result <= 12'b011111100010;
   14616: result <= 12'b011111100010;
   14617: result <= 12'b011111100010;
   14618: result <= 12'b011111100010;
   14619: result <= 12'b011111100010;
   14620: result <= 12'b011111100010;
   14621: result <= 12'b011111100010;
   14622: result <= 12'b011111100010;
   14623: result <= 12'b011111100010;
   14624: result <= 12'b011111100010;
   14625: result <= 12'b011111100010;
   14626: result <= 12'b011111100010;
   14627: result <= 12'b011111100011;
   14628: result <= 12'b011111100011;
   14629: result <= 12'b011111100011;
   14630: result <= 12'b011111100011;
   14631: result <= 12'b011111100011;
   14632: result <= 12'b011111100011;
   14633: result <= 12'b011111100011;
   14634: result <= 12'b011111100011;
   14635: result <= 12'b011111100011;
   14636: result <= 12'b011111100011;
   14637: result <= 12'b011111100011;
   14638: result <= 12'b011111100011;
   14639: result <= 12'b011111100011;
   14640: result <= 12'b011111100011;
   14641: result <= 12'b011111100011;
   14642: result <= 12'b011111100011;
   14643: result <= 12'b011111100011;
   14644: result <= 12'b011111100011;
   14645: result <= 12'b011111100011;
   14646: result <= 12'b011111100011;
   14647: result <= 12'b011111100011;
   14648: result <= 12'b011111100011;
   14649: result <= 12'b011111100011;
   14650: result <= 12'b011111100011;
   14651: result <= 12'b011111100011;
   14652: result <= 12'b011111100011;
   14653: result <= 12'b011111100011;
   14654: result <= 12'b011111100011;
   14655: result <= 12'b011111100011;
   14656: result <= 12'b011111100011;
   14657: result <= 12'b011111100011;
   14658: result <= 12'b011111100100;
   14659: result <= 12'b011111100100;
   14660: result <= 12'b011111100100;
   14661: result <= 12'b011111100100;
   14662: result <= 12'b011111100100;
   14663: result <= 12'b011111100100;
   14664: result <= 12'b011111100100;
   14665: result <= 12'b011111100100;
   14666: result <= 12'b011111100100;
   14667: result <= 12'b011111100100;
   14668: result <= 12'b011111100100;
   14669: result <= 12'b011111100100;
   14670: result <= 12'b011111100100;
   14671: result <= 12'b011111100100;
   14672: result <= 12'b011111100100;
   14673: result <= 12'b011111100100;
   14674: result <= 12'b011111100100;
   14675: result <= 12'b011111100100;
   14676: result <= 12'b011111100100;
   14677: result <= 12'b011111100100;
   14678: result <= 12'b011111100100;
   14679: result <= 12'b011111100100;
   14680: result <= 12'b011111100100;
   14681: result <= 12'b011111100100;
   14682: result <= 12'b011111100100;
   14683: result <= 12'b011111100100;
   14684: result <= 12'b011111100100;
   14685: result <= 12'b011111100100;
   14686: result <= 12'b011111100100;
   14687: result <= 12'b011111100100;
   14688: result <= 12'b011111100100;
   14689: result <= 12'b011111100101;
   14690: result <= 12'b011111100101;
   14691: result <= 12'b011111100101;
   14692: result <= 12'b011111100101;
   14693: result <= 12'b011111100101;
   14694: result <= 12'b011111100101;
   14695: result <= 12'b011111100101;
   14696: result <= 12'b011111100101;
   14697: result <= 12'b011111100101;
   14698: result <= 12'b011111100101;
   14699: result <= 12'b011111100101;
   14700: result <= 12'b011111100101;
   14701: result <= 12'b011111100101;
   14702: result <= 12'b011111100101;
   14703: result <= 12'b011111100101;
   14704: result <= 12'b011111100101;
   14705: result <= 12'b011111100101;
   14706: result <= 12'b011111100101;
   14707: result <= 12'b011111100101;
   14708: result <= 12'b011111100101;
   14709: result <= 12'b011111100101;
   14710: result <= 12'b011111100101;
   14711: result <= 12'b011111100101;
   14712: result <= 12'b011111100101;
   14713: result <= 12'b011111100101;
   14714: result <= 12'b011111100101;
   14715: result <= 12'b011111100101;
   14716: result <= 12'b011111100101;
   14717: result <= 12'b011111100101;
   14718: result <= 12'b011111100101;
   14719: result <= 12'b011111100101;
   14720: result <= 12'b011111100101;
   14721: result <= 12'b011111100110;
   14722: result <= 12'b011111100110;
   14723: result <= 12'b011111100110;
   14724: result <= 12'b011111100110;
   14725: result <= 12'b011111100110;
   14726: result <= 12'b011111100110;
   14727: result <= 12'b011111100110;
   14728: result <= 12'b011111100110;
   14729: result <= 12'b011111100110;
   14730: result <= 12'b011111100110;
   14731: result <= 12'b011111100110;
   14732: result <= 12'b011111100110;
   14733: result <= 12'b011111100110;
   14734: result <= 12'b011111100110;
   14735: result <= 12'b011111100110;
   14736: result <= 12'b011111100110;
   14737: result <= 12'b011111100110;
   14738: result <= 12'b011111100110;
   14739: result <= 12'b011111100110;
   14740: result <= 12'b011111100110;
   14741: result <= 12'b011111100110;
   14742: result <= 12'b011111100110;
   14743: result <= 12'b011111100110;
   14744: result <= 12'b011111100110;
   14745: result <= 12'b011111100110;
   14746: result <= 12'b011111100110;
   14747: result <= 12'b011111100110;
   14748: result <= 12'b011111100110;
   14749: result <= 12'b011111100110;
   14750: result <= 12'b011111100110;
   14751: result <= 12'b011111100110;
   14752: result <= 12'b011111100110;
   14753: result <= 12'b011111100111;
   14754: result <= 12'b011111100111;
   14755: result <= 12'b011111100111;
   14756: result <= 12'b011111100111;
   14757: result <= 12'b011111100111;
   14758: result <= 12'b011111100111;
   14759: result <= 12'b011111100111;
   14760: result <= 12'b011111100111;
   14761: result <= 12'b011111100111;
   14762: result <= 12'b011111100111;
   14763: result <= 12'b011111100111;
   14764: result <= 12'b011111100111;
   14765: result <= 12'b011111100111;
   14766: result <= 12'b011111100111;
   14767: result <= 12'b011111100111;
   14768: result <= 12'b011111100111;
   14769: result <= 12'b011111100111;
   14770: result <= 12'b011111100111;
   14771: result <= 12'b011111100111;
   14772: result <= 12'b011111100111;
   14773: result <= 12'b011111100111;
   14774: result <= 12'b011111100111;
   14775: result <= 12'b011111100111;
   14776: result <= 12'b011111100111;
   14777: result <= 12'b011111100111;
   14778: result <= 12'b011111100111;
   14779: result <= 12'b011111100111;
   14780: result <= 12'b011111100111;
   14781: result <= 12'b011111100111;
   14782: result <= 12'b011111100111;
   14783: result <= 12'b011111100111;
   14784: result <= 12'b011111100111;
   14785: result <= 12'b011111100111;
   14786: result <= 12'b011111101000;
   14787: result <= 12'b011111101000;
   14788: result <= 12'b011111101000;
   14789: result <= 12'b011111101000;
   14790: result <= 12'b011111101000;
   14791: result <= 12'b011111101000;
   14792: result <= 12'b011111101000;
   14793: result <= 12'b011111101000;
   14794: result <= 12'b011111101000;
   14795: result <= 12'b011111101000;
   14796: result <= 12'b011111101000;
   14797: result <= 12'b011111101000;
   14798: result <= 12'b011111101000;
   14799: result <= 12'b011111101000;
   14800: result <= 12'b011111101000;
   14801: result <= 12'b011111101000;
   14802: result <= 12'b011111101000;
   14803: result <= 12'b011111101000;
   14804: result <= 12'b011111101000;
   14805: result <= 12'b011111101000;
   14806: result <= 12'b011111101000;
   14807: result <= 12'b011111101000;
   14808: result <= 12'b011111101000;
   14809: result <= 12'b011111101000;
   14810: result <= 12'b011111101000;
   14811: result <= 12'b011111101000;
   14812: result <= 12'b011111101000;
   14813: result <= 12'b011111101000;
   14814: result <= 12'b011111101000;
   14815: result <= 12'b011111101000;
   14816: result <= 12'b011111101000;
   14817: result <= 12'b011111101000;
   14818: result <= 12'b011111101000;
   14819: result <= 12'b011111101000;
   14820: result <= 12'b011111101001;
   14821: result <= 12'b011111101001;
   14822: result <= 12'b011111101001;
   14823: result <= 12'b011111101001;
   14824: result <= 12'b011111101001;
   14825: result <= 12'b011111101001;
   14826: result <= 12'b011111101001;
   14827: result <= 12'b011111101001;
   14828: result <= 12'b011111101001;
   14829: result <= 12'b011111101001;
   14830: result <= 12'b011111101001;
   14831: result <= 12'b011111101001;
   14832: result <= 12'b011111101001;
   14833: result <= 12'b011111101001;
   14834: result <= 12'b011111101001;
   14835: result <= 12'b011111101001;
   14836: result <= 12'b011111101001;
   14837: result <= 12'b011111101001;
   14838: result <= 12'b011111101001;
   14839: result <= 12'b011111101001;
   14840: result <= 12'b011111101001;
   14841: result <= 12'b011111101001;
   14842: result <= 12'b011111101001;
   14843: result <= 12'b011111101001;
   14844: result <= 12'b011111101001;
   14845: result <= 12'b011111101001;
   14846: result <= 12'b011111101001;
   14847: result <= 12'b011111101001;
   14848: result <= 12'b011111101001;
   14849: result <= 12'b011111101001;
   14850: result <= 12'b011111101001;
   14851: result <= 12'b011111101001;
   14852: result <= 12'b011111101001;
   14853: result <= 12'b011111101001;
   14854: result <= 12'b011111101010;
   14855: result <= 12'b011111101010;
   14856: result <= 12'b011111101010;
   14857: result <= 12'b011111101010;
   14858: result <= 12'b011111101010;
   14859: result <= 12'b011111101010;
   14860: result <= 12'b011111101010;
   14861: result <= 12'b011111101010;
   14862: result <= 12'b011111101010;
   14863: result <= 12'b011111101010;
   14864: result <= 12'b011111101010;
   14865: result <= 12'b011111101010;
   14866: result <= 12'b011111101010;
   14867: result <= 12'b011111101010;
   14868: result <= 12'b011111101010;
   14869: result <= 12'b011111101010;
   14870: result <= 12'b011111101010;
   14871: result <= 12'b011111101010;
   14872: result <= 12'b011111101010;
   14873: result <= 12'b011111101010;
   14874: result <= 12'b011111101010;
   14875: result <= 12'b011111101010;
   14876: result <= 12'b011111101010;
   14877: result <= 12'b011111101010;
   14878: result <= 12'b011111101010;
   14879: result <= 12'b011111101010;
   14880: result <= 12'b011111101010;
   14881: result <= 12'b011111101010;
   14882: result <= 12'b011111101010;
   14883: result <= 12'b011111101010;
   14884: result <= 12'b011111101010;
   14885: result <= 12'b011111101010;
   14886: result <= 12'b011111101010;
   14887: result <= 12'b011111101010;
   14888: result <= 12'b011111101010;
   14889: result <= 12'b011111101010;
   14890: result <= 12'b011111101011;
   14891: result <= 12'b011111101011;
   14892: result <= 12'b011111101011;
   14893: result <= 12'b011111101011;
   14894: result <= 12'b011111101011;
   14895: result <= 12'b011111101011;
   14896: result <= 12'b011111101011;
   14897: result <= 12'b011111101011;
   14898: result <= 12'b011111101011;
   14899: result <= 12'b011111101011;
   14900: result <= 12'b011111101011;
   14901: result <= 12'b011111101011;
   14902: result <= 12'b011111101011;
   14903: result <= 12'b011111101011;
   14904: result <= 12'b011111101011;
   14905: result <= 12'b011111101011;
   14906: result <= 12'b011111101011;
   14907: result <= 12'b011111101011;
   14908: result <= 12'b011111101011;
   14909: result <= 12'b011111101011;
   14910: result <= 12'b011111101011;
   14911: result <= 12'b011111101011;
   14912: result <= 12'b011111101011;
   14913: result <= 12'b011111101011;
   14914: result <= 12'b011111101011;
   14915: result <= 12'b011111101011;
   14916: result <= 12'b011111101011;
   14917: result <= 12'b011111101011;
   14918: result <= 12'b011111101011;
   14919: result <= 12'b011111101011;
   14920: result <= 12'b011111101011;
   14921: result <= 12'b011111101011;
   14922: result <= 12'b011111101011;
   14923: result <= 12'b011111101011;
   14924: result <= 12'b011111101011;
   14925: result <= 12'b011111101011;
   14926: result <= 12'b011111101100;
   14927: result <= 12'b011111101100;
   14928: result <= 12'b011111101100;
   14929: result <= 12'b011111101100;
   14930: result <= 12'b011111101100;
   14931: result <= 12'b011111101100;
   14932: result <= 12'b011111101100;
   14933: result <= 12'b011111101100;
   14934: result <= 12'b011111101100;
   14935: result <= 12'b011111101100;
   14936: result <= 12'b011111101100;
   14937: result <= 12'b011111101100;
   14938: result <= 12'b011111101100;
   14939: result <= 12'b011111101100;
   14940: result <= 12'b011111101100;
   14941: result <= 12'b011111101100;
   14942: result <= 12'b011111101100;
   14943: result <= 12'b011111101100;
   14944: result <= 12'b011111101100;
   14945: result <= 12'b011111101100;
   14946: result <= 12'b011111101100;
   14947: result <= 12'b011111101100;
   14948: result <= 12'b011111101100;
   14949: result <= 12'b011111101100;
   14950: result <= 12'b011111101100;
   14951: result <= 12'b011111101100;
   14952: result <= 12'b011111101100;
   14953: result <= 12'b011111101100;
   14954: result <= 12'b011111101100;
   14955: result <= 12'b011111101100;
   14956: result <= 12'b011111101100;
   14957: result <= 12'b011111101100;
   14958: result <= 12'b011111101100;
   14959: result <= 12'b011111101100;
   14960: result <= 12'b011111101100;
   14961: result <= 12'b011111101100;
   14962: result <= 12'b011111101100;
   14963: result <= 12'b011111101101;
   14964: result <= 12'b011111101101;
   14965: result <= 12'b011111101101;
   14966: result <= 12'b011111101101;
   14967: result <= 12'b011111101101;
   14968: result <= 12'b011111101101;
   14969: result <= 12'b011111101101;
   14970: result <= 12'b011111101101;
   14971: result <= 12'b011111101101;
   14972: result <= 12'b011111101101;
   14973: result <= 12'b011111101101;
   14974: result <= 12'b011111101101;
   14975: result <= 12'b011111101101;
   14976: result <= 12'b011111101101;
   14977: result <= 12'b011111101101;
   14978: result <= 12'b011111101101;
   14979: result <= 12'b011111101101;
   14980: result <= 12'b011111101101;
   14981: result <= 12'b011111101101;
   14982: result <= 12'b011111101101;
   14983: result <= 12'b011111101101;
   14984: result <= 12'b011111101101;
   14985: result <= 12'b011111101101;
   14986: result <= 12'b011111101101;
   14987: result <= 12'b011111101101;
   14988: result <= 12'b011111101101;
   14989: result <= 12'b011111101101;
   14990: result <= 12'b011111101101;
   14991: result <= 12'b011111101101;
   14992: result <= 12'b011111101101;
   14993: result <= 12'b011111101101;
   14994: result <= 12'b011111101101;
   14995: result <= 12'b011111101101;
   14996: result <= 12'b011111101101;
   14997: result <= 12'b011111101101;
   14998: result <= 12'b011111101101;
   14999: result <= 12'b011111101101;
   15000: result <= 12'b011111101101;
   15001: result <= 12'b011111101110;
   15002: result <= 12'b011111101110;
   15003: result <= 12'b011111101110;
   15004: result <= 12'b011111101110;
   15005: result <= 12'b011111101110;
   15006: result <= 12'b011111101110;
   15007: result <= 12'b011111101110;
   15008: result <= 12'b011111101110;
   15009: result <= 12'b011111101110;
   15010: result <= 12'b011111101110;
   15011: result <= 12'b011111101110;
   15012: result <= 12'b011111101110;
   15013: result <= 12'b011111101110;
   15014: result <= 12'b011111101110;
   15015: result <= 12'b011111101110;
   15016: result <= 12'b011111101110;
   15017: result <= 12'b011111101110;
   15018: result <= 12'b011111101110;
   15019: result <= 12'b011111101110;
   15020: result <= 12'b011111101110;
   15021: result <= 12'b011111101110;
   15022: result <= 12'b011111101110;
   15023: result <= 12'b011111101110;
   15024: result <= 12'b011111101110;
   15025: result <= 12'b011111101110;
   15026: result <= 12'b011111101110;
   15027: result <= 12'b011111101110;
   15028: result <= 12'b011111101110;
   15029: result <= 12'b011111101110;
   15030: result <= 12'b011111101110;
   15031: result <= 12'b011111101110;
   15032: result <= 12'b011111101110;
   15033: result <= 12'b011111101110;
   15034: result <= 12'b011111101110;
   15035: result <= 12'b011111101110;
   15036: result <= 12'b011111101110;
   15037: result <= 12'b011111101110;
   15038: result <= 12'b011111101110;
   15039: result <= 12'b011111101110;
   15040: result <= 12'b011111101111;
   15041: result <= 12'b011111101111;
   15042: result <= 12'b011111101111;
   15043: result <= 12'b011111101111;
   15044: result <= 12'b011111101111;
   15045: result <= 12'b011111101111;
   15046: result <= 12'b011111101111;
   15047: result <= 12'b011111101111;
   15048: result <= 12'b011111101111;
   15049: result <= 12'b011111101111;
   15050: result <= 12'b011111101111;
   15051: result <= 12'b011111101111;
   15052: result <= 12'b011111101111;
   15053: result <= 12'b011111101111;
   15054: result <= 12'b011111101111;
   15055: result <= 12'b011111101111;
   15056: result <= 12'b011111101111;
   15057: result <= 12'b011111101111;
   15058: result <= 12'b011111101111;
   15059: result <= 12'b011111101111;
   15060: result <= 12'b011111101111;
   15061: result <= 12'b011111101111;
   15062: result <= 12'b011111101111;
   15063: result <= 12'b011111101111;
   15064: result <= 12'b011111101111;
   15065: result <= 12'b011111101111;
   15066: result <= 12'b011111101111;
   15067: result <= 12'b011111101111;
   15068: result <= 12'b011111101111;
   15069: result <= 12'b011111101111;
   15070: result <= 12'b011111101111;
   15071: result <= 12'b011111101111;
   15072: result <= 12'b011111101111;
   15073: result <= 12'b011111101111;
   15074: result <= 12'b011111101111;
   15075: result <= 12'b011111101111;
   15076: result <= 12'b011111101111;
   15077: result <= 12'b011111101111;
   15078: result <= 12'b011111101111;
   15079: result <= 12'b011111101111;
   15080: result <= 12'b011111110000;
   15081: result <= 12'b011111110000;
   15082: result <= 12'b011111110000;
   15083: result <= 12'b011111110000;
   15084: result <= 12'b011111110000;
   15085: result <= 12'b011111110000;
   15086: result <= 12'b011111110000;
   15087: result <= 12'b011111110000;
   15088: result <= 12'b011111110000;
   15089: result <= 12'b011111110000;
   15090: result <= 12'b011111110000;
   15091: result <= 12'b011111110000;
   15092: result <= 12'b011111110000;
   15093: result <= 12'b011111110000;
   15094: result <= 12'b011111110000;
   15095: result <= 12'b011111110000;
   15096: result <= 12'b011111110000;
   15097: result <= 12'b011111110000;
   15098: result <= 12'b011111110000;
   15099: result <= 12'b011111110000;
   15100: result <= 12'b011111110000;
   15101: result <= 12'b011111110000;
   15102: result <= 12'b011111110000;
   15103: result <= 12'b011111110000;
   15104: result <= 12'b011111110000;
   15105: result <= 12'b011111110000;
   15106: result <= 12'b011111110000;
   15107: result <= 12'b011111110000;
   15108: result <= 12'b011111110000;
   15109: result <= 12'b011111110000;
   15110: result <= 12'b011111110000;
   15111: result <= 12'b011111110000;
   15112: result <= 12'b011111110000;
   15113: result <= 12'b011111110000;
   15114: result <= 12'b011111110000;
   15115: result <= 12'b011111110000;
   15116: result <= 12'b011111110000;
   15117: result <= 12'b011111110000;
   15118: result <= 12'b011111110000;
   15119: result <= 12'b011111110000;
   15120: result <= 12'b011111110000;
   15121: result <= 12'b011111110001;
   15122: result <= 12'b011111110001;
   15123: result <= 12'b011111110001;
   15124: result <= 12'b011111110001;
   15125: result <= 12'b011111110001;
   15126: result <= 12'b011111110001;
   15127: result <= 12'b011111110001;
   15128: result <= 12'b011111110001;
   15129: result <= 12'b011111110001;
   15130: result <= 12'b011111110001;
   15131: result <= 12'b011111110001;
   15132: result <= 12'b011111110001;
   15133: result <= 12'b011111110001;
   15134: result <= 12'b011111110001;
   15135: result <= 12'b011111110001;
   15136: result <= 12'b011111110001;
   15137: result <= 12'b011111110001;
   15138: result <= 12'b011111110001;
   15139: result <= 12'b011111110001;
   15140: result <= 12'b011111110001;
   15141: result <= 12'b011111110001;
   15142: result <= 12'b011111110001;
   15143: result <= 12'b011111110001;
   15144: result <= 12'b011111110001;
   15145: result <= 12'b011111110001;
   15146: result <= 12'b011111110001;
   15147: result <= 12'b011111110001;
   15148: result <= 12'b011111110001;
   15149: result <= 12'b011111110001;
   15150: result <= 12'b011111110001;
   15151: result <= 12'b011111110001;
   15152: result <= 12'b011111110001;
   15153: result <= 12'b011111110001;
   15154: result <= 12'b011111110001;
   15155: result <= 12'b011111110001;
   15156: result <= 12'b011111110001;
   15157: result <= 12'b011111110001;
   15158: result <= 12'b011111110001;
   15159: result <= 12'b011111110001;
   15160: result <= 12'b011111110001;
   15161: result <= 12'b011111110001;
   15162: result <= 12'b011111110001;
   15163: result <= 12'b011111110001;
   15164: result <= 12'b011111110010;
   15165: result <= 12'b011111110010;
   15166: result <= 12'b011111110010;
   15167: result <= 12'b011111110010;
   15168: result <= 12'b011111110010;
   15169: result <= 12'b011111110010;
   15170: result <= 12'b011111110010;
   15171: result <= 12'b011111110010;
   15172: result <= 12'b011111110010;
   15173: result <= 12'b011111110010;
   15174: result <= 12'b011111110010;
   15175: result <= 12'b011111110010;
   15176: result <= 12'b011111110010;
   15177: result <= 12'b011111110010;
   15178: result <= 12'b011111110010;
   15179: result <= 12'b011111110010;
   15180: result <= 12'b011111110010;
   15181: result <= 12'b011111110010;
   15182: result <= 12'b011111110010;
   15183: result <= 12'b011111110010;
   15184: result <= 12'b011111110010;
   15185: result <= 12'b011111110010;
   15186: result <= 12'b011111110010;
   15187: result <= 12'b011111110010;
   15188: result <= 12'b011111110010;
   15189: result <= 12'b011111110010;
   15190: result <= 12'b011111110010;
   15191: result <= 12'b011111110010;
   15192: result <= 12'b011111110010;
   15193: result <= 12'b011111110010;
   15194: result <= 12'b011111110010;
   15195: result <= 12'b011111110010;
   15196: result <= 12'b011111110010;
   15197: result <= 12'b011111110010;
   15198: result <= 12'b011111110010;
   15199: result <= 12'b011111110010;
   15200: result <= 12'b011111110010;
   15201: result <= 12'b011111110010;
   15202: result <= 12'b011111110010;
   15203: result <= 12'b011111110010;
   15204: result <= 12'b011111110010;
   15205: result <= 12'b011111110010;
   15206: result <= 12'b011111110010;
   15207: result <= 12'b011111110010;
   15208: result <= 12'b011111110010;
   15209: result <= 12'b011111110011;
   15210: result <= 12'b011111110011;
   15211: result <= 12'b011111110011;
   15212: result <= 12'b011111110011;
   15213: result <= 12'b011111110011;
   15214: result <= 12'b011111110011;
   15215: result <= 12'b011111110011;
   15216: result <= 12'b011111110011;
   15217: result <= 12'b011111110011;
   15218: result <= 12'b011111110011;
   15219: result <= 12'b011111110011;
   15220: result <= 12'b011111110011;
   15221: result <= 12'b011111110011;
   15222: result <= 12'b011111110011;
   15223: result <= 12'b011111110011;
   15224: result <= 12'b011111110011;
   15225: result <= 12'b011111110011;
   15226: result <= 12'b011111110011;
   15227: result <= 12'b011111110011;
   15228: result <= 12'b011111110011;
   15229: result <= 12'b011111110011;
   15230: result <= 12'b011111110011;
   15231: result <= 12'b011111110011;
   15232: result <= 12'b011111110011;
   15233: result <= 12'b011111110011;
   15234: result <= 12'b011111110011;
   15235: result <= 12'b011111110011;
   15236: result <= 12'b011111110011;
   15237: result <= 12'b011111110011;
   15238: result <= 12'b011111110011;
   15239: result <= 12'b011111110011;
   15240: result <= 12'b011111110011;
   15241: result <= 12'b011111110011;
   15242: result <= 12'b011111110011;
   15243: result <= 12'b011111110011;
   15244: result <= 12'b011111110011;
   15245: result <= 12'b011111110011;
   15246: result <= 12'b011111110011;
   15247: result <= 12'b011111110011;
   15248: result <= 12'b011111110011;
   15249: result <= 12'b011111110011;
   15250: result <= 12'b011111110011;
   15251: result <= 12'b011111110011;
   15252: result <= 12'b011111110011;
   15253: result <= 12'b011111110011;
   15254: result <= 12'b011111110011;
   15255: result <= 12'b011111110100;
   15256: result <= 12'b011111110100;
   15257: result <= 12'b011111110100;
   15258: result <= 12'b011111110100;
   15259: result <= 12'b011111110100;
   15260: result <= 12'b011111110100;
   15261: result <= 12'b011111110100;
   15262: result <= 12'b011111110100;
   15263: result <= 12'b011111110100;
   15264: result <= 12'b011111110100;
   15265: result <= 12'b011111110100;
   15266: result <= 12'b011111110100;
   15267: result <= 12'b011111110100;
   15268: result <= 12'b011111110100;
   15269: result <= 12'b011111110100;
   15270: result <= 12'b011111110100;
   15271: result <= 12'b011111110100;
   15272: result <= 12'b011111110100;
   15273: result <= 12'b011111110100;
   15274: result <= 12'b011111110100;
   15275: result <= 12'b011111110100;
   15276: result <= 12'b011111110100;
   15277: result <= 12'b011111110100;
   15278: result <= 12'b011111110100;
   15279: result <= 12'b011111110100;
   15280: result <= 12'b011111110100;
   15281: result <= 12'b011111110100;
   15282: result <= 12'b011111110100;
   15283: result <= 12'b011111110100;
   15284: result <= 12'b011111110100;
   15285: result <= 12'b011111110100;
   15286: result <= 12'b011111110100;
   15287: result <= 12'b011111110100;
   15288: result <= 12'b011111110100;
   15289: result <= 12'b011111110100;
   15290: result <= 12'b011111110100;
   15291: result <= 12'b011111110100;
   15292: result <= 12'b011111110100;
   15293: result <= 12'b011111110100;
   15294: result <= 12'b011111110100;
   15295: result <= 12'b011111110100;
   15296: result <= 12'b011111110100;
   15297: result <= 12'b011111110100;
   15298: result <= 12'b011111110100;
   15299: result <= 12'b011111110100;
   15300: result <= 12'b011111110100;
   15301: result <= 12'b011111110100;
   15302: result <= 12'b011111110100;
   15303: result <= 12'b011111110101;
   15304: result <= 12'b011111110101;
   15305: result <= 12'b011111110101;
   15306: result <= 12'b011111110101;
   15307: result <= 12'b011111110101;
   15308: result <= 12'b011111110101;
   15309: result <= 12'b011111110101;
   15310: result <= 12'b011111110101;
   15311: result <= 12'b011111110101;
   15312: result <= 12'b011111110101;
   15313: result <= 12'b011111110101;
   15314: result <= 12'b011111110101;
   15315: result <= 12'b011111110101;
   15316: result <= 12'b011111110101;
   15317: result <= 12'b011111110101;
   15318: result <= 12'b011111110101;
   15319: result <= 12'b011111110101;
   15320: result <= 12'b011111110101;
   15321: result <= 12'b011111110101;
   15322: result <= 12'b011111110101;
   15323: result <= 12'b011111110101;
   15324: result <= 12'b011111110101;
   15325: result <= 12'b011111110101;
   15326: result <= 12'b011111110101;
   15327: result <= 12'b011111110101;
   15328: result <= 12'b011111110101;
   15329: result <= 12'b011111110101;
   15330: result <= 12'b011111110101;
   15331: result <= 12'b011111110101;
   15332: result <= 12'b011111110101;
   15333: result <= 12'b011111110101;
   15334: result <= 12'b011111110101;
   15335: result <= 12'b011111110101;
   15336: result <= 12'b011111110101;
   15337: result <= 12'b011111110101;
   15338: result <= 12'b011111110101;
   15339: result <= 12'b011111110101;
   15340: result <= 12'b011111110101;
   15341: result <= 12'b011111110101;
   15342: result <= 12'b011111110101;
   15343: result <= 12'b011111110101;
   15344: result <= 12'b011111110101;
   15345: result <= 12'b011111110101;
   15346: result <= 12'b011111110101;
   15347: result <= 12'b011111110101;
   15348: result <= 12'b011111110101;
   15349: result <= 12'b011111110101;
   15350: result <= 12'b011111110101;
   15351: result <= 12'b011111110101;
   15352: result <= 12'b011111110101;
   15353: result <= 12'b011111110110;
   15354: result <= 12'b011111110110;
   15355: result <= 12'b011111110110;
   15356: result <= 12'b011111110110;
   15357: result <= 12'b011111110110;
   15358: result <= 12'b011111110110;
   15359: result <= 12'b011111110110;
   15360: result <= 12'b011111110110;
   15361: result <= 12'b011111110110;
   15362: result <= 12'b011111110110;
   15363: result <= 12'b011111110110;
   15364: result <= 12'b011111110110;
   15365: result <= 12'b011111110110;
   15366: result <= 12'b011111110110;
   15367: result <= 12'b011111110110;
   15368: result <= 12'b011111110110;
   15369: result <= 12'b011111110110;
   15370: result <= 12'b011111110110;
   15371: result <= 12'b011111110110;
   15372: result <= 12'b011111110110;
   15373: result <= 12'b011111110110;
   15374: result <= 12'b011111110110;
   15375: result <= 12'b011111110110;
   15376: result <= 12'b011111110110;
   15377: result <= 12'b011111110110;
   15378: result <= 12'b011111110110;
   15379: result <= 12'b011111110110;
   15380: result <= 12'b011111110110;
   15381: result <= 12'b011111110110;
   15382: result <= 12'b011111110110;
   15383: result <= 12'b011111110110;
   15384: result <= 12'b011111110110;
   15385: result <= 12'b011111110110;
   15386: result <= 12'b011111110110;
   15387: result <= 12'b011111110110;
   15388: result <= 12'b011111110110;
   15389: result <= 12'b011111110110;
   15390: result <= 12'b011111110110;
   15391: result <= 12'b011111110110;
   15392: result <= 12'b011111110110;
   15393: result <= 12'b011111110110;
   15394: result <= 12'b011111110110;
   15395: result <= 12'b011111110110;
   15396: result <= 12'b011111110110;
   15397: result <= 12'b011111110110;
   15398: result <= 12'b011111110110;
   15399: result <= 12'b011111110110;
   15400: result <= 12'b011111110110;
   15401: result <= 12'b011111110110;
   15402: result <= 12'b011111110110;
   15403: result <= 12'b011111110110;
   15404: result <= 12'b011111110110;
   15405: result <= 12'b011111110110;
   15406: result <= 12'b011111110111;
   15407: result <= 12'b011111110111;
   15408: result <= 12'b011111110111;
   15409: result <= 12'b011111110111;
   15410: result <= 12'b011111110111;
   15411: result <= 12'b011111110111;
   15412: result <= 12'b011111110111;
   15413: result <= 12'b011111110111;
   15414: result <= 12'b011111110111;
   15415: result <= 12'b011111110111;
   15416: result <= 12'b011111110111;
   15417: result <= 12'b011111110111;
   15418: result <= 12'b011111110111;
   15419: result <= 12'b011111110111;
   15420: result <= 12'b011111110111;
   15421: result <= 12'b011111110111;
   15422: result <= 12'b011111110111;
   15423: result <= 12'b011111110111;
   15424: result <= 12'b011111110111;
   15425: result <= 12'b011111110111;
   15426: result <= 12'b011111110111;
   15427: result <= 12'b011111110111;
   15428: result <= 12'b011111110111;
   15429: result <= 12'b011111110111;
   15430: result <= 12'b011111110111;
   15431: result <= 12'b011111110111;
   15432: result <= 12'b011111110111;
   15433: result <= 12'b011111110111;
   15434: result <= 12'b011111110111;
   15435: result <= 12'b011111110111;
   15436: result <= 12'b011111110111;
   15437: result <= 12'b011111110111;
   15438: result <= 12'b011111110111;
   15439: result <= 12'b011111110111;
   15440: result <= 12'b011111110111;
   15441: result <= 12'b011111110111;
   15442: result <= 12'b011111110111;
   15443: result <= 12'b011111110111;
   15444: result <= 12'b011111110111;
   15445: result <= 12'b011111110111;
   15446: result <= 12'b011111110111;
   15447: result <= 12'b011111110111;
   15448: result <= 12'b011111110111;
   15449: result <= 12'b011111110111;
   15450: result <= 12'b011111110111;
   15451: result <= 12'b011111110111;
   15452: result <= 12'b011111110111;
   15453: result <= 12'b011111110111;
   15454: result <= 12'b011111110111;
   15455: result <= 12'b011111110111;
   15456: result <= 12'b011111110111;
   15457: result <= 12'b011111110111;
   15458: result <= 12'b011111110111;
   15459: result <= 12'b011111110111;
   15460: result <= 12'b011111110111;
   15461: result <= 12'b011111110111;
   15462: result <= 12'b011111111000;
   15463: result <= 12'b011111111000;
   15464: result <= 12'b011111111000;
   15465: result <= 12'b011111111000;
   15466: result <= 12'b011111111000;
   15467: result <= 12'b011111111000;
   15468: result <= 12'b011111111000;
   15469: result <= 12'b011111111000;
   15470: result <= 12'b011111111000;
   15471: result <= 12'b011111111000;
   15472: result <= 12'b011111111000;
   15473: result <= 12'b011111111000;
   15474: result <= 12'b011111111000;
   15475: result <= 12'b011111111000;
   15476: result <= 12'b011111111000;
   15477: result <= 12'b011111111000;
   15478: result <= 12'b011111111000;
   15479: result <= 12'b011111111000;
   15480: result <= 12'b011111111000;
   15481: result <= 12'b011111111000;
   15482: result <= 12'b011111111000;
   15483: result <= 12'b011111111000;
   15484: result <= 12'b011111111000;
   15485: result <= 12'b011111111000;
   15486: result <= 12'b011111111000;
   15487: result <= 12'b011111111000;
   15488: result <= 12'b011111111000;
   15489: result <= 12'b011111111000;
   15490: result <= 12'b011111111000;
   15491: result <= 12'b011111111000;
   15492: result <= 12'b011111111000;
   15493: result <= 12'b011111111000;
   15494: result <= 12'b011111111000;
   15495: result <= 12'b011111111000;
   15496: result <= 12'b011111111000;
   15497: result <= 12'b011111111000;
   15498: result <= 12'b011111111000;
   15499: result <= 12'b011111111000;
   15500: result <= 12'b011111111000;
   15501: result <= 12'b011111111000;
   15502: result <= 12'b011111111000;
   15503: result <= 12'b011111111000;
   15504: result <= 12'b011111111000;
   15505: result <= 12'b011111111000;
   15506: result <= 12'b011111111000;
   15507: result <= 12'b011111111000;
   15508: result <= 12'b011111111000;
   15509: result <= 12'b011111111000;
   15510: result <= 12'b011111111000;
   15511: result <= 12'b011111111000;
   15512: result <= 12'b011111111000;
   15513: result <= 12'b011111111000;
   15514: result <= 12'b011111111000;
   15515: result <= 12'b011111111000;
   15516: result <= 12'b011111111000;
   15517: result <= 12'b011111111000;
   15518: result <= 12'b011111111000;
   15519: result <= 12'b011111111000;
   15520: result <= 12'b011111111000;
   15521: result <= 12'b011111111000;
   15522: result <= 12'b011111111001;
   15523: result <= 12'b011111111001;
   15524: result <= 12'b011111111001;
   15525: result <= 12'b011111111001;
   15526: result <= 12'b011111111001;
   15527: result <= 12'b011111111001;
   15528: result <= 12'b011111111001;
   15529: result <= 12'b011111111001;
   15530: result <= 12'b011111111001;
   15531: result <= 12'b011111111001;
   15532: result <= 12'b011111111001;
   15533: result <= 12'b011111111001;
   15534: result <= 12'b011111111001;
   15535: result <= 12'b011111111001;
   15536: result <= 12'b011111111001;
   15537: result <= 12'b011111111001;
   15538: result <= 12'b011111111001;
   15539: result <= 12'b011111111001;
   15540: result <= 12'b011111111001;
   15541: result <= 12'b011111111001;
   15542: result <= 12'b011111111001;
   15543: result <= 12'b011111111001;
   15544: result <= 12'b011111111001;
   15545: result <= 12'b011111111001;
   15546: result <= 12'b011111111001;
   15547: result <= 12'b011111111001;
   15548: result <= 12'b011111111001;
   15549: result <= 12'b011111111001;
   15550: result <= 12'b011111111001;
   15551: result <= 12'b011111111001;
   15552: result <= 12'b011111111001;
   15553: result <= 12'b011111111001;
   15554: result <= 12'b011111111001;
   15555: result <= 12'b011111111001;
   15556: result <= 12'b011111111001;
   15557: result <= 12'b011111111001;
   15558: result <= 12'b011111111001;
   15559: result <= 12'b011111111001;
   15560: result <= 12'b011111111001;
   15561: result <= 12'b011111111001;
   15562: result <= 12'b011111111001;
   15563: result <= 12'b011111111001;
   15564: result <= 12'b011111111001;
   15565: result <= 12'b011111111001;
   15566: result <= 12'b011111111001;
   15567: result <= 12'b011111111001;
   15568: result <= 12'b011111111001;
   15569: result <= 12'b011111111001;
   15570: result <= 12'b011111111001;
   15571: result <= 12'b011111111001;
   15572: result <= 12'b011111111001;
   15573: result <= 12'b011111111001;
   15574: result <= 12'b011111111001;
   15575: result <= 12'b011111111001;
   15576: result <= 12'b011111111001;
   15577: result <= 12'b011111111001;
   15578: result <= 12'b011111111001;
   15579: result <= 12'b011111111001;
   15580: result <= 12'b011111111001;
   15581: result <= 12'b011111111001;
   15582: result <= 12'b011111111001;
   15583: result <= 12'b011111111001;
   15584: result <= 12'b011111111001;
   15585: result <= 12'b011111111001;
   15586: result <= 12'b011111111010;
   15587: result <= 12'b011111111010;
   15588: result <= 12'b011111111010;
   15589: result <= 12'b011111111010;
   15590: result <= 12'b011111111010;
   15591: result <= 12'b011111111010;
   15592: result <= 12'b011111111010;
   15593: result <= 12'b011111111010;
   15594: result <= 12'b011111111010;
   15595: result <= 12'b011111111010;
   15596: result <= 12'b011111111010;
   15597: result <= 12'b011111111010;
   15598: result <= 12'b011111111010;
   15599: result <= 12'b011111111010;
   15600: result <= 12'b011111111010;
   15601: result <= 12'b011111111010;
   15602: result <= 12'b011111111010;
   15603: result <= 12'b011111111010;
   15604: result <= 12'b011111111010;
   15605: result <= 12'b011111111010;
   15606: result <= 12'b011111111010;
   15607: result <= 12'b011111111010;
   15608: result <= 12'b011111111010;
   15609: result <= 12'b011111111010;
   15610: result <= 12'b011111111010;
   15611: result <= 12'b011111111010;
   15612: result <= 12'b011111111010;
   15613: result <= 12'b011111111010;
   15614: result <= 12'b011111111010;
   15615: result <= 12'b011111111010;
   15616: result <= 12'b011111111010;
   15617: result <= 12'b011111111010;
   15618: result <= 12'b011111111010;
   15619: result <= 12'b011111111010;
   15620: result <= 12'b011111111010;
   15621: result <= 12'b011111111010;
   15622: result <= 12'b011111111010;
   15623: result <= 12'b011111111010;
   15624: result <= 12'b011111111010;
   15625: result <= 12'b011111111010;
   15626: result <= 12'b011111111010;
   15627: result <= 12'b011111111010;
   15628: result <= 12'b011111111010;
   15629: result <= 12'b011111111010;
   15630: result <= 12'b011111111010;
   15631: result <= 12'b011111111010;
   15632: result <= 12'b011111111010;
   15633: result <= 12'b011111111010;
   15634: result <= 12'b011111111010;
   15635: result <= 12'b011111111010;
   15636: result <= 12'b011111111010;
   15637: result <= 12'b011111111010;
   15638: result <= 12'b011111111010;
   15639: result <= 12'b011111111010;
   15640: result <= 12'b011111111010;
   15641: result <= 12'b011111111010;
   15642: result <= 12'b011111111010;
   15643: result <= 12'b011111111010;
   15644: result <= 12'b011111111010;
   15645: result <= 12'b011111111010;
   15646: result <= 12'b011111111010;
   15647: result <= 12'b011111111010;
   15648: result <= 12'b011111111010;
   15649: result <= 12'b011111111010;
   15650: result <= 12'b011111111010;
   15651: result <= 12'b011111111010;
   15652: result <= 12'b011111111010;
   15653: result <= 12'b011111111010;
   15654: result <= 12'b011111111010;
   15655: result <= 12'b011111111010;
   15656: result <= 12'b011111111011;
   15657: result <= 12'b011111111011;
   15658: result <= 12'b011111111011;
   15659: result <= 12'b011111111011;
   15660: result <= 12'b011111111011;
   15661: result <= 12'b011111111011;
   15662: result <= 12'b011111111011;
   15663: result <= 12'b011111111011;
   15664: result <= 12'b011111111011;
   15665: result <= 12'b011111111011;
   15666: result <= 12'b011111111011;
   15667: result <= 12'b011111111011;
   15668: result <= 12'b011111111011;
   15669: result <= 12'b011111111011;
   15670: result <= 12'b011111111011;
   15671: result <= 12'b011111111011;
   15672: result <= 12'b011111111011;
   15673: result <= 12'b011111111011;
   15674: result <= 12'b011111111011;
   15675: result <= 12'b011111111011;
   15676: result <= 12'b011111111011;
   15677: result <= 12'b011111111011;
   15678: result <= 12'b011111111011;
   15679: result <= 12'b011111111011;
   15680: result <= 12'b011111111011;
   15681: result <= 12'b011111111011;
   15682: result <= 12'b011111111011;
   15683: result <= 12'b011111111011;
   15684: result <= 12'b011111111011;
   15685: result <= 12'b011111111011;
   15686: result <= 12'b011111111011;
   15687: result <= 12'b011111111011;
   15688: result <= 12'b011111111011;
   15689: result <= 12'b011111111011;
   15690: result <= 12'b011111111011;
   15691: result <= 12'b011111111011;
   15692: result <= 12'b011111111011;
   15693: result <= 12'b011111111011;
   15694: result <= 12'b011111111011;
   15695: result <= 12'b011111111011;
   15696: result <= 12'b011111111011;
   15697: result <= 12'b011111111011;
   15698: result <= 12'b011111111011;
   15699: result <= 12'b011111111011;
   15700: result <= 12'b011111111011;
   15701: result <= 12'b011111111011;
   15702: result <= 12'b011111111011;
   15703: result <= 12'b011111111011;
   15704: result <= 12'b011111111011;
   15705: result <= 12'b011111111011;
   15706: result <= 12'b011111111011;
   15707: result <= 12'b011111111011;
   15708: result <= 12'b011111111011;
   15709: result <= 12'b011111111011;
   15710: result <= 12'b011111111011;
   15711: result <= 12'b011111111011;
   15712: result <= 12'b011111111011;
   15713: result <= 12'b011111111011;
   15714: result <= 12'b011111111011;
   15715: result <= 12'b011111111011;
   15716: result <= 12'b011111111011;
   15717: result <= 12'b011111111011;
   15718: result <= 12'b011111111011;
   15719: result <= 12'b011111111011;
   15720: result <= 12'b011111111011;
   15721: result <= 12'b011111111011;
   15722: result <= 12'b011111111011;
   15723: result <= 12'b011111111011;
   15724: result <= 12'b011111111011;
   15725: result <= 12'b011111111011;
   15726: result <= 12'b011111111011;
   15727: result <= 12'b011111111011;
   15728: result <= 12'b011111111011;
   15729: result <= 12'b011111111011;
   15730: result <= 12'b011111111011;
   15731: result <= 12'b011111111011;
   15732: result <= 12'b011111111100;
   15733: result <= 12'b011111111100;
   15734: result <= 12'b011111111100;
   15735: result <= 12'b011111111100;
   15736: result <= 12'b011111111100;
   15737: result <= 12'b011111111100;
   15738: result <= 12'b011111111100;
   15739: result <= 12'b011111111100;
   15740: result <= 12'b011111111100;
   15741: result <= 12'b011111111100;
   15742: result <= 12'b011111111100;
   15743: result <= 12'b011111111100;
   15744: result <= 12'b011111111100;
   15745: result <= 12'b011111111100;
   15746: result <= 12'b011111111100;
   15747: result <= 12'b011111111100;
   15748: result <= 12'b011111111100;
   15749: result <= 12'b011111111100;
   15750: result <= 12'b011111111100;
   15751: result <= 12'b011111111100;
   15752: result <= 12'b011111111100;
   15753: result <= 12'b011111111100;
   15754: result <= 12'b011111111100;
   15755: result <= 12'b011111111100;
   15756: result <= 12'b011111111100;
   15757: result <= 12'b011111111100;
   15758: result <= 12'b011111111100;
   15759: result <= 12'b011111111100;
   15760: result <= 12'b011111111100;
   15761: result <= 12'b011111111100;
   15762: result <= 12'b011111111100;
   15763: result <= 12'b011111111100;
   15764: result <= 12'b011111111100;
   15765: result <= 12'b011111111100;
   15766: result <= 12'b011111111100;
   15767: result <= 12'b011111111100;
   15768: result <= 12'b011111111100;
   15769: result <= 12'b011111111100;
   15770: result <= 12'b011111111100;
   15771: result <= 12'b011111111100;
   15772: result <= 12'b011111111100;
   15773: result <= 12'b011111111100;
   15774: result <= 12'b011111111100;
   15775: result <= 12'b011111111100;
   15776: result <= 12'b011111111100;
   15777: result <= 12'b011111111100;
   15778: result <= 12'b011111111100;
   15779: result <= 12'b011111111100;
   15780: result <= 12'b011111111100;
   15781: result <= 12'b011111111100;
   15782: result <= 12'b011111111100;
   15783: result <= 12'b011111111100;
   15784: result <= 12'b011111111100;
   15785: result <= 12'b011111111100;
   15786: result <= 12'b011111111100;
   15787: result <= 12'b011111111100;
   15788: result <= 12'b011111111100;
   15789: result <= 12'b011111111100;
   15790: result <= 12'b011111111100;
   15791: result <= 12'b011111111100;
   15792: result <= 12'b011111111100;
   15793: result <= 12'b011111111100;
   15794: result <= 12'b011111111100;
   15795: result <= 12'b011111111100;
   15796: result <= 12'b011111111100;
   15797: result <= 12'b011111111100;
   15798: result <= 12'b011111111100;
   15799: result <= 12'b011111111100;
   15800: result <= 12'b011111111100;
   15801: result <= 12'b011111111100;
   15802: result <= 12'b011111111100;
   15803: result <= 12'b011111111100;
   15804: result <= 12'b011111111100;
   15805: result <= 12'b011111111100;
   15806: result <= 12'b011111111100;
   15807: result <= 12'b011111111100;
   15808: result <= 12'b011111111100;
   15809: result <= 12'b011111111100;
   15810: result <= 12'b011111111100;
   15811: result <= 12'b011111111100;
   15812: result <= 12'b011111111100;
   15813: result <= 12'b011111111100;
   15814: result <= 12'b011111111100;
   15815: result <= 12'b011111111100;
   15816: result <= 12'b011111111100;
   15817: result <= 12'b011111111100;
   15818: result <= 12'b011111111100;
   15819: result <= 12'b011111111100;
   15820: result <= 12'b011111111101;
   15821: result <= 12'b011111111101;
   15822: result <= 12'b011111111101;
   15823: result <= 12'b011111111101;
   15824: result <= 12'b011111111101;
   15825: result <= 12'b011111111101;
   15826: result <= 12'b011111111101;
   15827: result <= 12'b011111111101;
   15828: result <= 12'b011111111101;
   15829: result <= 12'b011111111101;
   15830: result <= 12'b011111111101;
   15831: result <= 12'b011111111101;
   15832: result <= 12'b011111111101;
   15833: result <= 12'b011111111101;
   15834: result <= 12'b011111111101;
   15835: result <= 12'b011111111101;
   15836: result <= 12'b011111111101;
   15837: result <= 12'b011111111101;
   15838: result <= 12'b011111111101;
   15839: result <= 12'b011111111101;
   15840: result <= 12'b011111111101;
   15841: result <= 12'b011111111101;
   15842: result <= 12'b011111111101;
   15843: result <= 12'b011111111101;
   15844: result <= 12'b011111111101;
   15845: result <= 12'b011111111101;
   15846: result <= 12'b011111111101;
   15847: result <= 12'b011111111101;
   15848: result <= 12'b011111111101;
   15849: result <= 12'b011111111101;
   15850: result <= 12'b011111111101;
   15851: result <= 12'b011111111101;
   15852: result <= 12'b011111111101;
   15853: result <= 12'b011111111101;
   15854: result <= 12'b011111111101;
   15855: result <= 12'b011111111101;
   15856: result <= 12'b011111111101;
   15857: result <= 12'b011111111101;
   15858: result <= 12'b011111111101;
   15859: result <= 12'b011111111101;
   15860: result <= 12'b011111111101;
   15861: result <= 12'b011111111101;
   15862: result <= 12'b011111111101;
   15863: result <= 12'b011111111101;
   15864: result <= 12'b011111111101;
   15865: result <= 12'b011111111101;
   15866: result <= 12'b011111111101;
   15867: result <= 12'b011111111101;
   15868: result <= 12'b011111111101;
   15869: result <= 12'b011111111101;
   15870: result <= 12'b011111111101;
   15871: result <= 12'b011111111101;
   15872: result <= 12'b011111111101;
   15873: result <= 12'b011111111101;
   15874: result <= 12'b011111111101;
   15875: result <= 12'b011111111101;
   15876: result <= 12'b011111111101;
   15877: result <= 12'b011111111101;
   15878: result <= 12'b011111111101;
   15879: result <= 12'b011111111101;
   15880: result <= 12'b011111111101;
   15881: result <= 12'b011111111101;
   15882: result <= 12'b011111111101;
   15883: result <= 12'b011111111101;
   15884: result <= 12'b011111111101;
   15885: result <= 12'b011111111101;
   15886: result <= 12'b011111111101;
   15887: result <= 12'b011111111101;
   15888: result <= 12'b011111111101;
   15889: result <= 12'b011111111101;
   15890: result <= 12'b011111111101;
   15891: result <= 12'b011111111101;
   15892: result <= 12'b011111111101;
   15893: result <= 12'b011111111101;
   15894: result <= 12'b011111111101;
   15895: result <= 12'b011111111101;
   15896: result <= 12'b011111111101;
   15897: result <= 12'b011111111101;
   15898: result <= 12'b011111111101;
   15899: result <= 12'b011111111101;
   15900: result <= 12'b011111111101;
   15901: result <= 12'b011111111101;
   15902: result <= 12'b011111111101;
   15903: result <= 12'b011111111101;
   15904: result <= 12'b011111111101;
   15905: result <= 12'b011111111101;
   15906: result <= 12'b011111111101;
   15907: result <= 12'b011111111101;
   15908: result <= 12'b011111111101;
   15909: result <= 12'b011111111101;
   15910: result <= 12'b011111111101;
   15911: result <= 12'b011111111101;
   15912: result <= 12'b011111111101;
   15913: result <= 12'b011111111101;
   15914: result <= 12'b011111111101;
   15915: result <= 12'b011111111101;
   15916: result <= 12'b011111111101;
   15917: result <= 12'b011111111101;
   15918: result <= 12'b011111111101;
   15919: result <= 12'b011111111101;
   15920: result <= 12'b011111111101;
   15921: result <= 12'b011111111101;
   15922: result <= 12'b011111111101;
   15923: result <= 12'b011111111101;
   15924: result <= 12'b011111111110;
   15925: result <= 12'b011111111110;
   15926: result <= 12'b011111111110;
   15927: result <= 12'b011111111110;
   15928: result <= 12'b011111111110;
   15929: result <= 12'b011111111110;
   15930: result <= 12'b011111111110;
   15931: result <= 12'b011111111110;
   15932: result <= 12'b011111111110;
   15933: result <= 12'b011111111110;
   15934: result <= 12'b011111111110;
   15935: result <= 12'b011111111110;
   15936: result <= 12'b011111111110;
   15937: result <= 12'b011111111110;
   15938: result <= 12'b011111111110;
   15939: result <= 12'b011111111110;
   15940: result <= 12'b011111111110;
   15941: result <= 12'b011111111110;
   15942: result <= 12'b011111111110;
   15943: result <= 12'b011111111110;
   15944: result <= 12'b011111111110;
   15945: result <= 12'b011111111110;
   15946: result <= 12'b011111111110;
   15947: result <= 12'b011111111110;
   15948: result <= 12'b011111111110;
   15949: result <= 12'b011111111110;
   15950: result <= 12'b011111111110;
   15951: result <= 12'b011111111110;
   15952: result <= 12'b011111111110;
   15953: result <= 12'b011111111110;
   15954: result <= 12'b011111111110;
   15955: result <= 12'b011111111110;
   15956: result <= 12'b011111111110;
   15957: result <= 12'b011111111110;
   15958: result <= 12'b011111111110;
   15959: result <= 12'b011111111110;
   15960: result <= 12'b011111111110;
   15961: result <= 12'b011111111110;
   15962: result <= 12'b011111111110;
   15963: result <= 12'b011111111110;
   15964: result <= 12'b011111111110;
   15965: result <= 12'b011111111110;
   15966: result <= 12'b011111111110;
   15967: result <= 12'b011111111110;
   15968: result <= 12'b011111111110;
   15969: result <= 12'b011111111110;
   15970: result <= 12'b011111111110;
   15971: result <= 12'b011111111110;
   15972: result <= 12'b011111111110;
   15973: result <= 12'b011111111110;
   15974: result <= 12'b011111111110;
   15975: result <= 12'b011111111110;
   15976: result <= 12'b011111111110;
   15977: result <= 12'b011111111110;
   15978: result <= 12'b011111111110;
   15979: result <= 12'b011111111110;
   15980: result <= 12'b011111111110;
   15981: result <= 12'b011111111110;
   15982: result <= 12'b011111111110;
   15983: result <= 12'b011111111110;
   15984: result <= 12'b011111111110;
   15985: result <= 12'b011111111110;
   15986: result <= 12'b011111111110;
   15987: result <= 12'b011111111110;
   15988: result <= 12'b011111111110;
   15989: result <= 12'b011111111110;
   15990: result <= 12'b011111111110;
   15991: result <= 12'b011111111110;
   15992: result <= 12'b011111111110;
   15993: result <= 12'b011111111110;
   15994: result <= 12'b011111111110;
   15995: result <= 12'b011111111110;
   15996: result <= 12'b011111111110;
   15997: result <= 12'b011111111110;
   15998: result <= 12'b011111111110;
   15999: result <= 12'b011111111110;
   16000: result <= 12'b011111111110;
   16001: result <= 12'b011111111110;
   16002: result <= 12'b011111111110;
   16003: result <= 12'b011111111110;
   16004: result <= 12'b011111111110;
   16005: result <= 12'b011111111110;
   16006: result <= 12'b011111111110;
   16007: result <= 12'b011111111110;
   16008: result <= 12'b011111111110;
   16009: result <= 12'b011111111110;
   16010: result <= 12'b011111111110;
   16011: result <= 12'b011111111110;
   16012: result <= 12'b011111111110;
   16013: result <= 12'b011111111110;
   16014: result <= 12'b011111111110;
   16015: result <= 12'b011111111110;
   16016: result <= 12'b011111111110;
   16017: result <= 12'b011111111110;
   16018: result <= 12'b011111111110;
   16019: result <= 12'b011111111110;
   16020: result <= 12'b011111111110;
   16021: result <= 12'b011111111110;
   16022: result <= 12'b011111111110;
   16023: result <= 12'b011111111110;
   16024: result <= 12'b011111111110;
   16025: result <= 12'b011111111110;
   16026: result <= 12'b011111111110;
   16027: result <= 12'b011111111110;
   16028: result <= 12'b011111111110;
   16029: result <= 12'b011111111110;
   16030: result <= 12'b011111111110;
   16031: result <= 12'b011111111110;
   16032: result <= 12'b011111111110;
   16033: result <= 12'b011111111110;
   16034: result <= 12'b011111111110;
   16035: result <= 12'b011111111110;
   16036: result <= 12'b011111111110;
   16037: result <= 12'b011111111110;
   16038: result <= 12'b011111111110;
   16039: result <= 12'b011111111110;
   16040: result <= 12'b011111111110;
   16041: result <= 12'b011111111110;
   16042: result <= 12'b011111111110;
   16043: result <= 12'b011111111110;
   16044: result <= 12'b011111111110;
   16045: result <= 12'b011111111110;
   16046: result <= 12'b011111111110;
   16047: result <= 12'b011111111110;
   16048: result <= 12'b011111111110;
   16049: result <= 12'b011111111110;
   16050: result <= 12'b011111111110;
   16051: result <= 12'b011111111110;
   16052: result <= 12'b011111111110;
   16053: result <= 12'b011111111110;
   16054: result <= 12'b011111111110;
   16055: result <= 12'b011111111110;
   16056: result <= 12'b011111111110;
   16057: result <= 12'b011111111110;
   16058: result <= 12'b011111111110;
   16059: result <= 12'b011111111111;
   16060: result <= 12'b011111111111;
   16061: result <= 12'b011111111111;
   16062: result <= 12'b011111111111;
   16063: result <= 12'b011111111111;
   16064: result <= 12'b011111111111;
   16065: result <= 12'b011111111111;
   16066: result <= 12'b011111111111;
   16067: result <= 12'b011111111111;
   16068: result <= 12'b011111111111;
   16069: result <= 12'b011111111111;
   16070: result <= 12'b011111111111;
   16071: result <= 12'b011111111111;
   16072: result <= 12'b011111111111;
   16073: result <= 12'b011111111111;
   16074: result <= 12'b011111111111;
   16075: result <= 12'b011111111111;
   16076: result <= 12'b011111111111;
   16077: result <= 12'b011111111111;
   16078: result <= 12'b011111111111;
   16079: result <= 12'b011111111111;
   16080: result <= 12'b011111111111;
   16081: result <= 12'b011111111111;
   16082: result <= 12'b011111111111;
   16083: result <= 12'b011111111111;
   16084: result <= 12'b011111111111;
   16085: result <= 12'b011111111111;
   16086: result <= 12'b011111111111;
   16087: result <= 12'b011111111111;
   16088: result <= 12'b011111111111;
   16089: result <= 12'b011111111111;
   16090: result <= 12'b011111111111;
   16091: result <= 12'b011111111111;
   16092: result <= 12'b011111111111;
   16093: result <= 12'b011111111111;
   16094: result <= 12'b011111111111;
   16095: result <= 12'b011111111111;
   16096: result <= 12'b011111111111;
   16097: result <= 12'b011111111111;
   16098: result <= 12'b011111111111;
   16099: result <= 12'b011111111111;
   16100: result <= 12'b011111111111;
   16101: result <= 12'b011111111111;
   16102: result <= 12'b011111111111;
   16103: result <= 12'b011111111111;
   16104: result <= 12'b011111111111;
   16105: result <= 12'b011111111111;
   16106: result <= 12'b011111111111;
   16107: result <= 12'b011111111111;
   16108: result <= 12'b011111111111;
   16109: result <= 12'b011111111111;
   16110: result <= 12'b011111111111;
   16111: result <= 12'b011111111111;
   16112: result <= 12'b011111111111;
   16113: result <= 12'b011111111111;
   16114: result <= 12'b011111111111;
   16115: result <= 12'b011111111111;
   16116: result <= 12'b011111111111;
   16117: result <= 12'b011111111111;
   16118: result <= 12'b011111111111;
   16119: result <= 12'b011111111111;
   16120: result <= 12'b011111111111;
   16121: result <= 12'b011111111111;
   16122: result <= 12'b011111111111;
   16123: result <= 12'b011111111111;
   16124: result <= 12'b011111111111;
   16125: result <= 12'b011111111111;
   16126: result <= 12'b011111111111;
   16127: result <= 12'b011111111111;
   16128: result <= 12'b011111111111;
   16129: result <= 12'b011111111111;
   16130: result <= 12'b011111111111;
   16131: result <= 12'b011111111111;
   16132: result <= 12'b011111111111;
   16133: result <= 12'b011111111111;
   16134: result <= 12'b011111111111;
   16135: result <= 12'b011111111111;
   16136: result <= 12'b011111111111;
   16137: result <= 12'b011111111111;
   16138: result <= 12'b011111111111;
   16139: result <= 12'b011111111111;
   16140: result <= 12'b011111111111;
   16141: result <= 12'b011111111111;
   16142: result <= 12'b011111111111;
   16143: result <= 12'b011111111111;
   16144: result <= 12'b011111111111;
   16145: result <= 12'b011111111111;
   16146: result <= 12'b011111111111;
   16147: result <= 12'b011111111111;
   16148: result <= 12'b011111111111;
   16149: result <= 12'b011111111111;
   16150: result <= 12'b011111111111;
   16151: result <= 12'b011111111111;
   16152: result <= 12'b011111111111;
   16153: result <= 12'b011111111111;
   16154: result <= 12'b011111111111;
   16155: result <= 12'b011111111111;
   16156: result <= 12'b011111111111;
   16157: result <= 12'b011111111111;
   16158: result <= 12'b011111111111;
   16159: result <= 12'b011111111111;
   16160: result <= 12'b011111111111;
   16161: result <= 12'b011111111111;
   16162: result <= 12'b011111111111;
   16163: result <= 12'b011111111111;
   16164: result <= 12'b011111111111;
   16165: result <= 12'b011111111111;
   16166: result <= 12'b011111111111;
   16167: result <= 12'b011111111111;
   16168: result <= 12'b011111111111;
   16169: result <= 12'b011111111111;
   16170: result <= 12'b011111111111;
   16171: result <= 12'b011111111111;
   16172: result <= 12'b011111111111;
   16173: result <= 12'b011111111111;
   16174: result <= 12'b011111111111;
   16175: result <= 12'b011111111111;
   16176: result <= 12'b011111111111;
   16177: result <= 12'b011111111111;
   16178: result <= 12'b011111111111;
   16179: result <= 12'b011111111111;
   16180: result <= 12'b011111111111;
   16181: result <= 12'b011111111111;
   16182: result <= 12'b011111111111;
   16183: result <= 12'b011111111111;
   16184: result <= 12'b011111111111;
   16185: result <= 12'b011111111111;
   16186: result <= 12'b011111111111;
   16187: result <= 12'b011111111111;
   16188: result <= 12'b011111111111;
   16189: result <= 12'b011111111111;
   16190: result <= 12'b011111111111;
   16191: result <= 12'b011111111111;
   16192: result <= 12'b011111111111;
   16193: result <= 12'b011111111111;
   16194: result <= 12'b011111111111;
   16195: result <= 12'b011111111111;
   16196: result <= 12'b011111111111;
   16197: result <= 12'b011111111111;
   16198: result <= 12'b011111111111;
   16199: result <= 12'b011111111111;
   16200: result <= 12'b011111111111;
   16201: result <= 12'b011111111111;
   16202: result <= 12'b011111111111;
   16203: result <= 12'b011111111111;
   16204: result <= 12'b011111111111;
   16205: result <= 12'b011111111111;
   16206: result <= 12'b011111111111;
   16207: result <= 12'b011111111111;
   16208: result <= 12'b011111111111;
   16209: result <= 12'b011111111111;
   16210: result <= 12'b011111111111;
   16211: result <= 12'b011111111111;
   16212: result <= 12'b011111111111;
   16213: result <= 12'b011111111111;
   16214: result <= 12'b011111111111;
   16215: result <= 12'b011111111111;
   16216: result <= 12'b011111111111;
   16217: result <= 12'b011111111111;
   16218: result <= 12'b011111111111;
   16219: result <= 12'b011111111111;
   16220: result <= 12'b011111111111;
   16221: result <= 12'b011111111111;
   16222: result <= 12'b011111111111;
   16223: result <= 12'b011111111111;
   16224: result <= 12'b011111111111;
   16225: result <= 12'b011111111111;
   16226: result <= 12'b011111111111;
   16227: result <= 12'b011111111111;
   16228: result <= 12'b011111111111;
   16229: result <= 12'b011111111111;
   16230: result <= 12'b011111111111;
   16231: result <= 12'b011111111111;
   16232: result <= 12'b011111111111;
   16233: result <= 12'b011111111111;
   16234: result <= 12'b011111111111;
   16235: result <= 12'b011111111111;
   16236: result <= 12'b011111111111;
   16237: result <= 12'b011111111111;
   16238: result <= 12'b011111111111;
   16239: result <= 12'b011111111111;
   16240: result <= 12'b011111111111;
   16241: result <= 12'b011111111111;
   16242: result <= 12'b011111111111;
   16243: result <= 12'b011111111111;
   16244: result <= 12'b011111111111;
   16245: result <= 12'b011111111111;
   16246: result <= 12'b011111111111;
   16247: result <= 12'b011111111111;
   16248: result <= 12'b011111111111;
   16249: result <= 12'b011111111111;
   16250: result <= 12'b011111111111;
   16251: result <= 12'b011111111111;
   16252: result <= 12'b011111111111;
   16253: result <= 12'b011111111111;
   16254: result <= 12'b011111111111;
   16255: result <= 12'b011111111111;
   16256: result <= 12'b011111111111;
   16257: result <= 12'b011111111111;
   16258: result <= 12'b011111111111;
   16259: result <= 12'b011111111111;
   16260: result <= 12'b011111111111;
   16261: result <= 12'b011111111111;
   16262: result <= 12'b011111111111;
   16263: result <= 12'b011111111111;
   16264: result <= 12'b011111111111;
   16265: result <= 12'b011111111111;
   16266: result <= 12'b011111111111;
   16267: result <= 12'b011111111111;
   16268: result <= 12'b011111111111;
   16269: result <= 12'b011111111111;
   16270: result <= 12'b011111111111;
   16271: result <= 12'b011111111111;
   16272: result <= 12'b011111111111;
   16273: result <= 12'b011111111111;
   16274: result <= 12'b011111111111;
   16275: result <= 12'b011111111111;
   16276: result <= 12'b011111111111;
   16277: result <= 12'b011111111111;
   16278: result <= 12'b011111111111;
   16279: result <= 12'b011111111111;
   16280: result <= 12'b011111111111;
   16281: result <= 12'b011111111111;
   16282: result <= 12'b011111111111;
   16283: result <= 12'b011111111111;
   16284: result <= 12'b011111111111;
   16285: result <= 12'b011111111111;
   16286: result <= 12'b011111111111;
   16287: result <= 12'b011111111111;
   16288: result <= 12'b011111111111;
   16289: result <= 12'b011111111111;
   16290: result <= 12'b011111111111;
   16291: result <= 12'b011111111111;
   16292: result <= 12'b011111111111;
   16293: result <= 12'b011111111111;
   16294: result <= 12'b011111111111;
   16295: result <= 12'b011111111111;
   16296: result <= 12'b011111111111;
   16297: result <= 12'b011111111111;
   16298: result <= 12'b011111111111;
   16299: result <= 12'b011111111111;
   16300: result <= 12'b011111111111;
   16301: result <= 12'b011111111111;
   16302: result <= 12'b011111111111;
   16303: result <= 12'b011111111111;
   16304: result <= 12'b011111111111;
   16305: result <= 12'b011111111111;
   16306: result <= 12'b011111111111;
   16307: result <= 12'b011111111111;
   16308: result <= 12'b011111111111;
   16309: result <= 12'b011111111111;
   16310: result <= 12'b011111111111;
   16311: result <= 12'b011111111111;
   16312: result <= 12'b011111111111;
   16313: result <= 12'b011111111111;
   16314: result <= 12'b011111111111;
   16315: result <= 12'b011111111111;
   16316: result <= 12'b011111111111;
   16317: result <= 12'b011111111111;
   16318: result <= 12'b011111111111;
   16319: result <= 12'b011111111111;
   16320: result <= 12'b011111111111;
   16321: result <= 12'b011111111111;
   16322: result <= 12'b011111111111;
   16323: result <= 12'b011111111111;
   16324: result <= 12'b011111111111;
   16325: result <= 12'b011111111111;
   16326: result <= 12'b011111111111;
   16327: result <= 12'b011111111111;
   16328: result <= 12'b011111111111;
   16329: result <= 12'b011111111111;
   16330: result <= 12'b011111111111;
   16331: result <= 12'b011111111111;
   16332: result <= 12'b011111111111;
   16333: result <= 12'b011111111111;
   16334: result <= 12'b011111111111;
   16335: result <= 12'b011111111111;
   16336: result <= 12'b011111111111;
   16337: result <= 12'b011111111111;
   16338: result <= 12'b011111111111;
   16339: result <= 12'b011111111111;
   16340: result <= 12'b011111111111;
   16341: result <= 12'b011111111111;
   16342: result <= 12'b011111111111;
   16343: result <= 12'b011111111111;
   16344: result <= 12'b011111111111;
   16345: result <= 12'b011111111111;
   16346: result <= 12'b011111111111;
   16347: result <= 12'b011111111111;
   16348: result <= 12'b011111111111;
   16349: result <= 12'b011111111111;
   16350: result <= 12'b011111111111;
   16351: result <= 12'b011111111111;
   16352: result <= 12'b011111111111;
   16353: result <= 12'b011111111111;
   16354: result <= 12'b011111111111;
   16355: result <= 12'b011111111111;
   16356: result <= 12'b011111111111;
   16357: result <= 12'b011111111111;
   16358: result <= 12'b011111111111;
   16359: result <= 12'b011111111111;
   16360: result <= 12'b011111111111;
   16361: result <= 12'b011111111111;
   16362: result <= 12'b011111111111;
   16363: result <= 12'b011111111111;
   16364: result <= 12'b011111111111;
   16365: result <= 12'b011111111111;
   16366: result <= 12'b011111111111;
   16367: result <= 12'b011111111111;
   16368: result <= 12'b011111111111;
   16369: result <= 12'b011111111111;
   16370: result <= 12'b011111111111;
   16371: result <= 12'b011111111111;
   16372: result <= 12'b011111111111;
   16373: result <= 12'b011111111111;
   16374: result <= 12'b011111111111;
   16375: result <= 12'b011111111111;
   16376: result <= 12'b011111111111;
   16377: result <= 12'b011111111111;
   16378: result <= 12'b011111111111;
   16379: result <= 12'b011111111111;
   16380: result <= 12'b011111111111;
   16381: result <= 12'b011111111111;
   16382: result <= 12'b011111111111;
   16383: result <= 12'b011111111111;
   16384: result <= 12'b100000000000;
   16385: result <= 12'b011111111111;
   16386: result <= 12'b011111111111;
   16387: result <= 12'b011111111111;
   16388: result <= 12'b011111111111;
   16389: result <= 12'b011111111111;
   16390: result <= 12'b011111111111;
   16391: result <= 12'b011111111111;
   16392: result <= 12'b011111111111;
   16393: result <= 12'b011111111111;
   16394: result <= 12'b011111111111;
   16395: result <= 12'b011111111111;
   16396: result <= 12'b011111111111;
   16397: result <= 12'b011111111111;
   16398: result <= 12'b011111111111;
   16399: result <= 12'b011111111111;
   16400: result <= 12'b011111111111;
   16401: result <= 12'b011111111111;
   16402: result <= 12'b011111111111;
   16403: result <= 12'b011111111111;
   16404: result <= 12'b011111111111;
   16405: result <= 12'b011111111111;
   16406: result <= 12'b011111111111;
   16407: result <= 12'b011111111111;
   16408: result <= 12'b011111111111;
   16409: result <= 12'b011111111111;
   16410: result <= 12'b011111111111;
   16411: result <= 12'b011111111111;
   16412: result <= 12'b011111111111;
   16413: result <= 12'b011111111111;
   16414: result <= 12'b011111111111;
   16415: result <= 12'b011111111111;
   16416: result <= 12'b011111111111;
   16417: result <= 12'b011111111111;
   16418: result <= 12'b011111111111;
   16419: result <= 12'b011111111111;
   16420: result <= 12'b011111111111;
   16421: result <= 12'b011111111111;
   16422: result <= 12'b011111111111;
   16423: result <= 12'b011111111111;
   16424: result <= 12'b011111111111;
   16425: result <= 12'b011111111111;
   16426: result <= 12'b011111111111;
   16427: result <= 12'b011111111111;
   16428: result <= 12'b011111111111;
   16429: result <= 12'b011111111111;
   16430: result <= 12'b011111111111;
   16431: result <= 12'b011111111111;
   16432: result <= 12'b011111111111;
   16433: result <= 12'b011111111111;
   16434: result <= 12'b011111111111;
   16435: result <= 12'b011111111111;
   16436: result <= 12'b011111111111;
   16437: result <= 12'b011111111111;
   16438: result <= 12'b011111111111;
   16439: result <= 12'b011111111111;
   16440: result <= 12'b011111111111;
   16441: result <= 12'b011111111111;
   16442: result <= 12'b011111111111;
   16443: result <= 12'b011111111111;
   16444: result <= 12'b011111111111;
   16445: result <= 12'b011111111111;
   16446: result <= 12'b011111111111;
   16447: result <= 12'b011111111111;
   16448: result <= 12'b011111111111;
   16449: result <= 12'b011111111111;
   16450: result <= 12'b011111111111;
   16451: result <= 12'b011111111111;
   16452: result <= 12'b011111111111;
   16453: result <= 12'b011111111111;
   16454: result <= 12'b011111111111;
   16455: result <= 12'b011111111111;
   16456: result <= 12'b011111111111;
   16457: result <= 12'b011111111111;
   16458: result <= 12'b011111111111;
   16459: result <= 12'b011111111111;
   16460: result <= 12'b011111111111;
   16461: result <= 12'b011111111111;
   16462: result <= 12'b011111111111;
   16463: result <= 12'b011111111111;
   16464: result <= 12'b011111111111;
   16465: result <= 12'b011111111111;
   16466: result <= 12'b011111111111;
   16467: result <= 12'b011111111111;
   16468: result <= 12'b011111111111;
   16469: result <= 12'b011111111111;
   16470: result <= 12'b011111111111;
   16471: result <= 12'b011111111111;
   16472: result <= 12'b011111111111;
   16473: result <= 12'b011111111111;
   16474: result <= 12'b011111111111;
   16475: result <= 12'b011111111111;
   16476: result <= 12'b011111111111;
   16477: result <= 12'b011111111111;
   16478: result <= 12'b011111111111;
   16479: result <= 12'b011111111111;
   16480: result <= 12'b011111111111;
   16481: result <= 12'b011111111111;
   16482: result <= 12'b011111111111;
   16483: result <= 12'b011111111111;
   16484: result <= 12'b011111111111;
   16485: result <= 12'b011111111111;
   16486: result <= 12'b011111111111;
   16487: result <= 12'b011111111111;
   16488: result <= 12'b011111111111;
   16489: result <= 12'b011111111111;
   16490: result <= 12'b011111111111;
   16491: result <= 12'b011111111111;
   16492: result <= 12'b011111111111;
   16493: result <= 12'b011111111111;
   16494: result <= 12'b011111111111;
   16495: result <= 12'b011111111111;
   16496: result <= 12'b011111111111;
   16497: result <= 12'b011111111111;
   16498: result <= 12'b011111111111;
   16499: result <= 12'b011111111111;
   16500: result <= 12'b011111111111;
   16501: result <= 12'b011111111111;
   16502: result <= 12'b011111111111;
   16503: result <= 12'b011111111111;
   16504: result <= 12'b011111111111;
   16505: result <= 12'b011111111111;
   16506: result <= 12'b011111111111;
   16507: result <= 12'b011111111111;
   16508: result <= 12'b011111111111;
   16509: result <= 12'b011111111111;
   16510: result <= 12'b011111111111;
   16511: result <= 12'b011111111111;
   16512: result <= 12'b011111111111;
   16513: result <= 12'b011111111111;
   16514: result <= 12'b011111111111;
   16515: result <= 12'b011111111111;
   16516: result <= 12'b011111111111;
   16517: result <= 12'b011111111111;
   16518: result <= 12'b011111111111;
   16519: result <= 12'b011111111111;
   16520: result <= 12'b011111111111;
   16521: result <= 12'b011111111111;
   16522: result <= 12'b011111111111;
   16523: result <= 12'b011111111111;
   16524: result <= 12'b011111111111;
   16525: result <= 12'b011111111111;
   16526: result <= 12'b011111111111;
   16527: result <= 12'b011111111111;
   16528: result <= 12'b011111111111;
   16529: result <= 12'b011111111111;
   16530: result <= 12'b011111111111;
   16531: result <= 12'b011111111111;
   16532: result <= 12'b011111111111;
   16533: result <= 12'b011111111111;
   16534: result <= 12'b011111111111;
   16535: result <= 12'b011111111111;
   16536: result <= 12'b011111111111;
   16537: result <= 12'b011111111111;
   16538: result <= 12'b011111111111;
   16539: result <= 12'b011111111111;
   16540: result <= 12'b011111111111;
   16541: result <= 12'b011111111111;
   16542: result <= 12'b011111111111;
   16543: result <= 12'b011111111111;
   16544: result <= 12'b011111111111;
   16545: result <= 12'b011111111111;
   16546: result <= 12'b011111111111;
   16547: result <= 12'b011111111111;
   16548: result <= 12'b011111111111;
   16549: result <= 12'b011111111111;
   16550: result <= 12'b011111111111;
   16551: result <= 12'b011111111111;
   16552: result <= 12'b011111111111;
   16553: result <= 12'b011111111111;
   16554: result <= 12'b011111111111;
   16555: result <= 12'b011111111111;
   16556: result <= 12'b011111111111;
   16557: result <= 12'b011111111111;
   16558: result <= 12'b011111111111;
   16559: result <= 12'b011111111111;
   16560: result <= 12'b011111111111;
   16561: result <= 12'b011111111111;
   16562: result <= 12'b011111111111;
   16563: result <= 12'b011111111111;
   16564: result <= 12'b011111111111;
   16565: result <= 12'b011111111111;
   16566: result <= 12'b011111111111;
   16567: result <= 12'b011111111111;
   16568: result <= 12'b011111111111;
   16569: result <= 12'b011111111111;
   16570: result <= 12'b011111111111;
   16571: result <= 12'b011111111111;
   16572: result <= 12'b011111111111;
   16573: result <= 12'b011111111111;
   16574: result <= 12'b011111111111;
   16575: result <= 12'b011111111111;
   16576: result <= 12'b011111111111;
   16577: result <= 12'b011111111111;
   16578: result <= 12'b011111111111;
   16579: result <= 12'b011111111111;
   16580: result <= 12'b011111111111;
   16581: result <= 12'b011111111111;
   16582: result <= 12'b011111111111;
   16583: result <= 12'b011111111111;
   16584: result <= 12'b011111111111;
   16585: result <= 12'b011111111111;
   16586: result <= 12'b011111111111;
   16587: result <= 12'b011111111111;
   16588: result <= 12'b011111111111;
   16589: result <= 12'b011111111111;
   16590: result <= 12'b011111111111;
   16591: result <= 12'b011111111111;
   16592: result <= 12'b011111111111;
   16593: result <= 12'b011111111111;
   16594: result <= 12'b011111111111;
   16595: result <= 12'b011111111111;
   16596: result <= 12'b011111111111;
   16597: result <= 12'b011111111111;
   16598: result <= 12'b011111111111;
   16599: result <= 12'b011111111111;
   16600: result <= 12'b011111111111;
   16601: result <= 12'b011111111111;
   16602: result <= 12'b011111111111;
   16603: result <= 12'b011111111111;
   16604: result <= 12'b011111111111;
   16605: result <= 12'b011111111111;
   16606: result <= 12'b011111111111;
   16607: result <= 12'b011111111111;
   16608: result <= 12'b011111111111;
   16609: result <= 12'b011111111111;
   16610: result <= 12'b011111111111;
   16611: result <= 12'b011111111111;
   16612: result <= 12'b011111111111;
   16613: result <= 12'b011111111111;
   16614: result <= 12'b011111111111;
   16615: result <= 12'b011111111111;
   16616: result <= 12'b011111111111;
   16617: result <= 12'b011111111111;
   16618: result <= 12'b011111111111;
   16619: result <= 12'b011111111111;
   16620: result <= 12'b011111111111;
   16621: result <= 12'b011111111111;
   16622: result <= 12'b011111111111;
   16623: result <= 12'b011111111111;
   16624: result <= 12'b011111111111;
   16625: result <= 12'b011111111111;
   16626: result <= 12'b011111111111;
   16627: result <= 12'b011111111111;
   16628: result <= 12'b011111111111;
   16629: result <= 12'b011111111111;
   16630: result <= 12'b011111111111;
   16631: result <= 12'b011111111111;
   16632: result <= 12'b011111111111;
   16633: result <= 12'b011111111111;
   16634: result <= 12'b011111111111;
   16635: result <= 12'b011111111111;
   16636: result <= 12'b011111111111;
   16637: result <= 12'b011111111111;
   16638: result <= 12'b011111111111;
   16639: result <= 12'b011111111111;
   16640: result <= 12'b011111111111;
   16641: result <= 12'b011111111111;
   16642: result <= 12'b011111111111;
   16643: result <= 12'b011111111111;
   16644: result <= 12'b011111111111;
   16645: result <= 12'b011111111111;
   16646: result <= 12'b011111111111;
   16647: result <= 12'b011111111111;
   16648: result <= 12'b011111111111;
   16649: result <= 12'b011111111111;
   16650: result <= 12'b011111111111;
   16651: result <= 12'b011111111111;
   16652: result <= 12'b011111111111;
   16653: result <= 12'b011111111111;
   16654: result <= 12'b011111111111;
   16655: result <= 12'b011111111111;
   16656: result <= 12'b011111111111;
   16657: result <= 12'b011111111111;
   16658: result <= 12'b011111111111;
   16659: result <= 12'b011111111111;
   16660: result <= 12'b011111111111;
   16661: result <= 12'b011111111111;
   16662: result <= 12'b011111111111;
   16663: result <= 12'b011111111111;
   16664: result <= 12'b011111111111;
   16665: result <= 12'b011111111111;
   16666: result <= 12'b011111111111;
   16667: result <= 12'b011111111111;
   16668: result <= 12'b011111111111;
   16669: result <= 12'b011111111111;
   16670: result <= 12'b011111111111;
   16671: result <= 12'b011111111111;
   16672: result <= 12'b011111111111;
   16673: result <= 12'b011111111111;
   16674: result <= 12'b011111111111;
   16675: result <= 12'b011111111111;
   16676: result <= 12'b011111111111;
   16677: result <= 12'b011111111111;
   16678: result <= 12'b011111111111;
   16679: result <= 12'b011111111111;
   16680: result <= 12'b011111111111;
   16681: result <= 12'b011111111111;
   16682: result <= 12'b011111111111;
   16683: result <= 12'b011111111111;
   16684: result <= 12'b011111111111;
   16685: result <= 12'b011111111111;
   16686: result <= 12'b011111111111;
   16687: result <= 12'b011111111111;
   16688: result <= 12'b011111111111;
   16689: result <= 12'b011111111111;
   16690: result <= 12'b011111111111;
   16691: result <= 12'b011111111111;
   16692: result <= 12'b011111111111;
   16693: result <= 12'b011111111111;
   16694: result <= 12'b011111111111;
   16695: result <= 12'b011111111111;
   16696: result <= 12'b011111111111;
   16697: result <= 12'b011111111111;
   16698: result <= 12'b011111111111;
   16699: result <= 12'b011111111111;
   16700: result <= 12'b011111111111;
   16701: result <= 12'b011111111111;
   16702: result <= 12'b011111111111;
   16703: result <= 12'b011111111111;
   16704: result <= 12'b011111111111;
   16705: result <= 12'b011111111111;
   16706: result <= 12'b011111111111;
   16707: result <= 12'b011111111111;
   16708: result <= 12'b011111111111;
   16709: result <= 12'b011111111111;
   16710: result <= 12'b011111111110;
   16711: result <= 12'b011111111110;
   16712: result <= 12'b011111111110;
   16713: result <= 12'b011111111110;
   16714: result <= 12'b011111111110;
   16715: result <= 12'b011111111110;
   16716: result <= 12'b011111111110;
   16717: result <= 12'b011111111110;
   16718: result <= 12'b011111111110;
   16719: result <= 12'b011111111110;
   16720: result <= 12'b011111111110;
   16721: result <= 12'b011111111110;
   16722: result <= 12'b011111111110;
   16723: result <= 12'b011111111110;
   16724: result <= 12'b011111111110;
   16725: result <= 12'b011111111110;
   16726: result <= 12'b011111111110;
   16727: result <= 12'b011111111110;
   16728: result <= 12'b011111111110;
   16729: result <= 12'b011111111110;
   16730: result <= 12'b011111111110;
   16731: result <= 12'b011111111110;
   16732: result <= 12'b011111111110;
   16733: result <= 12'b011111111110;
   16734: result <= 12'b011111111110;
   16735: result <= 12'b011111111110;
   16736: result <= 12'b011111111110;
   16737: result <= 12'b011111111110;
   16738: result <= 12'b011111111110;
   16739: result <= 12'b011111111110;
   16740: result <= 12'b011111111110;
   16741: result <= 12'b011111111110;
   16742: result <= 12'b011111111110;
   16743: result <= 12'b011111111110;
   16744: result <= 12'b011111111110;
   16745: result <= 12'b011111111110;
   16746: result <= 12'b011111111110;
   16747: result <= 12'b011111111110;
   16748: result <= 12'b011111111110;
   16749: result <= 12'b011111111110;
   16750: result <= 12'b011111111110;
   16751: result <= 12'b011111111110;
   16752: result <= 12'b011111111110;
   16753: result <= 12'b011111111110;
   16754: result <= 12'b011111111110;
   16755: result <= 12'b011111111110;
   16756: result <= 12'b011111111110;
   16757: result <= 12'b011111111110;
   16758: result <= 12'b011111111110;
   16759: result <= 12'b011111111110;
   16760: result <= 12'b011111111110;
   16761: result <= 12'b011111111110;
   16762: result <= 12'b011111111110;
   16763: result <= 12'b011111111110;
   16764: result <= 12'b011111111110;
   16765: result <= 12'b011111111110;
   16766: result <= 12'b011111111110;
   16767: result <= 12'b011111111110;
   16768: result <= 12'b011111111110;
   16769: result <= 12'b011111111110;
   16770: result <= 12'b011111111110;
   16771: result <= 12'b011111111110;
   16772: result <= 12'b011111111110;
   16773: result <= 12'b011111111110;
   16774: result <= 12'b011111111110;
   16775: result <= 12'b011111111110;
   16776: result <= 12'b011111111110;
   16777: result <= 12'b011111111110;
   16778: result <= 12'b011111111110;
   16779: result <= 12'b011111111110;
   16780: result <= 12'b011111111110;
   16781: result <= 12'b011111111110;
   16782: result <= 12'b011111111110;
   16783: result <= 12'b011111111110;
   16784: result <= 12'b011111111110;
   16785: result <= 12'b011111111110;
   16786: result <= 12'b011111111110;
   16787: result <= 12'b011111111110;
   16788: result <= 12'b011111111110;
   16789: result <= 12'b011111111110;
   16790: result <= 12'b011111111110;
   16791: result <= 12'b011111111110;
   16792: result <= 12'b011111111110;
   16793: result <= 12'b011111111110;
   16794: result <= 12'b011111111110;
   16795: result <= 12'b011111111110;
   16796: result <= 12'b011111111110;
   16797: result <= 12'b011111111110;
   16798: result <= 12'b011111111110;
   16799: result <= 12'b011111111110;
   16800: result <= 12'b011111111110;
   16801: result <= 12'b011111111110;
   16802: result <= 12'b011111111110;
   16803: result <= 12'b011111111110;
   16804: result <= 12'b011111111110;
   16805: result <= 12'b011111111110;
   16806: result <= 12'b011111111110;
   16807: result <= 12'b011111111110;
   16808: result <= 12'b011111111110;
   16809: result <= 12'b011111111110;
   16810: result <= 12'b011111111110;
   16811: result <= 12'b011111111110;
   16812: result <= 12'b011111111110;
   16813: result <= 12'b011111111110;
   16814: result <= 12'b011111111110;
   16815: result <= 12'b011111111110;
   16816: result <= 12'b011111111110;
   16817: result <= 12'b011111111110;
   16818: result <= 12'b011111111110;
   16819: result <= 12'b011111111110;
   16820: result <= 12'b011111111110;
   16821: result <= 12'b011111111110;
   16822: result <= 12'b011111111110;
   16823: result <= 12'b011111111110;
   16824: result <= 12'b011111111110;
   16825: result <= 12'b011111111110;
   16826: result <= 12'b011111111110;
   16827: result <= 12'b011111111110;
   16828: result <= 12'b011111111110;
   16829: result <= 12'b011111111110;
   16830: result <= 12'b011111111110;
   16831: result <= 12'b011111111110;
   16832: result <= 12'b011111111110;
   16833: result <= 12'b011111111110;
   16834: result <= 12'b011111111110;
   16835: result <= 12'b011111111110;
   16836: result <= 12'b011111111110;
   16837: result <= 12'b011111111110;
   16838: result <= 12'b011111111110;
   16839: result <= 12'b011111111110;
   16840: result <= 12'b011111111110;
   16841: result <= 12'b011111111110;
   16842: result <= 12'b011111111110;
   16843: result <= 12'b011111111110;
   16844: result <= 12'b011111111110;
   16845: result <= 12'b011111111101;
   16846: result <= 12'b011111111101;
   16847: result <= 12'b011111111101;
   16848: result <= 12'b011111111101;
   16849: result <= 12'b011111111101;
   16850: result <= 12'b011111111101;
   16851: result <= 12'b011111111101;
   16852: result <= 12'b011111111101;
   16853: result <= 12'b011111111101;
   16854: result <= 12'b011111111101;
   16855: result <= 12'b011111111101;
   16856: result <= 12'b011111111101;
   16857: result <= 12'b011111111101;
   16858: result <= 12'b011111111101;
   16859: result <= 12'b011111111101;
   16860: result <= 12'b011111111101;
   16861: result <= 12'b011111111101;
   16862: result <= 12'b011111111101;
   16863: result <= 12'b011111111101;
   16864: result <= 12'b011111111101;
   16865: result <= 12'b011111111101;
   16866: result <= 12'b011111111101;
   16867: result <= 12'b011111111101;
   16868: result <= 12'b011111111101;
   16869: result <= 12'b011111111101;
   16870: result <= 12'b011111111101;
   16871: result <= 12'b011111111101;
   16872: result <= 12'b011111111101;
   16873: result <= 12'b011111111101;
   16874: result <= 12'b011111111101;
   16875: result <= 12'b011111111101;
   16876: result <= 12'b011111111101;
   16877: result <= 12'b011111111101;
   16878: result <= 12'b011111111101;
   16879: result <= 12'b011111111101;
   16880: result <= 12'b011111111101;
   16881: result <= 12'b011111111101;
   16882: result <= 12'b011111111101;
   16883: result <= 12'b011111111101;
   16884: result <= 12'b011111111101;
   16885: result <= 12'b011111111101;
   16886: result <= 12'b011111111101;
   16887: result <= 12'b011111111101;
   16888: result <= 12'b011111111101;
   16889: result <= 12'b011111111101;
   16890: result <= 12'b011111111101;
   16891: result <= 12'b011111111101;
   16892: result <= 12'b011111111101;
   16893: result <= 12'b011111111101;
   16894: result <= 12'b011111111101;
   16895: result <= 12'b011111111101;
   16896: result <= 12'b011111111101;
   16897: result <= 12'b011111111101;
   16898: result <= 12'b011111111101;
   16899: result <= 12'b011111111101;
   16900: result <= 12'b011111111101;
   16901: result <= 12'b011111111101;
   16902: result <= 12'b011111111101;
   16903: result <= 12'b011111111101;
   16904: result <= 12'b011111111101;
   16905: result <= 12'b011111111101;
   16906: result <= 12'b011111111101;
   16907: result <= 12'b011111111101;
   16908: result <= 12'b011111111101;
   16909: result <= 12'b011111111101;
   16910: result <= 12'b011111111101;
   16911: result <= 12'b011111111101;
   16912: result <= 12'b011111111101;
   16913: result <= 12'b011111111101;
   16914: result <= 12'b011111111101;
   16915: result <= 12'b011111111101;
   16916: result <= 12'b011111111101;
   16917: result <= 12'b011111111101;
   16918: result <= 12'b011111111101;
   16919: result <= 12'b011111111101;
   16920: result <= 12'b011111111101;
   16921: result <= 12'b011111111101;
   16922: result <= 12'b011111111101;
   16923: result <= 12'b011111111101;
   16924: result <= 12'b011111111101;
   16925: result <= 12'b011111111101;
   16926: result <= 12'b011111111101;
   16927: result <= 12'b011111111101;
   16928: result <= 12'b011111111101;
   16929: result <= 12'b011111111101;
   16930: result <= 12'b011111111101;
   16931: result <= 12'b011111111101;
   16932: result <= 12'b011111111101;
   16933: result <= 12'b011111111101;
   16934: result <= 12'b011111111101;
   16935: result <= 12'b011111111101;
   16936: result <= 12'b011111111101;
   16937: result <= 12'b011111111101;
   16938: result <= 12'b011111111101;
   16939: result <= 12'b011111111101;
   16940: result <= 12'b011111111101;
   16941: result <= 12'b011111111101;
   16942: result <= 12'b011111111101;
   16943: result <= 12'b011111111101;
   16944: result <= 12'b011111111101;
   16945: result <= 12'b011111111101;
   16946: result <= 12'b011111111101;
   16947: result <= 12'b011111111101;
   16948: result <= 12'b011111111101;
   16949: result <= 12'b011111111100;
   16950: result <= 12'b011111111100;
   16951: result <= 12'b011111111100;
   16952: result <= 12'b011111111100;
   16953: result <= 12'b011111111100;
   16954: result <= 12'b011111111100;
   16955: result <= 12'b011111111100;
   16956: result <= 12'b011111111100;
   16957: result <= 12'b011111111100;
   16958: result <= 12'b011111111100;
   16959: result <= 12'b011111111100;
   16960: result <= 12'b011111111100;
   16961: result <= 12'b011111111100;
   16962: result <= 12'b011111111100;
   16963: result <= 12'b011111111100;
   16964: result <= 12'b011111111100;
   16965: result <= 12'b011111111100;
   16966: result <= 12'b011111111100;
   16967: result <= 12'b011111111100;
   16968: result <= 12'b011111111100;
   16969: result <= 12'b011111111100;
   16970: result <= 12'b011111111100;
   16971: result <= 12'b011111111100;
   16972: result <= 12'b011111111100;
   16973: result <= 12'b011111111100;
   16974: result <= 12'b011111111100;
   16975: result <= 12'b011111111100;
   16976: result <= 12'b011111111100;
   16977: result <= 12'b011111111100;
   16978: result <= 12'b011111111100;
   16979: result <= 12'b011111111100;
   16980: result <= 12'b011111111100;
   16981: result <= 12'b011111111100;
   16982: result <= 12'b011111111100;
   16983: result <= 12'b011111111100;
   16984: result <= 12'b011111111100;
   16985: result <= 12'b011111111100;
   16986: result <= 12'b011111111100;
   16987: result <= 12'b011111111100;
   16988: result <= 12'b011111111100;
   16989: result <= 12'b011111111100;
   16990: result <= 12'b011111111100;
   16991: result <= 12'b011111111100;
   16992: result <= 12'b011111111100;
   16993: result <= 12'b011111111100;
   16994: result <= 12'b011111111100;
   16995: result <= 12'b011111111100;
   16996: result <= 12'b011111111100;
   16997: result <= 12'b011111111100;
   16998: result <= 12'b011111111100;
   16999: result <= 12'b011111111100;
   17000: result <= 12'b011111111100;
   17001: result <= 12'b011111111100;
   17002: result <= 12'b011111111100;
   17003: result <= 12'b011111111100;
   17004: result <= 12'b011111111100;
   17005: result <= 12'b011111111100;
   17006: result <= 12'b011111111100;
   17007: result <= 12'b011111111100;
   17008: result <= 12'b011111111100;
   17009: result <= 12'b011111111100;
   17010: result <= 12'b011111111100;
   17011: result <= 12'b011111111100;
   17012: result <= 12'b011111111100;
   17013: result <= 12'b011111111100;
   17014: result <= 12'b011111111100;
   17015: result <= 12'b011111111100;
   17016: result <= 12'b011111111100;
   17017: result <= 12'b011111111100;
   17018: result <= 12'b011111111100;
   17019: result <= 12'b011111111100;
   17020: result <= 12'b011111111100;
   17021: result <= 12'b011111111100;
   17022: result <= 12'b011111111100;
   17023: result <= 12'b011111111100;
   17024: result <= 12'b011111111100;
   17025: result <= 12'b011111111100;
   17026: result <= 12'b011111111100;
   17027: result <= 12'b011111111100;
   17028: result <= 12'b011111111100;
   17029: result <= 12'b011111111100;
   17030: result <= 12'b011111111100;
   17031: result <= 12'b011111111100;
   17032: result <= 12'b011111111100;
   17033: result <= 12'b011111111100;
   17034: result <= 12'b011111111100;
   17035: result <= 12'b011111111100;
   17036: result <= 12'b011111111100;
   17037: result <= 12'b011111111011;
   17038: result <= 12'b011111111011;
   17039: result <= 12'b011111111011;
   17040: result <= 12'b011111111011;
   17041: result <= 12'b011111111011;
   17042: result <= 12'b011111111011;
   17043: result <= 12'b011111111011;
   17044: result <= 12'b011111111011;
   17045: result <= 12'b011111111011;
   17046: result <= 12'b011111111011;
   17047: result <= 12'b011111111011;
   17048: result <= 12'b011111111011;
   17049: result <= 12'b011111111011;
   17050: result <= 12'b011111111011;
   17051: result <= 12'b011111111011;
   17052: result <= 12'b011111111011;
   17053: result <= 12'b011111111011;
   17054: result <= 12'b011111111011;
   17055: result <= 12'b011111111011;
   17056: result <= 12'b011111111011;
   17057: result <= 12'b011111111011;
   17058: result <= 12'b011111111011;
   17059: result <= 12'b011111111011;
   17060: result <= 12'b011111111011;
   17061: result <= 12'b011111111011;
   17062: result <= 12'b011111111011;
   17063: result <= 12'b011111111011;
   17064: result <= 12'b011111111011;
   17065: result <= 12'b011111111011;
   17066: result <= 12'b011111111011;
   17067: result <= 12'b011111111011;
   17068: result <= 12'b011111111011;
   17069: result <= 12'b011111111011;
   17070: result <= 12'b011111111011;
   17071: result <= 12'b011111111011;
   17072: result <= 12'b011111111011;
   17073: result <= 12'b011111111011;
   17074: result <= 12'b011111111011;
   17075: result <= 12'b011111111011;
   17076: result <= 12'b011111111011;
   17077: result <= 12'b011111111011;
   17078: result <= 12'b011111111011;
   17079: result <= 12'b011111111011;
   17080: result <= 12'b011111111011;
   17081: result <= 12'b011111111011;
   17082: result <= 12'b011111111011;
   17083: result <= 12'b011111111011;
   17084: result <= 12'b011111111011;
   17085: result <= 12'b011111111011;
   17086: result <= 12'b011111111011;
   17087: result <= 12'b011111111011;
   17088: result <= 12'b011111111011;
   17089: result <= 12'b011111111011;
   17090: result <= 12'b011111111011;
   17091: result <= 12'b011111111011;
   17092: result <= 12'b011111111011;
   17093: result <= 12'b011111111011;
   17094: result <= 12'b011111111011;
   17095: result <= 12'b011111111011;
   17096: result <= 12'b011111111011;
   17097: result <= 12'b011111111011;
   17098: result <= 12'b011111111011;
   17099: result <= 12'b011111111011;
   17100: result <= 12'b011111111011;
   17101: result <= 12'b011111111011;
   17102: result <= 12'b011111111011;
   17103: result <= 12'b011111111011;
   17104: result <= 12'b011111111011;
   17105: result <= 12'b011111111011;
   17106: result <= 12'b011111111011;
   17107: result <= 12'b011111111011;
   17108: result <= 12'b011111111011;
   17109: result <= 12'b011111111011;
   17110: result <= 12'b011111111011;
   17111: result <= 12'b011111111011;
   17112: result <= 12'b011111111011;
   17113: result <= 12'b011111111010;
   17114: result <= 12'b011111111010;
   17115: result <= 12'b011111111010;
   17116: result <= 12'b011111111010;
   17117: result <= 12'b011111111010;
   17118: result <= 12'b011111111010;
   17119: result <= 12'b011111111010;
   17120: result <= 12'b011111111010;
   17121: result <= 12'b011111111010;
   17122: result <= 12'b011111111010;
   17123: result <= 12'b011111111010;
   17124: result <= 12'b011111111010;
   17125: result <= 12'b011111111010;
   17126: result <= 12'b011111111010;
   17127: result <= 12'b011111111010;
   17128: result <= 12'b011111111010;
   17129: result <= 12'b011111111010;
   17130: result <= 12'b011111111010;
   17131: result <= 12'b011111111010;
   17132: result <= 12'b011111111010;
   17133: result <= 12'b011111111010;
   17134: result <= 12'b011111111010;
   17135: result <= 12'b011111111010;
   17136: result <= 12'b011111111010;
   17137: result <= 12'b011111111010;
   17138: result <= 12'b011111111010;
   17139: result <= 12'b011111111010;
   17140: result <= 12'b011111111010;
   17141: result <= 12'b011111111010;
   17142: result <= 12'b011111111010;
   17143: result <= 12'b011111111010;
   17144: result <= 12'b011111111010;
   17145: result <= 12'b011111111010;
   17146: result <= 12'b011111111010;
   17147: result <= 12'b011111111010;
   17148: result <= 12'b011111111010;
   17149: result <= 12'b011111111010;
   17150: result <= 12'b011111111010;
   17151: result <= 12'b011111111010;
   17152: result <= 12'b011111111010;
   17153: result <= 12'b011111111010;
   17154: result <= 12'b011111111010;
   17155: result <= 12'b011111111010;
   17156: result <= 12'b011111111010;
   17157: result <= 12'b011111111010;
   17158: result <= 12'b011111111010;
   17159: result <= 12'b011111111010;
   17160: result <= 12'b011111111010;
   17161: result <= 12'b011111111010;
   17162: result <= 12'b011111111010;
   17163: result <= 12'b011111111010;
   17164: result <= 12'b011111111010;
   17165: result <= 12'b011111111010;
   17166: result <= 12'b011111111010;
   17167: result <= 12'b011111111010;
   17168: result <= 12'b011111111010;
   17169: result <= 12'b011111111010;
   17170: result <= 12'b011111111010;
   17171: result <= 12'b011111111010;
   17172: result <= 12'b011111111010;
   17173: result <= 12'b011111111010;
   17174: result <= 12'b011111111010;
   17175: result <= 12'b011111111010;
   17176: result <= 12'b011111111010;
   17177: result <= 12'b011111111010;
   17178: result <= 12'b011111111010;
   17179: result <= 12'b011111111010;
   17180: result <= 12'b011111111010;
   17181: result <= 12'b011111111010;
   17182: result <= 12'b011111111010;
   17183: result <= 12'b011111111001;
   17184: result <= 12'b011111111001;
   17185: result <= 12'b011111111001;
   17186: result <= 12'b011111111001;
   17187: result <= 12'b011111111001;
   17188: result <= 12'b011111111001;
   17189: result <= 12'b011111111001;
   17190: result <= 12'b011111111001;
   17191: result <= 12'b011111111001;
   17192: result <= 12'b011111111001;
   17193: result <= 12'b011111111001;
   17194: result <= 12'b011111111001;
   17195: result <= 12'b011111111001;
   17196: result <= 12'b011111111001;
   17197: result <= 12'b011111111001;
   17198: result <= 12'b011111111001;
   17199: result <= 12'b011111111001;
   17200: result <= 12'b011111111001;
   17201: result <= 12'b011111111001;
   17202: result <= 12'b011111111001;
   17203: result <= 12'b011111111001;
   17204: result <= 12'b011111111001;
   17205: result <= 12'b011111111001;
   17206: result <= 12'b011111111001;
   17207: result <= 12'b011111111001;
   17208: result <= 12'b011111111001;
   17209: result <= 12'b011111111001;
   17210: result <= 12'b011111111001;
   17211: result <= 12'b011111111001;
   17212: result <= 12'b011111111001;
   17213: result <= 12'b011111111001;
   17214: result <= 12'b011111111001;
   17215: result <= 12'b011111111001;
   17216: result <= 12'b011111111001;
   17217: result <= 12'b011111111001;
   17218: result <= 12'b011111111001;
   17219: result <= 12'b011111111001;
   17220: result <= 12'b011111111001;
   17221: result <= 12'b011111111001;
   17222: result <= 12'b011111111001;
   17223: result <= 12'b011111111001;
   17224: result <= 12'b011111111001;
   17225: result <= 12'b011111111001;
   17226: result <= 12'b011111111001;
   17227: result <= 12'b011111111001;
   17228: result <= 12'b011111111001;
   17229: result <= 12'b011111111001;
   17230: result <= 12'b011111111001;
   17231: result <= 12'b011111111001;
   17232: result <= 12'b011111111001;
   17233: result <= 12'b011111111001;
   17234: result <= 12'b011111111001;
   17235: result <= 12'b011111111001;
   17236: result <= 12'b011111111001;
   17237: result <= 12'b011111111001;
   17238: result <= 12'b011111111001;
   17239: result <= 12'b011111111001;
   17240: result <= 12'b011111111001;
   17241: result <= 12'b011111111001;
   17242: result <= 12'b011111111001;
   17243: result <= 12'b011111111001;
   17244: result <= 12'b011111111001;
   17245: result <= 12'b011111111001;
   17246: result <= 12'b011111111001;
   17247: result <= 12'b011111111000;
   17248: result <= 12'b011111111000;
   17249: result <= 12'b011111111000;
   17250: result <= 12'b011111111000;
   17251: result <= 12'b011111111000;
   17252: result <= 12'b011111111000;
   17253: result <= 12'b011111111000;
   17254: result <= 12'b011111111000;
   17255: result <= 12'b011111111000;
   17256: result <= 12'b011111111000;
   17257: result <= 12'b011111111000;
   17258: result <= 12'b011111111000;
   17259: result <= 12'b011111111000;
   17260: result <= 12'b011111111000;
   17261: result <= 12'b011111111000;
   17262: result <= 12'b011111111000;
   17263: result <= 12'b011111111000;
   17264: result <= 12'b011111111000;
   17265: result <= 12'b011111111000;
   17266: result <= 12'b011111111000;
   17267: result <= 12'b011111111000;
   17268: result <= 12'b011111111000;
   17269: result <= 12'b011111111000;
   17270: result <= 12'b011111111000;
   17271: result <= 12'b011111111000;
   17272: result <= 12'b011111111000;
   17273: result <= 12'b011111111000;
   17274: result <= 12'b011111111000;
   17275: result <= 12'b011111111000;
   17276: result <= 12'b011111111000;
   17277: result <= 12'b011111111000;
   17278: result <= 12'b011111111000;
   17279: result <= 12'b011111111000;
   17280: result <= 12'b011111111000;
   17281: result <= 12'b011111111000;
   17282: result <= 12'b011111111000;
   17283: result <= 12'b011111111000;
   17284: result <= 12'b011111111000;
   17285: result <= 12'b011111111000;
   17286: result <= 12'b011111111000;
   17287: result <= 12'b011111111000;
   17288: result <= 12'b011111111000;
   17289: result <= 12'b011111111000;
   17290: result <= 12'b011111111000;
   17291: result <= 12'b011111111000;
   17292: result <= 12'b011111111000;
   17293: result <= 12'b011111111000;
   17294: result <= 12'b011111111000;
   17295: result <= 12'b011111111000;
   17296: result <= 12'b011111111000;
   17297: result <= 12'b011111111000;
   17298: result <= 12'b011111111000;
   17299: result <= 12'b011111111000;
   17300: result <= 12'b011111111000;
   17301: result <= 12'b011111111000;
   17302: result <= 12'b011111111000;
   17303: result <= 12'b011111111000;
   17304: result <= 12'b011111111000;
   17305: result <= 12'b011111111000;
   17306: result <= 12'b011111111000;
   17307: result <= 12'b011111110111;
   17308: result <= 12'b011111110111;
   17309: result <= 12'b011111110111;
   17310: result <= 12'b011111110111;
   17311: result <= 12'b011111110111;
   17312: result <= 12'b011111110111;
   17313: result <= 12'b011111110111;
   17314: result <= 12'b011111110111;
   17315: result <= 12'b011111110111;
   17316: result <= 12'b011111110111;
   17317: result <= 12'b011111110111;
   17318: result <= 12'b011111110111;
   17319: result <= 12'b011111110111;
   17320: result <= 12'b011111110111;
   17321: result <= 12'b011111110111;
   17322: result <= 12'b011111110111;
   17323: result <= 12'b011111110111;
   17324: result <= 12'b011111110111;
   17325: result <= 12'b011111110111;
   17326: result <= 12'b011111110111;
   17327: result <= 12'b011111110111;
   17328: result <= 12'b011111110111;
   17329: result <= 12'b011111110111;
   17330: result <= 12'b011111110111;
   17331: result <= 12'b011111110111;
   17332: result <= 12'b011111110111;
   17333: result <= 12'b011111110111;
   17334: result <= 12'b011111110111;
   17335: result <= 12'b011111110111;
   17336: result <= 12'b011111110111;
   17337: result <= 12'b011111110111;
   17338: result <= 12'b011111110111;
   17339: result <= 12'b011111110111;
   17340: result <= 12'b011111110111;
   17341: result <= 12'b011111110111;
   17342: result <= 12'b011111110111;
   17343: result <= 12'b011111110111;
   17344: result <= 12'b011111110111;
   17345: result <= 12'b011111110111;
   17346: result <= 12'b011111110111;
   17347: result <= 12'b011111110111;
   17348: result <= 12'b011111110111;
   17349: result <= 12'b011111110111;
   17350: result <= 12'b011111110111;
   17351: result <= 12'b011111110111;
   17352: result <= 12'b011111110111;
   17353: result <= 12'b011111110111;
   17354: result <= 12'b011111110111;
   17355: result <= 12'b011111110111;
   17356: result <= 12'b011111110111;
   17357: result <= 12'b011111110111;
   17358: result <= 12'b011111110111;
   17359: result <= 12'b011111110111;
   17360: result <= 12'b011111110111;
   17361: result <= 12'b011111110111;
   17362: result <= 12'b011111110111;
   17363: result <= 12'b011111110110;
   17364: result <= 12'b011111110110;
   17365: result <= 12'b011111110110;
   17366: result <= 12'b011111110110;
   17367: result <= 12'b011111110110;
   17368: result <= 12'b011111110110;
   17369: result <= 12'b011111110110;
   17370: result <= 12'b011111110110;
   17371: result <= 12'b011111110110;
   17372: result <= 12'b011111110110;
   17373: result <= 12'b011111110110;
   17374: result <= 12'b011111110110;
   17375: result <= 12'b011111110110;
   17376: result <= 12'b011111110110;
   17377: result <= 12'b011111110110;
   17378: result <= 12'b011111110110;
   17379: result <= 12'b011111110110;
   17380: result <= 12'b011111110110;
   17381: result <= 12'b011111110110;
   17382: result <= 12'b011111110110;
   17383: result <= 12'b011111110110;
   17384: result <= 12'b011111110110;
   17385: result <= 12'b011111110110;
   17386: result <= 12'b011111110110;
   17387: result <= 12'b011111110110;
   17388: result <= 12'b011111110110;
   17389: result <= 12'b011111110110;
   17390: result <= 12'b011111110110;
   17391: result <= 12'b011111110110;
   17392: result <= 12'b011111110110;
   17393: result <= 12'b011111110110;
   17394: result <= 12'b011111110110;
   17395: result <= 12'b011111110110;
   17396: result <= 12'b011111110110;
   17397: result <= 12'b011111110110;
   17398: result <= 12'b011111110110;
   17399: result <= 12'b011111110110;
   17400: result <= 12'b011111110110;
   17401: result <= 12'b011111110110;
   17402: result <= 12'b011111110110;
   17403: result <= 12'b011111110110;
   17404: result <= 12'b011111110110;
   17405: result <= 12'b011111110110;
   17406: result <= 12'b011111110110;
   17407: result <= 12'b011111110110;
   17408: result <= 12'b011111110110;
   17409: result <= 12'b011111110110;
   17410: result <= 12'b011111110110;
   17411: result <= 12'b011111110110;
   17412: result <= 12'b011111110110;
   17413: result <= 12'b011111110110;
   17414: result <= 12'b011111110110;
   17415: result <= 12'b011111110110;
   17416: result <= 12'b011111110101;
   17417: result <= 12'b011111110101;
   17418: result <= 12'b011111110101;
   17419: result <= 12'b011111110101;
   17420: result <= 12'b011111110101;
   17421: result <= 12'b011111110101;
   17422: result <= 12'b011111110101;
   17423: result <= 12'b011111110101;
   17424: result <= 12'b011111110101;
   17425: result <= 12'b011111110101;
   17426: result <= 12'b011111110101;
   17427: result <= 12'b011111110101;
   17428: result <= 12'b011111110101;
   17429: result <= 12'b011111110101;
   17430: result <= 12'b011111110101;
   17431: result <= 12'b011111110101;
   17432: result <= 12'b011111110101;
   17433: result <= 12'b011111110101;
   17434: result <= 12'b011111110101;
   17435: result <= 12'b011111110101;
   17436: result <= 12'b011111110101;
   17437: result <= 12'b011111110101;
   17438: result <= 12'b011111110101;
   17439: result <= 12'b011111110101;
   17440: result <= 12'b011111110101;
   17441: result <= 12'b011111110101;
   17442: result <= 12'b011111110101;
   17443: result <= 12'b011111110101;
   17444: result <= 12'b011111110101;
   17445: result <= 12'b011111110101;
   17446: result <= 12'b011111110101;
   17447: result <= 12'b011111110101;
   17448: result <= 12'b011111110101;
   17449: result <= 12'b011111110101;
   17450: result <= 12'b011111110101;
   17451: result <= 12'b011111110101;
   17452: result <= 12'b011111110101;
   17453: result <= 12'b011111110101;
   17454: result <= 12'b011111110101;
   17455: result <= 12'b011111110101;
   17456: result <= 12'b011111110101;
   17457: result <= 12'b011111110101;
   17458: result <= 12'b011111110101;
   17459: result <= 12'b011111110101;
   17460: result <= 12'b011111110101;
   17461: result <= 12'b011111110101;
   17462: result <= 12'b011111110101;
   17463: result <= 12'b011111110101;
   17464: result <= 12'b011111110101;
   17465: result <= 12'b011111110101;
   17466: result <= 12'b011111110100;
   17467: result <= 12'b011111110100;
   17468: result <= 12'b011111110100;
   17469: result <= 12'b011111110100;
   17470: result <= 12'b011111110100;
   17471: result <= 12'b011111110100;
   17472: result <= 12'b011111110100;
   17473: result <= 12'b011111110100;
   17474: result <= 12'b011111110100;
   17475: result <= 12'b011111110100;
   17476: result <= 12'b011111110100;
   17477: result <= 12'b011111110100;
   17478: result <= 12'b011111110100;
   17479: result <= 12'b011111110100;
   17480: result <= 12'b011111110100;
   17481: result <= 12'b011111110100;
   17482: result <= 12'b011111110100;
   17483: result <= 12'b011111110100;
   17484: result <= 12'b011111110100;
   17485: result <= 12'b011111110100;
   17486: result <= 12'b011111110100;
   17487: result <= 12'b011111110100;
   17488: result <= 12'b011111110100;
   17489: result <= 12'b011111110100;
   17490: result <= 12'b011111110100;
   17491: result <= 12'b011111110100;
   17492: result <= 12'b011111110100;
   17493: result <= 12'b011111110100;
   17494: result <= 12'b011111110100;
   17495: result <= 12'b011111110100;
   17496: result <= 12'b011111110100;
   17497: result <= 12'b011111110100;
   17498: result <= 12'b011111110100;
   17499: result <= 12'b011111110100;
   17500: result <= 12'b011111110100;
   17501: result <= 12'b011111110100;
   17502: result <= 12'b011111110100;
   17503: result <= 12'b011111110100;
   17504: result <= 12'b011111110100;
   17505: result <= 12'b011111110100;
   17506: result <= 12'b011111110100;
   17507: result <= 12'b011111110100;
   17508: result <= 12'b011111110100;
   17509: result <= 12'b011111110100;
   17510: result <= 12'b011111110100;
   17511: result <= 12'b011111110100;
   17512: result <= 12'b011111110100;
   17513: result <= 12'b011111110100;
   17514: result <= 12'b011111110011;
   17515: result <= 12'b011111110011;
   17516: result <= 12'b011111110011;
   17517: result <= 12'b011111110011;
   17518: result <= 12'b011111110011;
   17519: result <= 12'b011111110011;
   17520: result <= 12'b011111110011;
   17521: result <= 12'b011111110011;
   17522: result <= 12'b011111110011;
   17523: result <= 12'b011111110011;
   17524: result <= 12'b011111110011;
   17525: result <= 12'b011111110011;
   17526: result <= 12'b011111110011;
   17527: result <= 12'b011111110011;
   17528: result <= 12'b011111110011;
   17529: result <= 12'b011111110011;
   17530: result <= 12'b011111110011;
   17531: result <= 12'b011111110011;
   17532: result <= 12'b011111110011;
   17533: result <= 12'b011111110011;
   17534: result <= 12'b011111110011;
   17535: result <= 12'b011111110011;
   17536: result <= 12'b011111110011;
   17537: result <= 12'b011111110011;
   17538: result <= 12'b011111110011;
   17539: result <= 12'b011111110011;
   17540: result <= 12'b011111110011;
   17541: result <= 12'b011111110011;
   17542: result <= 12'b011111110011;
   17543: result <= 12'b011111110011;
   17544: result <= 12'b011111110011;
   17545: result <= 12'b011111110011;
   17546: result <= 12'b011111110011;
   17547: result <= 12'b011111110011;
   17548: result <= 12'b011111110011;
   17549: result <= 12'b011111110011;
   17550: result <= 12'b011111110011;
   17551: result <= 12'b011111110011;
   17552: result <= 12'b011111110011;
   17553: result <= 12'b011111110011;
   17554: result <= 12'b011111110011;
   17555: result <= 12'b011111110011;
   17556: result <= 12'b011111110011;
   17557: result <= 12'b011111110011;
   17558: result <= 12'b011111110011;
   17559: result <= 12'b011111110011;
   17560: result <= 12'b011111110010;
   17561: result <= 12'b011111110010;
   17562: result <= 12'b011111110010;
   17563: result <= 12'b011111110010;
   17564: result <= 12'b011111110010;
   17565: result <= 12'b011111110010;
   17566: result <= 12'b011111110010;
   17567: result <= 12'b011111110010;
   17568: result <= 12'b011111110010;
   17569: result <= 12'b011111110010;
   17570: result <= 12'b011111110010;
   17571: result <= 12'b011111110010;
   17572: result <= 12'b011111110010;
   17573: result <= 12'b011111110010;
   17574: result <= 12'b011111110010;
   17575: result <= 12'b011111110010;
   17576: result <= 12'b011111110010;
   17577: result <= 12'b011111110010;
   17578: result <= 12'b011111110010;
   17579: result <= 12'b011111110010;
   17580: result <= 12'b011111110010;
   17581: result <= 12'b011111110010;
   17582: result <= 12'b011111110010;
   17583: result <= 12'b011111110010;
   17584: result <= 12'b011111110010;
   17585: result <= 12'b011111110010;
   17586: result <= 12'b011111110010;
   17587: result <= 12'b011111110010;
   17588: result <= 12'b011111110010;
   17589: result <= 12'b011111110010;
   17590: result <= 12'b011111110010;
   17591: result <= 12'b011111110010;
   17592: result <= 12'b011111110010;
   17593: result <= 12'b011111110010;
   17594: result <= 12'b011111110010;
   17595: result <= 12'b011111110010;
   17596: result <= 12'b011111110010;
   17597: result <= 12'b011111110010;
   17598: result <= 12'b011111110010;
   17599: result <= 12'b011111110010;
   17600: result <= 12'b011111110010;
   17601: result <= 12'b011111110010;
   17602: result <= 12'b011111110010;
   17603: result <= 12'b011111110010;
   17604: result <= 12'b011111110010;
   17605: result <= 12'b011111110001;
   17606: result <= 12'b011111110001;
   17607: result <= 12'b011111110001;
   17608: result <= 12'b011111110001;
   17609: result <= 12'b011111110001;
   17610: result <= 12'b011111110001;
   17611: result <= 12'b011111110001;
   17612: result <= 12'b011111110001;
   17613: result <= 12'b011111110001;
   17614: result <= 12'b011111110001;
   17615: result <= 12'b011111110001;
   17616: result <= 12'b011111110001;
   17617: result <= 12'b011111110001;
   17618: result <= 12'b011111110001;
   17619: result <= 12'b011111110001;
   17620: result <= 12'b011111110001;
   17621: result <= 12'b011111110001;
   17622: result <= 12'b011111110001;
   17623: result <= 12'b011111110001;
   17624: result <= 12'b011111110001;
   17625: result <= 12'b011111110001;
   17626: result <= 12'b011111110001;
   17627: result <= 12'b011111110001;
   17628: result <= 12'b011111110001;
   17629: result <= 12'b011111110001;
   17630: result <= 12'b011111110001;
   17631: result <= 12'b011111110001;
   17632: result <= 12'b011111110001;
   17633: result <= 12'b011111110001;
   17634: result <= 12'b011111110001;
   17635: result <= 12'b011111110001;
   17636: result <= 12'b011111110001;
   17637: result <= 12'b011111110001;
   17638: result <= 12'b011111110001;
   17639: result <= 12'b011111110001;
   17640: result <= 12'b011111110001;
   17641: result <= 12'b011111110001;
   17642: result <= 12'b011111110001;
   17643: result <= 12'b011111110001;
   17644: result <= 12'b011111110001;
   17645: result <= 12'b011111110001;
   17646: result <= 12'b011111110001;
   17647: result <= 12'b011111110001;
   17648: result <= 12'b011111110000;
   17649: result <= 12'b011111110000;
   17650: result <= 12'b011111110000;
   17651: result <= 12'b011111110000;
   17652: result <= 12'b011111110000;
   17653: result <= 12'b011111110000;
   17654: result <= 12'b011111110000;
   17655: result <= 12'b011111110000;
   17656: result <= 12'b011111110000;
   17657: result <= 12'b011111110000;
   17658: result <= 12'b011111110000;
   17659: result <= 12'b011111110000;
   17660: result <= 12'b011111110000;
   17661: result <= 12'b011111110000;
   17662: result <= 12'b011111110000;
   17663: result <= 12'b011111110000;
   17664: result <= 12'b011111110000;
   17665: result <= 12'b011111110000;
   17666: result <= 12'b011111110000;
   17667: result <= 12'b011111110000;
   17668: result <= 12'b011111110000;
   17669: result <= 12'b011111110000;
   17670: result <= 12'b011111110000;
   17671: result <= 12'b011111110000;
   17672: result <= 12'b011111110000;
   17673: result <= 12'b011111110000;
   17674: result <= 12'b011111110000;
   17675: result <= 12'b011111110000;
   17676: result <= 12'b011111110000;
   17677: result <= 12'b011111110000;
   17678: result <= 12'b011111110000;
   17679: result <= 12'b011111110000;
   17680: result <= 12'b011111110000;
   17681: result <= 12'b011111110000;
   17682: result <= 12'b011111110000;
   17683: result <= 12'b011111110000;
   17684: result <= 12'b011111110000;
   17685: result <= 12'b011111110000;
   17686: result <= 12'b011111110000;
   17687: result <= 12'b011111110000;
   17688: result <= 12'b011111110000;
   17689: result <= 12'b011111101111;
   17690: result <= 12'b011111101111;
   17691: result <= 12'b011111101111;
   17692: result <= 12'b011111101111;
   17693: result <= 12'b011111101111;
   17694: result <= 12'b011111101111;
   17695: result <= 12'b011111101111;
   17696: result <= 12'b011111101111;
   17697: result <= 12'b011111101111;
   17698: result <= 12'b011111101111;
   17699: result <= 12'b011111101111;
   17700: result <= 12'b011111101111;
   17701: result <= 12'b011111101111;
   17702: result <= 12'b011111101111;
   17703: result <= 12'b011111101111;
   17704: result <= 12'b011111101111;
   17705: result <= 12'b011111101111;
   17706: result <= 12'b011111101111;
   17707: result <= 12'b011111101111;
   17708: result <= 12'b011111101111;
   17709: result <= 12'b011111101111;
   17710: result <= 12'b011111101111;
   17711: result <= 12'b011111101111;
   17712: result <= 12'b011111101111;
   17713: result <= 12'b011111101111;
   17714: result <= 12'b011111101111;
   17715: result <= 12'b011111101111;
   17716: result <= 12'b011111101111;
   17717: result <= 12'b011111101111;
   17718: result <= 12'b011111101111;
   17719: result <= 12'b011111101111;
   17720: result <= 12'b011111101111;
   17721: result <= 12'b011111101111;
   17722: result <= 12'b011111101111;
   17723: result <= 12'b011111101111;
   17724: result <= 12'b011111101111;
   17725: result <= 12'b011111101111;
   17726: result <= 12'b011111101111;
   17727: result <= 12'b011111101111;
   17728: result <= 12'b011111101111;
   17729: result <= 12'b011111101110;
   17730: result <= 12'b011111101110;
   17731: result <= 12'b011111101110;
   17732: result <= 12'b011111101110;
   17733: result <= 12'b011111101110;
   17734: result <= 12'b011111101110;
   17735: result <= 12'b011111101110;
   17736: result <= 12'b011111101110;
   17737: result <= 12'b011111101110;
   17738: result <= 12'b011111101110;
   17739: result <= 12'b011111101110;
   17740: result <= 12'b011111101110;
   17741: result <= 12'b011111101110;
   17742: result <= 12'b011111101110;
   17743: result <= 12'b011111101110;
   17744: result <= 12'b011111101110;
   17745: result <= 12'b011111101110;
   17746: result <= 12'b011111101110;
   17747: result <= 12'b011111101110;
   17748: result <= 12'b011111101110;
   17749: result <= 12'b011111101110;
   17750: result <= 12'b011111101110;
   17751: result <= 12'b011111101110;
   17752: result <= 12'b011111101110;
   17753: result <= 12'b011111101110;
   17754: result <= 12'b011111101110;
   17755: result <= 12'b011111101110;
   17756: result <= 12'b011111101110;
   17757: result <= 12'b011111101110;
   17758: result <= 12'b011111101110;
   17759: result <= 12'b011111101110;
   17760: result <= 12'b011111101110;
   17761: result <= 12'b011111101110;
   17762: result <= 12'b011111101110;
   17763: result <= 12'b011111101110;
   17764: result <= 12'b011111101110;
   17765: result <= 12'b011111101110;
   17766: result <= 12'b011111101110;
   17767: result <= 12'b011111101110;
   17768: result <= 12'b011111101101;
   17769: result <= 12'b011111101101;
   17770: result <= 12'b011111101101;
   17771: result <= 12'b011111101101;
   17772: result <= 12'b011111101101;
   17773: result <= 12'b011111101101;
   17774: result <= 12'b011111101101;
   17775: result <= 12'b011111101101;
   17776: result <= 12'b011111101101;
   17777: result <= 12'b011111101101;
   17778: result <= 12'b011111101101;
   17779: result <= 12'b011111101101;
   17780: result <= 12'b011111101101;
   17781: result <= 12'b011111101101;
   17782: result <= 12'b011111101101;
   17783: result <= 12'b011111101101;
   17784: result <= 12'b011111101101;
   17785: result <= 12'b011111101101;
   17786: result <= 12'b011111101101;
   17787: result <= 12'b011111101101;
   17788: result <= 12'b011111101101;
   17789: result <= 12'b011111101101;
   17790: result <= 12'b011111101101;
   17791: result <= 12'b011111101101;
   17792: result <= 12'b011111101101;
   17793: result <= 12'b011111101101;
   17794: result <= 12'b011111101101;
   17795: result <= 12'b011111101101;
   17796: result <= 12'b011111101101;
   17797: result <= 12'b011111101101;
   17798: result <= 12'b011111101101;
   17799: result <= 12'b011111101101;
   17800: result <= 12'b011111101101;
   17801: result <= 12'b011111101101;
   17802: result <= 12'b011111101101;
   17803: result <= 12'b011111101101;
   17804: result <= 12'b011111101101;
   17805: result <= 12'b011111101101;
   17806: result <= 12'b011111101100;
   17807: result <= 12'b011111101100;
   17808: result <= 12'b011111101100;
   17809: result <= 12'b011111101100;
   17810: result <= 12'b011111101100;
   17811: result <= 12'b011111101100;
   17812: result <= 12'b011111101100;
   17813: result <= 12'b011111101100;
   17814: result <= 12'b011111101100;
   17815: result <= 12'b011111101100;
   17816: result <= 12'b011111101100;
   17817: result <= 12'b011111101100;
   17818: result <= 12'b011111101100;
   17819: result <= 12'b011111101100;
   17820: result <= 12'b011111101100;
   17821: result <= 12'b011111101100;
   17822: result <= 12'b011111101100;
   17823: result <= 12'b011111101100;
   17824: result <= 12'b011111101100;
   17825: result <= 12'b011111101100;
   17826: result <= 12'b011111101100;
   17827: result <= 12'b011111101100;
   17828: result <= 12'b011111101100;
   17829: result <= 12'b011111101100;
   17830: result <= 12'b011111101100;
   17831: result <= 12'b011111101100;
   17832: result <= 12'b011111101100;
   17833: result <= 12'b011111101100;
   17834: result <= 12'b011111101100;
   17835: result <= 12'b011111101100;
   17836: result <= 12'b011111101100;
   17837: result <= 12'b011111101100;
   17838: result <= 12'b011111101100;
   17839: result <= 12'b011111101100;
   17840: result <= 12'b011111101100;
   17841: result <= 12'b011111101100;
   17842: result <= 12'b011111101100;
   17843: result <= 12'b011111101011;
   17844: result <= 12'b011111101011;
   17845: result <= 12'b011111101011;
   17846: result <= 12'b011111101011;
   17847: result <= 12'b011111101011;
   17848: result <= 12'b011111101011;
   17849: result <= 12'b011111101011;
   17850: result <= 12'b011111101011;
   17851: result <= 12'b011111101011;
   17852: result <= 12'b011111101011;
   17853: result <= 12'b011111101011;
   17854: result <= 12'b011111101011;
   17855: result <= 12'b011111101011;
   17856: result <= 12'b011111101011;
   17857: result <= 12'b011111101011;
   17858: result <= 12'b011111101011;
   17859: result <= 12'b011111101011;
   17860: result <= 12'b011111101011;
   17861: result <= 12'b011111101011;
   17862: result <= 12'b011111101011;
   17863: result <= 12'b011111101011;
   17864: result <= 12'b011111101011;
   17865: result <= 12'b011111101011;
   17866: result <= 12'b011111101011;
   17867: result <= 12'b011111101011;
   17868: result <= 12'b011111101011;
   17869: result <= 12'b011111101011;
   17870: result <= 12'b011111101011;
   17871: result <= 12'b011111101011;
   17872: result <= 12'b011111101011;
   17873: result <= 12'b011111101011;
   17874: result <= 12'b011111101011;
   17875: result <= 12'b011111101011;
   17876: result <= 12'b011111101011;
   17877: result <= 12'b011111101011;
   17878: result <= 12'b011111101011;
   17879: result <= 12'b011111101010;
   17880: result <= 12'b011111101010;
   17881: result <= 12'b011111101010;
   17882: result <= 12'b011111101010;
   17883: result <= 12'b011111101010;
   17884: result <= 12'b011111101010;
   17885: result <= 12'b011111101010;
   17886: result <= 12'b011111101010;
   17887: result <= 12'b011111101010;
   17888: result <= 12'b011111101010;
   17889: result <= 12'b011111101010;
   17890: result <= 12'b011111101010;
   17891: result <= 12'b011111101010;
   17892: result <= 12'b011111101010;
   17893: result <= 12'b011111101010;
   17894: result <= 12'b011111101010;
   17895: result <= 12'b011111101010;
   17896: result <= 12'b011111101010;
   17897: result <= 12'b011111101010;
   17898: result <= 12'b011111101010;
   17899: result <= 12'b011111101010;
   17900: result <= 12'b011111101010;
   17901: result <= 12'b011111101010;
   17902: result <= 12'b011111101010;
   17903: result <= 12'b011111101010;
   17904: result <= 12'b011111101010;
   17905: result <= 12'b011111101010;
   17906: result <= 12'b011111101010;
   17907: result <= 12'b011111101010;
   17908: result <= 12'b011111101010;
   17909: result <= 12'b011111101010;
   17910: result <= 12'b011111101010;
   17911: result <= 12'b011111101010;
   17912: result <= 12'b011111101010;
   17913: result <= 12'b011111101010;
   17914: result <= 12'b011111101010;
   17915: result <= 12'b011111101001;
   17916: result <= 12'b011111101001;
   17917: result <= 12'b011111101001;
   17918: result <= 12'b011111101001;
   17919: result <= 12'b011111101001;
   17920: result <= 12'b011111101001;
   17921: result <= 12'b011111101001;
   17922: result <= 12'b011111101001;
   17923: result <= 12'b011111101001;
   17924: result <= 12'b011111101001;
   17925: result <= 12'b011111101001;
   17926: result <= 12'b011111101001;
   17927: result <= 12'b011111101001;
   17928: result <= 12'b011111101001;
   17929: result <= 12'b011111101001;
   17930: result <= 12'b011111101001;
   17931: result <= 12'b011111101001;
   17932: result <= 12'b011111101001;
   17933: result <= 12'b011111101001;
   17934: result <= 12'b011111101001;
   17935: result <= 12'b011111101001;
   17936: result <= 12'b011111101001;
   17937: result <= 12'b011111101001;
   17938: result <= 12'b011111101001;
   17939: result <= 12'b011111101001;
   17940: result <= 12'b011111101001;
   17941: result <= 12'b011111101001;
   17942: result <= 12'b011111101001;
   17943: result <= 12'b011111101001;
   17944: result <= 12'b011111101001;
   17945: result <= 12'b011111101001;
   17946: result <= 12'b011111101001;
   17947: result <= 12'b011111101001;
   17948: result <= 12'b011111101001;
   17949: result <= 12'b011111101000;
   17950: result <= 12'b011111101000;
   17951: result <= 12'b011111101000;
   17952: result <= 12'b011111101000;
   17953: result <= 12'b011111101000;
   17954: result <= 12'b011111101000;
   17955: result <= 12'b011111101000;
   17956: result <= 12'b011111101000;
   17957: result <= 12'b011111101000;
   17958: result <= 12'b011111101000;
   17959: result <= 12'b011111101000;
   17960: result <= 12'b011111101000;
   17961: result <= 12'b011111101000;
   17962: result <= 12'b011111101000;
   17963: result <= 12'b011111101000;
   17964: result <= 12'b011111101000;
   17965: result <= 12'b011111101000;
   17966: result <= 12'b011111101000;
   17967: result <= 12'b011111101000;
   17968: result <= 12'b011111101000;
   17969: result <= 12'b011111101000;
   17970: result <= 12'b011111101000;
   17971: result <= 12'b011111101000;
   17972: result <= 12'b011111101000;
   17973: result <= 12'b011111101000;
   17974: result <= 12'b011111101000;
   17975: result <= 12'b011111101000;
   17976: result <= 12'b011111101000;
   17977: result <= 12'b011111101000;
   17978: result <= 12'b011111101000;
   17979: result <= 12'b011111101000;
   17980: result <= 12'b011111101000;
   17981: result <= 12'b011111101000;
   17982: result <= 12'b011111101000;
   17983: result <= 12'b011111100111;
   17984: result <= 12'b011111100111;
   17985: result <= 12'b011111100111;
   17986: result <= 12'b011111100111;
   17987: result <= 12'b011111100111;
   17988: result <= 12'b011111100111;
   17989: result <= 12'b011111100111;
   17990: result <= 12'b011111100111;
   17991: result <= 12'b011111100111;
   17992: result <= 12'b011111100111;
   17993: result <= 12'b011111100111;
   17994: result <= 12'b011111100111;
   17995: result <= 12'b011111100111;
   17996: result <= 12'b011111100111;
   17997: result <= 12'b011111100111;
   17998: result <= 12'b011111100111;
   17999: result <= 12'b011111100111;
   18000: result <= 12'b011111100111;
   18001: result <= 12'b011111100111;
   18002: result <= 12'b011111100111;
   18003: result <= 12'b011111100111;
   18004: result <= 12'b011111100111;
   18005: result <= 12'b011111100111;
   18006: result <= 12'b011111100111;
   18007: result <= 12'b011111100111;
   18008: result <= 12'b011111100111;
   18009: result <= 12'b011111100111;
   18010: result <= 12'b011111100111;
   18011: result <= 12'b011111100111;
   18012: result <= 12'b011111100111;
   18013: result <= 12'b011111100111;
   18014: result <= 12'b011111100111;
   18015: result <= 12'b011111100111;
   18016: result <= 12'b011111100110;
   18017: result <= 12'b011111100110;
   18018: result <= 12'b011111100110;
   18019: result <= 12'b011111100110;
   18020: result <= 12'b011111100110;
   18021: result <= 12'b011111100110;
   18022: result <= 12'b011111100110;
   18023: result <= 12'b011111100110;
   18024: result <= 12'b011111100110;
   18025: result <= 12'b011111100110;
   18026: result <= 12'b011111100110;
   18027: result <= 12'b011111100110;
   18028: result <= 12'b011111100110;
   18029: result <= 12'b011111100110;
   18030: result <= 12'b011111100110;
   18031: result <= 12'b011111100110;
   18032: result <= 12'b011111100110;
   18033: result <= 12'b011111100110;
   18034: result <= 12'b011111100110;
   18035: result <= 12'b011111100110;
   18036: result <= 12'b011111100110;
   18037: result <= 12'b011111100110;
   18038: result <= 12'b011111100110;
   18039: result <= 12'b011111100110;
   18040: result <= 12'b011111100110;
   18041: result <= 12'b011111100110;
   18042: result <= 12'b011111100110;
   18043: result <= 12'b011111100110;
   18044: result <= 12'b011111100110;
   18045: result <= 12'b011111100110;
   18046: result <= 12'b011111100110;
   18047: result <= 12'b011111100110;
   18048: result <= 12'b011111100101;
   18049: result <= 12'b011111100101;
   18050: result <= 12'b011111100101;
   18051: result <= 12'b011111100101;
   18052: result <= 12'b011111100101;
   18053: result <= 12'b011111100101;
   18054: result <= 12'b011111100101;
   18055: result <= 12'b011111100101;
   18056: result <= 12'b011111100101;
   18057: result <= 12'b011111100101;
   18058: result <= 12'b011111100101;
   18059: result <= 12'b011111100101;
   18060: result <= 12'b011111100101;
   18061: result <= 12'b011111100101;
   18062: result <= 12'b011111100101;
   18063: result <= 12'b011111100101;
   18064: result <= 12'b011111100101;
   18065: result <= 12'b011111100101;
   18066: result <= 12'b011111100101;
   18067: result <= 12'b011111100101;
   18068: result <= 12'b011111100101;
   18069: result <= 12'b011111100101;
   18070: result <= 12'b011111100101;
   18071: result <= 12'b011111100101;
   18072: result <= 12'b011111100101;
   18073: result <= 12'b011111100101;
   18074: result <= 12'b011111100101;
   18075: result <= 12'b011111100101;
   18076: result <= 12'b011111100101;
   18077: result <= 12'b011111100101;
   18078: result <= 12'b011111100101;
   18079: result <= 12'b011111100101;
   18080: result <= 12'b011111100100;
   18081: result <= 12'b011111100100;
   18082: result <= 12'b011111100100;
   18083: result <= 12'b011111100100;
   18084: result <= 12'b011111100100;
   18085: result <= 12'b011111100100;
   18086: result <= 12'b011111100100;
   18087: result <= 12'b011111100100;
   18088: result <= 12'b011111100100;
   18089: result <= 12'b011111100100;
   18090: result <= 12'b011111100100;
   18091: result <= 12'b011111100100;
   18092: result <= 12'b011111100100;
   18093: result <= 12'b011111100100;
   18094: result <= 12'b011111100100;
   18095: result <= 12'b011111100100;
   18096: result <= 12'b011111100100;
   18097: result <= 12'b011111100100;
   18098: result <= 12'b011111100100;
   18099: result <= 12'b011111100100;
   18100: result <= 12'b011111100100;
   18101: result <= 12'b011111100100;
   18102: result <= 12'b011111100100;
   18103: result <= 12'b011111100100;
   18104: result <= 12'b011111100100;
   18105: result <= 12'b011111100100;
   18106: result <= 12'b011111100100;
   18107: result <= 12'b011111100100;
   18108: result <= 12'b011111100100;
   18109: result <= 12'b011111100100;
   18110: result <= 12'b011111100100;
   18111: result <= 12'b011111100011;
   18112: result <= 12'b011111100011;
   18113: result <= 12'b011111100011;
   18114: result <= 12'b011111100011;
   18115: result <= 12'b011111100011;
   18116: result <= 12'b011111100011;
   18117: result <= 12'b011111100011;
   18118: result <= 12'b011111100011;
   18119: result <= 12'b011111100011;
   18120: result <= 12'b011111100011;
   18121: result <= 12'b011111100011;
   18122: result <= 12'b011111100011;
   18123: result <= 12'b011111100011;
   18124: result <= 12'b011111100011;
   18125: result <= 12'b011111100011;
   18126: result <= 12'b011111100011;
   18127: result <= 12'b011111100011;
   18128: result <= 12'b011111100011;
   18129: result <= 12'b011111100011;
   18130: result <= 12'b011111100011;
   18131: result <= 12'b011111100011;
   18132: result <= 12'b011111100011;
   18133: result <= 12'b011111100011;
   18134: result <= 12'b011111100011;
   18135: result <= 12'b011111100011;
   18136: result <= 12'b011111100011;
   18137: result <= 12'b011111100011;
   18138: result <= 12'b011111100011;
   18139: result <= 12'b011111100011;
   18140: result <= 12'b011111100011;
   18141: result <= 12'b011111100011;
   18142: result <= 12'b011111100010;
   18143: result <= 12'b011111100010;
   18144: result <= 12'b011111100010;
   18145: result <= 12'b011111100010;
   18146: result <= 12'b011111100010;
   18147: result <= 12'b011111100010;
   18148: result <= 12'b011111100010;
   18149: result <= 12'b011111100010;
   18150: result <= 12'b011111100010;
   18151: result <= 12'b011111100010;
   18152: result <= 12'b011111100010;
   18153: result <= 12'b011111100010;
   18154: result <= 12'b011111100010;
   18155: result <= 12'b011111100010;
   18156: result <= 12'b011111100010;
   18157: result <= 12'b011111100010;
   18158: result <= 12'b011111100010;
   18159: result <= 12'b011111100010;
   18160: result <= 12'b011111100010;
   18161: result <= 12'b011111100010;
   18162: result <= 12'b011111100010;
   18163: result <= 12'b011111100010;
   18164: result <= 12'b011111100010;
   18165: result <= 12'b011111100010;
   18166: result <= 12'b011111100010;
   18167: result <= 12'b011111100010;
   18168: result <= 12'b011111100010;
   18169: result <= 12'b011111100010;
   18170: result <= 12'b011111100010;
   18171: result <= 12'b011111100010;
   18172: result <= 12'b011111100001;
   18173: result <= 12'b011111100001;
   18174: result <= 12'b011111100001;
   18175: result <= 12'b011111100001;
   18176: result <= 12'b011111100001;
   18177: result <= 12'b011111100001;
   18178: result <= 12'b011111100001;
   18179: result <= 12'b011111100001;
   18180: result <= 12'b011111100001;
   18181: result <= 12'b011111100001;
   18182: result <= 12'b011111100001;
   18183: result <= 12'b011111100001;
   18184: result <= 12'b011111100001;
   18185: result <= 12'b011111100001;
   18186: result <= 12'b011111100001;
   18187: result <= 12'b011111100001;
   18188: result <= 12'b011111100001;
   18189: result <= 12'b011111100001;
   18190: result <= 12'b011111100001;
   18191: result <= 12'b011111100001;
   18192: result <= 12'b011111100001;
   18193: result <= 12'b011111100001;
   18194: result <= 12'b011111100001;
   18195: result <= 12'b011111100001;
   18196: result <= 12'b011111100001;
   18197: result <= 12'b011111100001;
   18198: result <= 12'b011111100001;
   18199: result <= 12'b011111100001;
   18200: result <= 12'b011111100001;
   18201: result <= 12'b011111100001;
   18202: result <= 12'b011111100000;
   18203: result <= 12'b011111100000;
   18204: result <= 12'b011111100000;
   18205: result <= 12'b011111100000;
   18206: result <= 12'b011111100000;
   18207: result <= 12'b011111100000;
   18208: result <= 12'b011111100000;
   18209: result <= 12'b011111100000;
   18210: result <= 12'b011111100000;
   18211: result <= 12'b011111100000;
   18212: result <= 12'b011111100000;
   18213: result <= 12'b011111100000;
   18214: result <= 12'b011111100000;
   18215: result <= 12'b011111100000;
   18216: result <= 12'b011111100000;
   18217: result <= 12'b011111100000;
   18218: result <= 12'b011111100000;
   18219: result <= 12'b011111100000;
   18220: result <= 12'b011111100000;
   18221: result <= 12'b011111100000;
   18222: result <= 12'b011111100000;
   18223: result <= 12'b011111100000;
   18224: result <= 12'b011111100000;
   18225: result <= 12'b011111100000;
   18226: result <= 12'b011111100000;
   18227: result <= 12'b011111100000;
   18228: result <= 12'b011111100000;
   18229: result <= 12'b011111100000;
   18230: result <= 12'b011111100000;
   18231: result <= 12'b011111011111;
   18232: result <= 12'b011111011111;
   18233: result <= 12'b011111011111;
   18234: result <= 12'b011111011111;
   18235: result <= 12'b011111011111;
   18236: result <= 12'b011111011111;
   18237: result <= 12'b011111011111;
   18238: result <= 12'b011111011111;
   18239: result <= 12'b011111011111;
   18240: result <= 12'b011111011111;
   18241: result <= 12'b011111011111;
   18242: result <= 12'b011111011111;
   18243: result <= 12'b011111011111;
   18244: result <= 12'b011111011111;
   18245: result <= 12'b011111011111;
   18246: result <= 12'b011111011111;
   18247: result <= 12'b011111011111;
   18248: result <= 12'b011111011111;
   18249: result <= 12'b011111011111;
   18250: result <= 12'b011111011111;
   18251: result <= 12'b011111011111;
   18252: result <= 12'b011111011111;
   18253: result <= 12'b011111011111;
   18254: result <= 12'b011111011111;
   18255: result <= 12'b011111011111;
   18256: result <= 12'b011111011111;
   18257: result <= 12'b011111011111;
   18258: result <= 12'b011111011111;
   18259: result <= 12'b011111011110;
   18260: result <= 12'b011111011110;
   18261: result <= 12'b011111011110;
   18262: result <= 12'b011111011110;
   18263: result <= 12'b011111011110;
   18264: result <= 12'b011111011110;
   18265: result <= 12'b011111011110;
   18266: result <= 12'b011111011110;
   18267: result <= 12'b011111011110;
   18268: result <= 12'b011111011110;
   18269: result <= 12'b011111011110;
   18270: result <= 12'b011111011110;
   18271: result <= 12'b011111011110;
   18272: result <= 12'b011111011110;
   18273: result <= 12'b011111011110;
   18274: result <= 12'b011111011110;
   18275: result <= 12'b011111011110;
   18276: result <= 12'b011111011110;
   18277: result <= 12'b011111011110;
   18278: result <= 12'b011111011110;
   18279: result <= 12'b011111011110;
   18280: result <= 12'b011111011110;
   18281: result <= 12'b011111011110;
   18282: result <= 12'b011111011110;
   18283: result <= 12'b011111011110;
   18284: result <= 12'b011111011110;
   18285: result <= 12'b011111011110;
   18286: result <= 12'b011111011110;
   18287: result <= 12'b011111011110;
   18288: result <= 12'b011111011101;
   18289: result <= 12'b011111011101;
   18290: result <= 12'b011111011101;
   18291: result <= 12'b011111011101;
   18292: result <= 12'b011111011101;
   18293: result <= 12'b011111011101;
   18294: result <= 12'b011111011101;
   18295: result <= 12'b011111011101;
   18296: result <= 12'b011111011101;
   18297: result <= 12'b011111011101;
   18298: result <= 12'b011111011101;
   18299: result <= 12'b011111011101;
   18300: result <= 12'b011111011101;
   18301: result <= 12'b011111011101;
   18302: result <= 12'b011111011101;
   18303: result <= 12'b011111011101;
   18304: result <= 12'b011111011101;
   18305: result <= 12'b011111011101;
   18306: result <= 12'b011111011101;
   18307: result <= 12'b011111011101;
   18308: result <= 12'b011111011101;
   18309: result <= 12'b011111011101;
   18310: result <= 12'b011111011101;
   18311: result <= 12'b011111011101;
   18312: result <= 12'b011111011101;
   18313: result <= 12'b011111011101;
   18314: result <= 12'b011111011101;
   18315: result <= 12'b011111011101;
   18316: result <= 12'b011111011100;
   18317: result <= 12'b011111011100;
   18318: result <= 12'b011111011100;
   18319: result <= 12'b011111011100;
   18320: result <= 12'b011111011100;
   18321: result <= 12'b011111011100;
   18322: result <= 12'b011111011100;
   18323: result <= 12'b011111011100;
   18324: result <= 12'b011111011100;
   18325: result <= 12'b011111011100;
   18326: result <= 12'b011111011100;
   18327: result <= 12'b011111011100;
   18328: result <= 12'b011111011100;
   18329: result <= 12'b011111011100;
   18330: result <= 12'b011111011100;
   18331: result <= 12'b011111011100;
   18332: result <= 12'b011111011100;
   18333: result <= 12'b011111011100;
   18334: result <= 12'b011111011100;
   18335: result <= 12'b011111011100;
   18336: result <= 12'b011111011100;
   18337: result <= 12'b011111011100;
   18338: result <= 12'b011111011100;
   18339: result <= 12'b011111011100;
   18340: result <= 12'b011111011100;
   18341: result <= 12'b011111011100;
   18342: result <= 12'b011111011100;
   18343: result <= 12'b011111011011;
   18344: result <= 12'b011111011011;
   18345: result <= 12'b011111011011;
   18346: result <= 12'b011111011011;
   18347: result <= 12'b011111011011;
   18348: result <= 12'b011111011011;
   18349: result <= 12'b011111011011;
   18350: result <= 12'b011111011011;
   18351: result <= 12'b011111011011;
   18352: result <= 12'b011111011011;
   18353: result <= 12'b011111011011;
   18354: result <= 12'b011111011011;
   18355: result <= 12'b011111011011;
   18356: result <= 12'b011111011011;
   18357: result <= 12'b011111011011;
   18358: result <= 12'b011111011011;
   18359: result <= 12'b011111011011;
   18360: result <= 12'b011111011011;
   18361: result <= 12'b011111011011;
   18362: result <= 12'b011111011011;
   18363: result <= 12'b011111011011;
   18364: result <= 12'b011111011011;
   18365: result <= 12'b011111011011;
   18366: result <= 12'b011111011011;
   18367: result <= 12'b011111011011;
   18368: result <= 12'b011111011011;
   18369: result <= 12'b011111011011;
   18370: result <= 12'b011111011010;
   18371: result <= 12'b011111011010;
   18372: result <= 12'b011111011010;
   18373: result <= 12'b011111011010;
   18374: result <= 12'b011111011010;
   18375: result <= 12'b011111011010;
   18376: result <= 12'b011111011010;
   18377: result <= 12'b011111011010;
   18378: result <= 12'b011111011010;
   18379: result <= 12'b011111011010;
   18380: result <= 12'b011111011010;
   18381: result <= 12'b011111011010;
   18382: result <= 12'b011111011010;
   18383: result <= 12'b011111011010;
   18384: result <= 12'b011111011010;
   18385: result <= 12'b011111011010;
   18386: result <= 12'b011111011010;
   18387: result <= 12'b011111011010;
   18388: result <= 12'b011111011010;
   18389: result <= 12'b011111011010;
   18390: result <= 12'b011111011010;
   18391: result <= 12'b011111011010;
   18392: result <= 12'b011111011010;
   18393: result <= 12'b011111011010;
   18394: result <= 12'b011111011010;
   18395: result <= 12'b011111011010;
   18396: result <= 12'b011111011010;
   18397: result <= 12'b011111011001;
   18398: result <= 12'b011111011001;
   18399: result <= 12'b011111011001;
   18400: result <= 12'b011111011001;
   18401: result <= 12'b011111011001;
   18402: result <= 12'b011111011001;
   18403: result <= 12'b011111011001;
   18404: result <= 12'b011111011001;
   18405: result <= 12'b011111011001;
   18406: result <= 12'b011111011001;
   18407: result <= 12'b011111011001;
   18408: result <= 12'b011111011001;
   18409: result <= 12'b011111011001;
   18410: result <= 12'b011111011001;
   18411: result <= 12'b011111011001;
   18412: result <= 12'b011111011001;
   18413: result <= 12'b011111011001;
   18414: result <= 12'b011111011001;
   18415: result <= 12'b011111011001;
   18416: result <= 12'b011111011001;
   18417: result <= 12'b011111011001;
   18418: result <= 12'b011111011001;
   18419: result <= 12'b011111011001;
   18420: result <= 12'b011111011001;
   18421: result <= 12'b011111011001;
   18422: result <= 12'b011111011001;
   18423: result <= 12'b011111011000;
   18424: result <= 12'b011111011000;
   18425: result <= 12'b011111011000;
   18426: result <= 12'b011111011000;
   18427: result <= 12'b011111011000;
   18428: result <= 12'b011111011000;
   18429: result <= 12'b011111011000;
   18430: result <= 12'b011111011000;
   18431: result <= 12'b011111011000;
   18432: result <= 12'b011111011000;
   18433: result <= 12'b011111011000;
   18434: result <= 12'b011111011000;
   18435: result <= 12'b011111011000;
   18436: result <= 12'b011111011000;
   18437: result <= 12'b011111011000;
   18438: result <= 12'b011111011000;
   18439: result <= 12'b011111011000;
   18440: result <= 12'b011111011000;
   18441: result <= 12'b011111011000;
   18442: result <= 12'b011111011000;
   18443: result <= 12'b011111011000;
   18444: result <= 12'b011111011000;
   18445: result <= 12'b011111011000;
   18446: result <= 12'b011111011000;
   18447: result <= 12'b011111011000;
   18448: result <= 12'b011111011000;
   18449: result <= 12'b011111010111;
   18450: result <= 12'b011111010111;
   18451: result <= 12'b011111010111;
   18452: result <= 12'b011111010111;
   18453: result <= 12'b011111010111;
   18454: result <= 12'b011111010111;
   18455: result <= 12'b011111010111;
   18456: result <= 12'b011111010111;
   18457: result <= 12'b011111010111;
   18458: result <= 12'b011111010111;
   18459: result <= 12'b011111010111;
   18460: result <= 12'b011111010111;
   18461: result <= 12'b011111010111;
   18462: result <= 12'b011111010111;
   18463: result <= 12'b011111010111;
   18464: result <= 12'b011111010111;
   18465: result <= 12'b011111010111;
   18466: result <= 12'b011111010111;
   18467: result <= 12'b011111010111;
   18468: result <= 12'b011111010111;
   18469: result <= 12'b011111010111;
   18470: result <= 12'b011111010111;
   18471: result <= 12'b011111010111;
   18472: result <= 12'b011111010111;
   18473: result <= 12'b011111010111;
   18474: result <= 12'b011111010111;
   18475: result <= 12'b011111010110;
   18476: result <= 12'b011111010110;
   18477: result <= 12'b011111010110;
   18478: result <= 12'b011111010110;
   18479: result <= 12'b011111010110;
   18480: result <= 12'b011111010110;
   18481: result <= 12'b011111010110;
   18482: result <= 12'b011111010110;
   18483: result <= 12'b011111010110;
   18484: result <= 12'b011111010110;
   18485: result <= 12'b011111010110;
   18486: result <= 12'b011111010110;
   18487: result <= 12'b011111010110;
   18488: result <= 12'b011111010110;
   18489: result <= 12'b011111010110;
   18490: result <= 12'b011111010110;
   18491: result <= 12'b011111010110;
   18492: result <= 12'b011111010110;
   18493: result <= 12'b011111010110;
   18494: result <= 12'b011111010110;
   18495: result <= 12'b011111010110;
   18496: result <= 12'b011111010110;
   18497: result <= 12'b011111010110;
   18498: result <= 12'b011111010110;
   18499: result <= 12'b011111010110;
   18500: result <= 12'b011111010110;
   18501: result <= 12'b011111010101;
   18502: result <= 12'b011111010101;
   18503: result <= 12'b011111010101;
   18504: result <= 12'b011111010101;
   18505: result <= 12'b011111010101;
   18506: result <= 12'b011111010101;
   18507: result <= 12'b011111010101;
   18508: result <= 12'b011111010101;
   18509: result <= 12'b011111010101;
   18510: result <= 12'b011111010101;
   18511: result <= 12'b011111010101;
   18512: result <= 12'b011111010101;
   18513: result <= 12'b011111010101;
   18514: result <= 12'b011111010101;
   18515: result <= 12'b011111010101;
   18516: result <= 12'b011111010101;
   18517: result <= 12'b011111010101;
   18518: result <= 12'b011111010101;
   18519: result <= 12'b011111010101;
   18520: result <= 12'b011111010101;
   18521: result <= 12'b011111010101;
   18522: result <= 12'b011111010101;
   18523: result <= 12'b011111010101;
   18524: result <= 12'b011111010101;
   18525: result <= 12'b011111010101;
   18526: result <= 12'b011111010100;
   18527: result <= 12'b011111010100;
   18528: result <= 12'b011111010100;
   18529: result <= 12'b011111010100;
   18530: result <= 12'b011111010100;
   18531: result <= 12'b011111010100;
   18532: result <= 12'b011111010100;
   18533: result <= 12'b011111010100;
   18534: result <= 12'b011111010100;
   18535: result <= 12'b011111010100;
   18536: result <= 12'b011111010100;
   18537: result <= 12'b011111010100;
   18538: result <= 12'b011111010100;
   18539: result <= 12'b011111010100;
   18540: result <= 12'b011111010100;
   18541: result <= 12'b011111010100;
   18542: result <= 12'b011111010100;
   18543: result <= 12'b011111010100;
   18544: result <= 12'b011111010100;
   18545: result <= 12'b011111010100;
   18546: result <= 12'b011111010100;
   18547: result <= 12'b011111010100;
   18548: result <= 12'b011111010100;
   18549: result <= 12'b011111010100;
   18550: result <= 12'b011111010011;
   18551: result <= 12'b011111010011;
   18552: result <= 12'b011111010011;
   18553: result <= 12'b011111010011;
   18554: result <= 12'b011111010011;
   18555: result <= 12'b011111010011;
   18556: result <= 12'b011111010011;
   18557: result <= 12'b011111010011;
   18558: result <= 12'b011111010011;
   18559: result <= 12'b011111010011;
   18560: result <= 12'b011111010011;
   18561: result <= 12'b011111010011;
   18562: result <= 12'b011111010011;
   18563: result <= 12'b011111010011;
   18564: result <= 12'b011111010011;
   18565: result <= 12'b011111010011;
   18566: result <= 12'b011111010011;
   18567: result <= 12'b011111010011;
   18568: result <= 12'b011111010011;
   18569: result <= 12'b011111010011;
   18570: result <= 12'b011111010011;
   18571: result <= 12'b011111010011;
   18572: result <= 12'b011111010011;
   18573: result <= 12'b011111010011;
   18574: result <= 12'b011111010011;
   18575: result <= 12'b011111010010;
   18576: result <= 12'b011111010010;
   18577: result <= 12'b011111010010;
   18578: result <= 12'b011111010010;
   18579: result <= 12'b011111010010;
   18580: result <= 12'b011111010010;
   18581: result <= 12'b011111010010;
   18582: result <= 12'b011111010010;
   18583: result <= 12'b011111010010;
   18584: result <= 12'b011111010010;
   18585: result <= 12'b011111010010;
   18586: result <= 12'b011111010010;
   18587: result <= 12'b011111010010;
   18588: result <= 12'b011111010010;
   18589: result <= 12'b011111010010;
   18590: result <= 12'b011111010010;
   18591: result <= 12'b011111010010;
   18592: result <= 12'b011111010010;
   18593: result <= 12'b011111010010;
   18594: result <= 12'b011111010010;
   18595: result <= 12'b011111010010;
   18596: result <= 12'b011111010010;
   18597: result <= 12'b011111010010;
   18598: result <= 12'b011111010010;
   18599: result <= 12'b011111010001;
   18600: result <= 12'b011111010001;
   18601: result <= 12'b011111010001;
   18602: result <= 12'b011111010001;
   18603: result <= 12'b011111010001;
   18604: result <= 12'b011111010001;
   18605: result <= 12'b011111010001;
   18606: result <= 12'b011111010001;
   18607: result <= 12'b011111010001;
   18608: result <= 12'b011111010001;
   18609: result <= 12'b011111010001;
   18610: result <= 12'b011111010001;
   18611: result <= 12'b011111010001;
   18612: result <= 12'b011111010001;
   18613: result <= 12'b011111010001;
   18614: result <= 12'b011111010001;
   18615: result <= 12'b011111010001;
   18616: result <= 12'b011111010001;
   18617: result <= 12'b011111010001;
   18618: result <= 12'b011111010001;
   18619: result <= 12'b011111010001;
   18620: result <= 12'b011111010001;
   18621: result <= 12'b011111010001;
   18622: result <= 12'b011111010001;
   18623: result <= 12'b011111010000;
   18624: result <= 12'b011111010000;
   18625: result <= 12'b011111010000;
   18626: result <= 12'b011111010000;
   18627: result <= 12'b011111010000;
   18628: result <= 12'b011111010000;
   18629: result <= 12'b011111010000;
   18630: result <= 12'b011111010000;
   18631: result <= 12'b011111010000;
   18632: result <= 12'b011111010000;
   18633: result <= 12'b011111010000;
   18634: result <= 12'b011111010000;
   18635: result <= 12'b011111010000;
   18636: result <= 12'b011111010000;
   18637: result <= 12'b011111010000;
   18638: result <= 12'b011111010000;
   18639: result <= 12'b011111010000;
   18640: result <= 12'b011111010000;
   18641: result <= 12'b011111010000;
   18642: result <= 12'b011111010000;
   18643: result <= 12'b011111010000;
   18644: result <= 12'b011111010000;
   18645: result <= 12'b011111010000;
   18646: result <= 12'b011111010000;
   18647: result <= 12'b011111001111;
   18648: result <= 12'b011111001111;
   18649: result <= 12'b011111001111;
   18650: result <= 12'b011111001111;
   18651: result <= 12'b011111001111;
   18652: result <= 12'b011111001111;
   18653: result <= 12'b011111001111;
   18654: result <= 12'b011111001111;
   18655: result <= 12'b011111001111;
   18656: result <= 12'b011111001111;
   18657: result <= 12'b011111001111;
   18658: result <= 12'b011111001111;
   18659: result <= 12'b011111001111;
   18660: result <= 12'b011111001111;
   18661: result <= 12'b011111001111;
   18662: result <= 12'b011111001111;
   18663: result <= 12'b011111001111;
   18664: result <= 12'b011111001111;
   18665: result <= 12'b011111001111;
   18666: result <= 12'b011111001111;
   18667: result <= 12'b011111001111;
   18668: result <= 12'b011111001111;
   18669: result <= 12'b011111001111;
   18670: result <= 12'b011111001111;
   18671: result <= 12'b011111001110;
   18672: result <= 12'b011111001110;
   18673: result <= 12'b011111001110;
   18674: result <= 12'b011111001110;
   18675: result <= 12'b011111001110;
   18676: result <= 12'b011111001110;
   18677: result <= 12'b011111001110;
   18678: result <= 12'b011111001110;
   18679: result <= 12'b011111001110;
   18680: result <= 12'b011111001110;
   18681: result <= 12'b011111001110;
   18682: result <= 12'b011111001110;
   18683: result <= 12'b011111001110;
   18684: result <= 12'b011111001110;
   18685: result <= 12'b011111001110;
   18686: result <= 12'b011111001110;
   18687: result <= 12'b011111001110;
   18688: result <= 12'b011111001110;
   18689: result <= 12'b011111001110;
   18690: result <= 12'b011111001110;
   18691: result <= 12'b011111001110;
   18692: result <= 12'b011111001110;
   18693: result <= 12'b011111001110;
   18694: result <= 12'b011111001101;
   18695: result <= 12'b011111001101;
   18696: result <= 12'b011111001101;
   18697: result <= 12'b011111001101;
   18698: result <= 12'b011111001101;
   18699: result <= 12'b011111001101;
   18700: result <= 12'b011111001101;
   18701: result <= 12'b011111001101;
   18702: result <= 12'b011111001101;
   18703: result <= 12'b011111001101;
   18704: result <= 12'b011111001101;
   18705: result <= 12'b011111001101;
   18706: result <= 12'b011111001101;
   18707: result <= 12'b011111001101;
   18708: result <= 12'b011111001101;
   18709: result <= 12'b011111001101;
   18710: result <= 12'b011111001101;
   18711: result <= 12'b011111001101;
   18712: result <= 12'b011111001101;
   18713: result <= 12'b011111001101;
   18714: result <= 12'b011111001101;
   18715: result <= 12'b011111001101;
   18716: result <= 12'b011111001101;
   18717: result <= 12'b011111001100;
   18718: result <= 12'b011111001100;
   18719: result <= 12'b011111001100;
   18720: result <= 12'b011111001100;
   18721: result <= 12'b011111001100;
   18722: result <= 12'b011111001100;
   18723: result <= 12'b011111001100;
   18724: result <= 12'b011111001100;
   18725: result <= 12'b011111001100;
   18726: result <= 12'b011111001100;
   18727: result <= 12'b011111001100;
   18728: result <= 12'b011111001100;
   18729: result <= 12'b011111001100;
   18730: result <= 12'b011111001100;
   18731: result <= 12'b011111001100;
   18732: result <= 12'b011111001100;
   18733: result <= 12'b011111001100;
   18734: result <= 12'b011111001100;
   18735: result <= 12'b011111001100;
   18736: result <= 12'b011111001100;
   18737: result <= 12'b011111001100;
   18738: result <= 12'b011111001100;
   18739: result <= 12'b011111001100;
   18740: result <= 12'b011111001011;
   18741: result <= 12'b011111001011;
   18742: result <= 12'b011111001011;
   18743: result <= 12'b011111001011;
   18744: result <= 12'b011111001011;
   18745: result <= 12'b011111001011;
   18746: result <= 12'b011111001011;
   18747: result <= 12'b011111001011;
   18748: result <= 12'b011111001011;
   18749: result <= 12'b011111001011;
   18750: result <= 12'b011111001011;
   18751: result <= 12'b011111001011;
   18752: result <= 12'b011111001011;
   18753: result <= 12'b011111001011;
   18754: result <= 12'b011111001011;
   18755: result <= 12'b011111001011;
   18756: result <= 12'b011111001011;
   18757: result <= 12'b011111001011;
   18758: result <= 12'b011111001011;
   18759: result <= 12'b011111001011;
   18760: result <= 12'b011111001011;
   18761: result <= 12'b011111001011;
   18762: result <= 12'b011111001011;
   18763: result <= 12'b011111001010;
   18764: result <= 12'b011111001010;
   18765: result <= 12'b011111001010;
   18766: result <= 12'b011111001010;
   18767: result <= 12'b011111001010;
   18768: result <= 12'b011111001010;
   18769: result <= 12'b011111001010;
   18770: result <= 12'b011111001010;
   18771: result <= 12'b011111001010;
   18772: result <= 12'b011111001010;
   18773: result <= 12'b011111001010;
   18774: result <= 12'b011111001010;
   18775: result <= 12'b011111001010;
   18776: result <= 12'b011111001010;
   18777: result <= 12'b011111001010;
   18778: result <= 12'b011111001010;
   18779: result <= 12'b011111001010;
   18780: result <= 12'b011111001010;
   18781: result <= 12'b011111001010;
   18782: result <= 12'b011111001010;
   18783: result <= 12'b011111001010;
   18784: result <= 12'b011111001010;
   18785: result <= 12'b011111001001;
   18786: result <= 12'b011111001001;
   18787: result <= 12'b011111001001;
   18788: result <= 12'b011111001001;
   18789: result <= 12'b011111001001;
   18790: result <= 12'b011111001001;
   18791: result <= 12'b011111001001;
   18792: result <= 12'b011111001001;
   18793: result <= 12'b011111001001;
   18794: result <= 12'b011111001001;
   18795: result <= 12'b011111001001;
   18796: result <= 12'b011111001001;
   18797: result <= 12'b011111001001;
   18798: result <= 12'b011111001001;
   18799: result <= 12'b011111001001;
   18800: result <= 12'b011111001001;
   18801: result <= 12'b011111001001;
   18802: result <= 12'b011111001001;
   18803: result <= 12'b011111001001;
   18804: result <= 12'b011111001001;
   18805: result <= 12'b011111001001;
   18806: result <= 12'b011111001001;
   18807: result <= 12'b011111001000;
   18808: result <= 12'b011111001000;
   18809: result <= 12'b011111001000;
   18810: result <= 12'b011111001000;
   18811: result <= 12'b011111001000;
   18812: result <= 12'b011111001000;
   18813: result <= 12'b011111001000;
   18814: result <= 12'b011111001000;
   18815: result <= 12'b011111001000;
   18816: result <= 12'b011111001000;
   18817: result <= 12'b011111001000;
   18818: result <= 12'b011111001000;
   18819: result <= 12'b011111001000;
   18820: result <= 12'b011111001000;
   18821: result <= 12'b011111001000;
   18822: result <= 12'b011111001000;
   18823: result <= 12'b011111001000;
   18824: result <= 12'b011111001000;
   18825: result <= 12'b011111001000;
   18826: result <= 12'b011111001000;
   18827: result <= 12'b011111001000;
   18828: result <= 12'b011111001000;
   18829: result <= 12'b011111000111;
   18830: result <= 12'b011111000111;
   18831: result <= 12'b011111000111;
   18832: result <= 12'b011111000111;
   18833: result <= 12'b011111000111;
   18834: result <= 12'b011111000111;
   18835: result <= 12'b011111000111;
   18836: result <= 12'b011111000111;
   18837: result <= 12'b011111000111;
   18838: result <= 12'b011111000111;
   18839: result <= 12'b011111000111;
   18840: result <= 12'b011111000111;
   18841: result <= 12'b011111000111;
   18842: result <= 12'b011111000111;
   18843: result <= 12'b011111000111;
   18844: result <= 12'b011111000111;
   18845: result <= 12'b011111000111;
   18846: result <= 12'b011111000111;
   18847: result <= 12'b011111000111;
   18848: result <= 12'b011111000111;
   18849: result <= 12'b011111000111;
   18850: result <= 12'b011111000111;
   18851: result <= 12'b011111000110;
   18852: result <= 12'b011111000110;
   18853: result <= 12'b011111000110;
   18854: result <= 12'b011111000110;
   18855: result <= 12'b011111000110;
   18856: result <= 12'b011111000110;
   18857: result <= 12'b011111000110;
   18858: result <= 12'b011111000110;
   18859: result <= 12'b011111000110;
   18860: result <= 12'b011111000110;
   18861: result <= 12'b011111000110;
   18862: result <= 12'b011111000110;
   18863: result <= 12'b011111000110;
   18864: result <= 12'b011111000110;
   18865: result <= 12'b011111000110;
   18866: result <= 12'b011111000110;
   18867: result <= 12'b011111000110;
   18868: result <= 12'b011111000110;
   18869: result <= 12'b011111000110;
   18870: result <= 12'b011111000110;
   18871: result <= 12'b011111000110;
   18872: result <= 12'b011111000110;
   18873: result <= 12'b011111000101;
   18874: result <= 12'b011111000101;
   18875: result <= 12'b011111000101;
   18876: result <= 12'b011111000101;
   18877: result <= 12'b011111000101;
   18878: result <= 12'b011111000101;
   18879: result <= 12'b011111000101;
   18880: result <= 12'b011111000101;
   18881: result <= 12'b011111000101;
   18882: result <= 12'b011111000101;
   18883: result <= 12'b011111000101;
   18884: result <= 12'b011111000101;
   18885: result <= 12'b011111000101;
   18886: result <= 12'b011111000101;
   18887: result <= 12'b011111000101;
   18888: result <= 12'b011111000101;
   18889: result <= 12'b011111000101;
   18890: result <= 12'b011111000101;
   18891: result <= 12'b011111000101;
   18892: result <= 12'b011111000101;
   18893: result <= 12'b011111000101;
   18894: result <= 12'b011111000100;
   18895: result <= 12'b011111000100;
   18896: result <= 12'b011111000100;
   18897: result <= 12'b011111000100;
   18898: result <= 12'b011111000100;
   18899: result <= 12'b011111000100;
   18900: result <= 12'b011111000100;
   18901: result <= 12'b011111000100;
   18902: result <= 12'b011111000100;
   18903: result <= 12'b011111000100;
   18904: result <= 12'b011111000100;
   18905: result <= 12'b011111000100;
   18906: result <= 12'b011111000100;
   18907: result <= 12'b011111000100;
   18908: result <= 12'b011111000100;
   18909: result <= 12'b011111000100;
   18910: result <= 12'b011111000100;
   18911: result <= 12'b011111000100;
   18912: result <= 12'b011111000100;
   18913: result <= 12'b011111000100;
   18914: result <= 12'b011111000100;
   18915: result <= 12'b011111000011;
   18916: result <= 12'b011111000011;
   18917: result <= 12'b011111000011;
   18918: result <= 12'b011111000011;
   18919: result <= 12'b011111000011;
   18920: result <= 12'b011111000011;
   18921: result <= 12'b011111000011;
   18922: result <= 12'b011111000011;
   18923: result <= 12'b011111000011;
   18924: result <= 12'b011111000011;
   18925: result <= 12'b011111000011;
   18926: result <= 12'b011111000011;
   18927: result <= 12'b011111000011;
   18928: result <= 12'b011111000011;
   18929: result <= 12'b011111000011;
   18930: result <= 12'b011111000011;
   18931: result <= 12'b011111000011;
   18932: result <= 12'b011111000011;
   18933: result <= 12'b011111000011;
   18934: result <= 12'b011111000011;
   18935: result <= 12'b011111000011;
   18936: result <= 12'b011111000011;
   18937: result <= 12'b011111000010;
   18938: result <= 12'b011111000010;
   18939: result <= 12'b011111000010;
   18940: result <= 12'b011111000010;
   18941: result <= 12'b011111000010;
   18942: result <= 12'b011111000010;
   18943: result <= 12'b011111000010;
   18944: result <= 12'b011111000010;
   18945: result <= 12'b011111000010;
   18946: result <= 12'b011111000010;
   18947: result <= 12'b011111000010;
   18948: result <= 12'b011111000010;
   18949: result <= 12'b011111000010;
   18950: result <= 12'b011111000010;
   18951: result <= 12'b011111000010;
   18952: result <= 12'b011111000010;
   18953: result <= 12'b011111000010;
   18954: result <= 12'b011111000010;
   18955: result <= 12'b011111000010;
   18956: result <= 12'b011111000010;
   18957: result <= 12'b011111000010;
   18958: result <= 12'b011111000001;
   18959: result <= 12'b011111000001;
   18960: result <= 12'b011111000001;
   18961: result <= 12'b011111000001;
   18962: result <= 12'b011111000001;
   18963: result <= 12'b011111000001;
   18964: result <= 12'b011111000001;
   18965: result <= 12'b011111000001;
   18966: result <= 12'b011111000001;
   18967: result <= 12'b011111000001;
   18968: result <= 12'b011111000001;
   18969: result <= 12'b011111000001;
   18970: result <= 12'b011111000001;
   18971: result <= 12'b011111000001;
   18972: result <= 12'b011111000001;
   18973: result <= 12'b011111000001;
   18974: result <= 12'b011111000001;
   18975: result <= 12'b011111000001;
   18976: result <= 12'b011111000001;
   18977: result <= 12'b011111000001;
   18978: result <= 12'b011111000000;
   18979: result <= 12'b011111000000;
   18980: result <= 12'b011111000000;
   18981: result <= 12'b011111000000;
   18982: result <= 12'b011111000000;
   18983: result <= 12'b011111000000;
   18984: result <= 12'b011111000000;
   18985: result <= 12'b011111000000;
   18986: result <= 12'b011111000000;
   18987: result <= 12'b011111000000;
   18988: result <= 12'b011111000000;
   18989: result <= 12'b011111000000;
   18990: result <= 12'b011111000000;
   18991: result <= 12'b011111000000;
   18992: result <= 12'b011111000000;
   18993: result <= 12'b011111000000;
   18994: result <= 12'b011111000000;
   18995: result <= 12'b011111000000;
   18996: result <= 12'b011111000000;
   18997: result <= 12'b011111000000;
   18998: result <= 12'b011111000000;
   18999: result <= 12'b011110111111;
   19000: result <= 12'b011110111111;
   19001: result <= 12'b011110111111;
   19002: result <= 12'b011110111111;
   19003: result <= 12'b011110111111;
   19004: result <= 12'b011110111111;
   19005: result <= 12'b011110111111;
   19006: result <= 12'b011110111111;
   19007: result <= 12'b011110111111;
   19008: result <= 12'b011110111111;
   19009: result <= 12'b011110111111;
   19010: result <= 12'b011110111111;
   19011: result <= 12'b011110111111;
   19012: result <= 12'b011110111111;
   19013: result <= 12'b011110111111;
   19014: result <= 12'b011110111111;
   19015: result <= 12'b011110111111;
   19016: result <= 12'b011110111111;
   19017: result <= 12'b011110111111;
   19018: result <= 12'b011110111111;
   19019: result <= 12'b011110111110;
   19020: result <= 12'b011110111110;
   19021: result <= 12'b011110111110;
   19022: result <= 12'b011110111110;
   19023: result <= 12'b011110111110;
   19024: result <= 12'b011110111110;
   19025: result <= 12'b011110111110;
   19026: result <= 12'b011110111110;
   19027: result <= 12'b011110111110;
   19028: result <= 12'b011110111110;
   19029: result <= 12'b011110111110;
   19030: result <= 12'b011110111110;
   19031: result <= 12'b011110111110;
   19032: result <= 12'b011110111110;
   19033: result <= 12'b011110111110;
   19034: result <= 12'b011110111110;
   19035: result <= 12'b011110111110;
   19036: result <= 12'b011110111110;
   19037: result <= 12'b011110111110;
   19038: result <= 12'b011110111110;
   19039: result <= 12'b011110111110;
   19040: result <= 12'b011110111101;
   19041: result <= 12'b011110111101;
   19042: result <= 12'b011110111101;
   19043: result <= 12'b011110111101;
   19044: result <= 12'b011110111101;
   19045: result <= 12'b011110111101;
   19046: result <= 12'b011110111101;
   19047: result <= 12'b011110111101;
   19048: result <= 12'b011110111101;
   19049: result <= 12'b011110111101;
   19050: result <= 12'b011110111101;
   19051: result <= 12'b011110111101;
   19052: result <= 12'b011110111101;
   19053: result <= 12'b011110111101;
   19054: result <= 12'b011110111101;
   19055: result <= 12'b011110111101;
   19056: result <= 12'b011110111101;
   19057: result <= 12'b011110111101;
   19058: result <= 12'b011110111101;
   19059: result <= 12'b011110111101;
   19060: result <= 12'b011110111100;
   19061: result <= 12'b011110111100;
   19062: result <= 12'b011110111100;
   19063: result <= 12'b011110111100;
   19064: result <= 12'b011110111100;
   19065: result <= 12'b011110111100;
   19066: result <= 12'b011110111100;
   19067: result <= 12'b011110111100;
   19068: result <= 12'b011110111100;
   19069: result <= 12'b011110111100;
   19070: result <= 12'b011110111100;
   19071: result <= 12'b011110111100;
   19072: result <= 12'b011110111100;
   19073: result <= 12'b011110111100;
   19074: result <= 12'b011110111100;
   19075: result <= 12'b011110111100;
   19076: result <= 12'b011110111100;
   19077: result <= 12'b011110111100;
   19078: result <= 12'b011110111100;
   19079: result <= 12'b011110111100;
   19080: result <= 12'b011110111011;
   19081: result <= 12'b011110111011;
   19082: result <= 12'b011110111011;
   19083: result <= 12'b011110111011;
   19084: result <= 12'b011110111011;
   19085: result <= 12'b011110111011;
   19086: result <= 12'b011110111011;
   19087: result <= 12'b011110111011;
   19088: result <= 12'b011110111011;
   19089: result <= 12'b011110111011;
   19090: result <= 12'b011110111011;
   19091: result <= 12'b011110111011;
   19092: result <= 12'b011110111011;
   19093: result <= 12'b011110111011;
   19094: result <= 12'b011110111011;
   19095: result <= 12'b011110111011;
   19096: result <= 12'b011110111011;
   19097: result <= 12'b011110111011;
   19098: result <= 12'b011110111011;
   19099: result <= 12'b011110111011;
   19100: result <= 12'b011110111010;
   19101: result <= 12'b011110111010;
   19102: result <= 12'b011110111010;
   19103: result <= 12'b011110111010;
   19104: result <= 12'b011110111010;
   19105: result <= 12'b011110111010;
   19106: result <= 12'b011110111010;
   19107: result <= 12'b011110111010;
   19108: result <= 12'b011110111010;
   19109: result <= 12'b011110111010;
   19110: result <= 12'b011110111010;
   19111: result <= 12'b011110111010;
   19112: result <= 12'b011110111010;
   19113: result <= 12'b011110111010;
   19114: result <= 12'b011110111010;
   19115: result <= 12'b011110111010;
   19116: result <= 12'b011110111010;
   19117: result <= 12'b011110111010;
   19118: result <= 12'b011110111010;
   19119: result <= 12'b011110111001;
   19120: result <= 12'b011110111001;
   19121: result <= 12'b011110111001;
   19122: result <= 12'b011110111001;
   19123: result <= 12'b011110111001;
   19124: result <= 12'b011110111001;
   19125: result <= 12'b011110111001;
   19126: result <= 12'b011110111001;
   19127: result <= 12'b011110111001;
   19128: result <= 12'b011110111001;
   19129: result <= 12'b011110111001;
   19130: result <= 12'b011110111001;
   19131: result <= 12'b011110111001;
   19132: result <= 12'b011110111001;
   19133: result <= 12'b011110111001;
   19134: result <= 12'b011110111001;
   19135: result <= 12'b011110111001;
   19136: result <= 12'b011110111001;
   19137: result <= 12'b011110111001;
   19138: result <= 12'b011110111001;
   19139: result <= 12'b011110111000;
   19140: result <= 12'b011110111000;
   19141: result <= 12'b011110111000;
   19142: result <= 12'b011110111000;
   19143: result <= 12'b011110111000;
   19144: result <= 12'b011110111000;
   19145: result <= 12'b011110111000;
   19146: result <= 12'b011110111000;
   19147: result <= 12'b011110111000;
   19148: result <= 12'b011110111000;
   19149: result <= 12'b011110111000;
   19150: result <= 12'b011110111000;
   19151: result <= 12'b011110111000;
   19152: result <= 12'b011110111000;
   19153: result <= 12'b011110111000;
   19154: result <= 12'b011110111000;
   19155: result <= 12'b011110111000;
   19156: result <= 12'b011110111000;
   19157: result <= 12'b011110111000;
   19158: result <= 12'b011110110111;
   19159: result <= 12'b011110110111;
   19160: result <= 12'b011110110111;
   19161: result <= 12'b011110110111;
   19162: result <= 12'b011110110111;
   19163: result <= 12'b011110110111;
   19164: result <= 12'b011110110111;
   19165: result <= 12'b011110110111;
   19166: result <= 12'b011110110111;
   19167: result <= 12'b011110110111;
   19168: result <= 12'b011110110111;
   19169: result <= 12'b011110110111;
   19170: result <= 12'b011110110111;
   19171: result <= 12'b011110110111;
   19172: result <= 12'b011110110111;
   19173: result <= 12'b011110110111;
   19174: result <= 12'b011110110111;
   19175: result <= 12'b011110110111;
   19176: result <= 12'b011110110111;
   19177: result <= 12'b011110110111;
   19178: result <= 12'b011110110110;
   19179: result <= 12'b011110110110;
   19180: result <= 12'b011110110110;
   19181: result <= 12'b011110110110;
   19182: result <= 12'b011110110110;
   19183: result <= 12'b011110110110;
   19184: result <= 12'b011110110110;
   19185: result <= 12'b011110110110;
   19186: result <= 12'b011110110110;
   19187: result <= 12'b011110110110;
   19188: result <= 12'b011110110110;
   19189: result <= 12'b011110110110;
   19190: result <= 12'b011110110110;
   19191: result <= 12'b011110110110;
   19192: result <= 12'b011110110110;
   19193: result <= 12'b011110110110;
   19194: result <= 12'b011110110110;
   19195: result <= 12'b011110110110;
   19196: result <= 12'b011110110110;
   19197: result <= 12'b011110110101;
   19198: result <= 12'b011110110101;
   19199: result <= 12'b011110110101;
   19200: result <= 12'b011110110101;
   19201: result <= 12'b011110110101;
   19202: result <= 12'b011110110101;
   19203: result <= 12'b011110110101;
   19204: result <= 12'b011110110101;
   19205: result <= 12'b011110110101;
   19206: result <= 12'b011110110101;
   19207: result <= 12'b011110110101;
   19208: result <= 12'b011110110101;
   19209: result <= 12'b011110110101;
   19210: result <= 12'b011110110101;
   19211: result <= 12'b011110110101;
   19212: result <= 12'b011110110101;
   19213: result <= 12'b011110110101;
   19214: result <= 12'b011110110101;
   19215: result <= 12'b011110110101;
   19216: result <= 12'b011110110100;
   19217: result <= 12'b011110110100;
   19218: result <= 12'b011110110100;
   19219: result <= 12'b011110110100;
   19220: result <= 12'b011110110100;
   19221: result <= 12'b011110110100;
   19222: result <= 12'b011110110100;
   19223: result <= 12'b011110110100;
   19224: result <= 12'b011110110100;
   19225: result <= 12'b011110110100;
   19226: result <= 12'b011110110100;
   19227: result <= 12'b011110110100;
   19228: result <= 12'b011110110100;
   19229: result <= 12'b011110110100;
   19230: result <= 12'b011110110100;
   19231: result <= 12'b011110110100;
   19232: result <= 12'b011110110100;
   19233: result <= 12'b011110110100;
   19234: result <= 12'b011110110100;
   19235: result <= 12'b011110110011;
   19236: result <= 12'b011110110011;
   19237: result <= 12'b011110110011;
   19238: result <= 12'b011110110011;
   19239: result <= 12'b011110110011;
   19240: result <= 12'b011110110011;
   19241: result <= 12'b011110110011;
   19242: result <= 12'b011110110011;
   19243: result <= 12'b011110110011;
   19244: result <= 12'b011110110011;
   19245: result <= 12'b011110110011;
   19246: result <= 12'b011110110011;
   19247: result <= 12'b011110110011;
   19248: result <= 12'b011110110011;
   19249: result <= 12'b011110110011;
   19250: result <= 12'b011110110011;
   19251: result <= 12'b011110110011;
   19252: result <= 12'b011110110011;
   19253: result <= 12'b011110110011;
   19254: result <= 12'b011110110010;
   19255: result <= 12'b011110110010;
   19256: result <= 12'b011110110010;
   19257: result <= 12'b011110110010;
   19258: result <= 12'b011110110010;
   19259: result <= 12'b011110110010;
   19260: result <= 12'b011110110010;
   19261: result <= 12'b011110110010;
   19262: result <= 12'b011110110010;
   19263: result <= 12'b011110110010;
   19264: result <= 12'b011110110010;
   19265: result <= 12'b011110110010;
   19266: result <= 12'b011110110010;
   19267: result <= 12'b011110110010;
   19268: result <= 12'b011110110010;
   19269: result <= 12'b011110110010;
   19270: result <= 12'b011110110010;
   19271: result <= 12'b011110110010;
   19272: result <= 12'b011110110001;
   19273: result <= 12'b011110110001;
   19274: result <= 12'b011110110001;
   19275: result <= 12'b011110110001;
   19276: result <= 12'b011110110001;
   19277: result <= 12'b011110110001;
   19278: result <= 12'b011110110001;
   19279: result <= 12'b011110110001;
   19280: result <= 12'b011110110001;
   19281: result <= 12'b011110110001;
   19282: result <= 12'b011110110001;
   19283: result <= 12'b011110110001;
   19284: result <= 12'b011110110001;
   19285: result <= 12'b011110110001;
   19286: result <= 12'b011110110001;
   19287: result <= 12'b011110110001;
   19288: result <= 12'b011110110001;
   19289: result <= 12'b011110110001;
   19290: result <= 12'b011110110001;
   19291: result <= 12'b011110110000;
   19292: result <= 12'b011110110000;
   19293: result <= 12'b011110110000;
   19294: result <= 12'b011110110000;
   19295: result <= 12'b011110110000;
   19296: result <= 12'b011110110000;
   19297: result <= 12'b011110110000;
   19298: result <= 12'b011110110000;
   19299: result <= 12'b011110110000;
   19300: result <= 12'b011110110000;
   19301: result <= 12'b011110110000;
   19302: result <= 12'b011110110000;
   19303: result <= 12'b011110110000;
   19304: result <= 12'b011110110000;
   19305: result <= 12'b011110110000;
   19306: result <= 12'b011110110000;
   19307: result <= 12'b011110110000;
   19308: result <= 12'b011110110000;
   19309: result <= 12'b011110101111;
   19310: result <= 12'b011110101111;
   19311: result <= 12'b011110101111;
   19312: result <= 12'b011110101111;
   19313: result <= 12'b011110101111;
   19314: result <= 12'b011110101111;
   19315: result <= 12'b011110101111;
   19316: result <= 12'b011110101111;
   19317: result <= 12'b011110101111;
   19318: result <= 12'b011110101111;
   19319: result <= 12'b011110101111;
   19320: result <= 12'b011110101111;
   19321: result <= 12'b011110101111;
   19322: result <= 12'b011110101111;
   19323: result <= 12'b011110101111;
   19324: result <= 12'b011110101111;
   19325: result <= 12'b011110101111;
   19326: result <= 12'b011110101111;
   19327: result <= 12'b011110101111;
   19328: result <= 12'b011110101110;
   19329: result <= 12'b011110101110;
   19330: result <= 12'b011110101110;
   19331: result <= 12'b011110101110;
   19332: result <= 12'b011110101110;
   19333: result <= 12'b011110101110;
   19334: result <= 12'b011110101110;
   19335: result <= 12'b011110101110;
   19336: result <= 12'b011110101110;
   19337: result <= 12'b011110101110;
   19338: result <= 12'b011110101110;
   19339: result <= 12'b011110101110;
   19340: result <= 12'b011110101110;
   19341: result <= 12'b011110101110;
   19342: result <= 12'b011110101110;
   19343: result <= 12'b011110101110;
   19344: result <= 12'b011110101110;
   19345: result <= 12'b011110101110;
   19346: result <= 12'b011110101101;
   19347: result <= 12'b011110101101;
   19348: result <= 12'b011110101101;
   19349: result <= 12'b011110101101;
   19350: result <= 12'b011110101101;
   19351: result <= 12'b011110101101;
   19352: result <= 12'b011110101101;
   19353: result <= 12'b011110101101;
   19354: result <= 12'b011110101101;
   19355: result <= 12'b011110101101;
   19356: result <= 12'b011110101101;
   19357: result <= 12'b011110101101;
   19358: result <= 12'b011110101101;
   19359: result <= 12'b011110101101;
   19360: result <= 12'b011110101101;
   19361: result <= 12'b011110101101;
   19362: result <= 12'b011110101101;
   19363: result <= 12'b011110101101;
   19364: result <= 12'b011110101100;
   19365: result <= 12'b011110101100;
   19366: result <= 12'b011110101100;
   19367: result <= 12'b011110101100;
   19368: result <= 12'b011110101100;
   19369: result <= 12'b011110101100;
   19370: result <= 12'b011110101100;
   19371: result <= 12'b011110101100;
   19372: result <= 12'b011110101100;
   19373: result <= 12'b011110101100;
   19374: result <= 12'b011110101100;
   19375: result <= 12'b011110101100;
   19376: result <= 12'b011110101100;
   19377: result <= 12'b011110101100;
   19378: result <= 12'b011110101100;
   19379: result <= 12'b011110101100;
   19380: result <= 12'b011110101100;
   19381: result <= 12'b011110101100;
   19382: result <= 12'b011110101011;
   19383: result <= 12'b011110101011;
   19384: result <= 12'b011110101011;
   19385: result <= 12'b011110101011;
   19386: result <= 12'b011110101011;
   19387: result <= 12'b011110101011;
   19388: result <= 12'b011110101011;
   19389: result <= 12'b011110101011;
   19390: result <= 12'b011110101011;
   19391: result <= 12'b011110101011;
   19392: result <= 12'b011110101011;
   19393: result <= 12'b011110101011;
   19394: result <= 12'b011110101011;
   19395: result <= 12'b011110101011;
   19396: result <= 12'b011110101011;
   19397: result <= 12'b011110101011;
   19398: result <= 12'b011110101011;
   19399: result <= 12'b011110101011;
   19400: result <= 12'b011110101010;
   19401: result <= 12'b011110101010;
   19402: result <= 12'b011110101010;
   19403: result <= 12'b011110101010;
   19404: result <= 12'b011110101010;
   19405: result <= 12'b011110101010;
   19406: result <= 12'b011110101010;
   19407: result <= 12'b011110101010;
   19408: result <= 12'b011110101010;
   19409: result <= 12'b011110101010;
   19410: result <= 12'b011110101010;
   19411: result <= 12'b011110101010;
   19412: result <= 12'b011110101010;
   19413: result <= 12'b011110101010;
   19414: result <= 12'b011110101010;
   19415: result <= 12'b011110101010;
   19416: result <= 12'b011110101010;
   19417: result <= 12'b011110101010;
   19418: result <= 12'b011110101001;
   19419: result <= 12'b011110101001;
   19420: result <= 12'b011110101001;
   19421: result <= 12'b011110101001;
   19422: result <= 12'b011110101001;
   19423: result <= 12'b011110101001;
   19424: result <= 12'b011110101001;
   19425: result <= 12'b011110101001;
   19426: result <= 12'b011110101001;
   19427: result <= 12'b011110101001;
   19428: result <= 12'b011110101001;
   19429: result <= 12'b011110101001;
   19430: result <= 12'b011110101001;
   19431: result <= 12'b011110101001;
   19432: result <= 12'b011110101001;
   19433: result <= 12'b011110101001;
   19434: result <= 12'b011110101001;
   19435: result <= 12'b011110101001;
   19436: result <= 12'b011110101000;
   19437: result <= 12'b011110101000;
   19438: result <= 12'b011110101000;
   19439: result <= 12'b011110101000;
   19440: result <= 12'b011110101000;
   19441: result <= 12'b011110101000;
   19442: result <= 12'b011110101000;
   19443: result <= 12'b011110101000;
   19444: result <= 12'b011110101000;
   19445: result <= 12'b011110101000;
   19446: result <= 12'b011110101000;
   19447: result <= 12'b011110101000;
   19448: result <= 12'b011110101000;
   19449: result <= 12'b011110101000;
   19450: result <= 12'b011110101000;
   19451: result <= 12'b011110101000;
   19452: result <= 12'b011110101000;
   19453: result <= 12'b011110100111;
   19454: result <= 12'b011110100111;
   19455: result <= 12'b011110100111;
   19456: result <= 12'b011110100111;
   19457: result <= 12'b011110100111;
   19458: result <= 12'b011110100111;
   19459: result <= 12'b011110100111;
   19460: result <= 12'b011110100111;
   19461: result <= 12'b011110100111;
   19462: result <= 12'b011110100111;
   19463: result <= 12'b011110100111;
   19464: result <= 12'b011110100111;
   19465: result <= 12'b011110100111;
   19466: result <= 12'b011110100111;
   19467: result <= 12'b011110100111;
   19468: result <= 12'b011110100111;
   19469: result <= 12'b011110100111;
   19470: result <= 12'b011110100111;
   19471: result <= 12'b011110100110;
   19472: result <= 12'b011110100110;
   19473: result <= 12'b011110100110;
   19474: result <= 12'b011110100110;
   19475: result <= 12'b011110100110;
   19476: result <= 12'b011110100110;
   19477: result <= 12'b011110100110;
   19478: result <= 12'b011110100110;
   19479: result <= 12'b011110100110;
   19480: result <= 12'b011110100110;
   19481: result <= 12'b011110100110;
   19482: result <= 12'b011110100110;
   19483: result <= 12'b011110100110;
   19484: result <= 12'b011110100110;
   19485: result <= 12'b011110100110;
   19486: result <= 12'b011110100110;
   19487: result <= 12'b011110100110;
   19488: result <= 12'b011110100101;
   19489: result <= 12'b011110100101;
   19490: result <= 12'b011110100101;
   19491: result <= 12'b011110100101;
   19492: result <= 12'b011110100101;
   19493: result <= 12'b011110100101;
   19494: result <= 12'b011110100101;
   19495: result <= 12'b011110100101;
   19496: result <= 12'b011110100101;
   19497: result <= 12'b011110100101;
   19498: result <= 12'b011110100101;
   19499: result <= 12'b011110100101;
   19500: result <= 12'b011110100101;
   19501: result <= 12'b011110100101;
   19502: result <= 12'b011110100101;
   19503: result <= 12'b011110100101;
   19504: result <= 12'b011110100101;
   19505: result <= 12'b011110100100;
   19506: result <= 12'b011110100100;
   19507: result <= 12'b011110100100;
   19508: result <= 12'b011110100100;
   19509: result <= 12'b011110100100;
   19510: result <= 12'b011110100100;
   19511: result <= 12'b011110100100;
   19512: result <= 12'b011110100100;
   19513: result <= 12'b011110100100;
   19514: result <= 12'b011110100100;
   19515: result <= 12'b011110100100;
   19516: result <= 12'b011110100100;
   19517: result <= 12'b011110100100;
   19518: result <= 12'b011110100100;
   19519: result <= 12'b011110100100;
   19520: result <= 12'b011110100100;
   19521: result <= 12'b011110100100;
   19522: result <= 12'b011110100100;
   19523: result <= 12'b011110100011;
   19524: result <= 12'b011110100011;
   19525: result <= 12'b011110100011;
   19526: result <= 12'b011110100011;
   19527: result <= 12'b011110100011;
   19528: result <= 12'b011110100011;
   19529: result <= 12'b011110100011;
   19530: result <= 12'b011110100011;
   19531: result <= 12'b011110100011;
   19532: result <= 12'b011110100011;
   19533: result <= 12'b011110100011;
   19534: result <= 12'b011110100011;
   19535: result <= 12'b011110100011;
   19536: result <= 12'b011110100011;
   19537: result <= 12'b011110100011;
   19538: result <= 12'b011110100011;
   19539: result <= 12'b011110100011;
   19540: result <= 12'b011110100010;
   19541: result <= 12'b011110100010;
   19542: result <= 12'b011110100010;
   19543: result <= 12'b011110100010;
   19544: result <= 12'b011110100010;
   19545: result <= 12'b011110100010;
   19546: result <= 12'b011110100010;
   19547: result <= 12'b011110100010;
   19548: result <= 12'b011110100010;
   19549: result <= 12'b011110100010;
   19550: result <= 12'b011110100010;
   19551: result <= 12'b011110100010;
   19552: result <= 12'b011110100010;
   19553: result <= 12'b011110100010;
   19554: result <= 12'b011110100010;
   19555: result <= 12'b011110100010;
   19556: result <= 12'b011110100010;
   19557: result <= 12'b011110100001;
   19558: result <= 12'b011110100001;
   19559: result <= 12'b011110100001;
   19560: result <= 12'b011110100001;
   19561: result <= 12'b011110100001;
   19562: result <= 12'b011110100001;
   19563: result <= 12'b011110100001;
   19564: result <= 12'b011110100001;
   19565: result <= 12'b011110100001;
   19566: result <= 12'b011110100001;
   19567: result <= 12'b011110100001;
   19568: result <= 12'b011110100001;
   19569: result <= 12'b011110100001;
   19570: result <= 12'b011110100001;
   19571: result <= 12'b011110100001;
   19572: result <= 12'b011110100001;
   19573: result <= 12'b011110100001;
   19574: result <= 12'b011110100000;
   19575: result <= 12'b011110100000;
   19576: result <= 12'b011110100000;
   19577: result <= 12'b011110100000;
   19578: result <= 12'b011110100000;
   19579: result <= 12'b011110100000;
   19580: result <= 12'b011110100000;
   19581: result <= 12'b011110100000;
   19582: result <= 12'b011110100000;
   19583: result <= 12'b011110100000;
   19584: result <= 12'b011110100000;
   19585: result <= 12'b011110100000;
   19586: result <= 12'b011110100000;
   19587: result <= 12'b011110100000;
   19588: result <= 12'b011110100000;
   19589: result <= 12'b011110100000;
   19590: result <= 12'b011110100000;
   19591: result <= 12'b011110011111;
   19592: result <= 12'b011110011111;
   19593: result <= 12'b011110011111;
   19594: result <= 12'b011110011111;
   19595: result <= 12'b011110011111;
   19596: result <= 12'b011110011111;
   19597: result <= 12'b011110011111;
   19598: result <= 12'b011110011111;
   19599: result <= 12'b011110011111;
   19600: result <= 12'b011110011111;
   19601: result <= 12'b011110011111;
   19602: result <= 12'b011110011111;
   19603: result <= 12'b011110011111;
   19604: result <= 12'b011110011111;
   19605: result <= 12'b011110011111;
   19606: result <= 12'b011110011111;
   19607: result <= 12'b011110011111;
   19608: result <= 12'b011110011110;
   19609: result <= 12'b011110011110;
   19610: result <= 12'b011110011110;
   19611: result <= 12'b011110011110;
   19612: result <= 12'b011110011110;
   19613: result <= 12'b011110011110;
   19614: result <= 12'b011110011110;
   19615: result <= 12'b011110011110;
   19616: result <= 12'b011110011110;
   19617: result <= 12'b011110011110;
   19618: result <= 12'b011110011110;
   19619: result <= 12'b011110011110;
   19620: result <= 12'b011110011110;
   19621: result <= 12'b011110011110;
   19622: result <= 12'b011110011110;
   19623: result <= 12'b011110011110;
   19624: result <= 12'b011110011101;
   19625: result <= 12'b011110011101;
   19626: result <= 12'b011110011101;
   19627: result <= 12'b011110011101;
   19628: result <= 12'b011110011101;
   19629: result <= 12'b011110011101;
   19630: result <= 12'b011110011101;
   19631: result <= 12'b011110011101;
   19632: result <= 12'b011110011101;
   19633: result <= 12'b011110011101;
   19634: result <= 12'b011110011101;
   19635: result <= 12'b011110011101;
   19636: result <= 12'b011110011101;
   19637: result <= 12'b011110011101;
   19638: result <= 12'b011110011101;
   19639: result <= 12'b011110011101;
   19640: result <= 12'b011110011101;
   19641: result <= 12'b011110011100;
   19642: result <= 12'b011110011100;
   19643: result <= 12'b011110011100;
   19644: result <= 12'b011110011100;
   19645: result <= 12'b011110011100;
   19646: result <= 12'b011110011100;
   19647: result <= 12'b011110011100;
   19648: result <= 12'b011110011100;
   19649: result <= 12'b011110011100;
   19650: result <= 12'b011110011100;
   19651: result <= 12'b011110011100;
   19652: result <= 12'b011110011100;
   19653: result <= 12'b011110011100;
   19654: result <= 12'b011110011100;
   19655: result <= 12'b011110011100;
   19656: result <= 12'b011110011100;
   19657: result <= 12'b011110011011;
   19658: result <= 12'b011110011011;
   19659: result <= 12'b011110011011;
   19660: result <= 12'b011110011011;
   19661: result <= 12'b011110011011;
   19662: result <= 12'b011110011011;
   19663: result <= 12'b011110011011;
   19664: result <= 12'b011110011011;
   19665: result <= 12'b011110011011;
   19666: result <= 12'b011110011011;
   19667: result <= 12'b011110011011;
   19668: result <= 12'b011110011011;
   19669: result <= 12'b011110011011;
   19670: result <= 12'b011110011011;
   19671: result <= 12'b011110011011;
   19672: result <= 12'b011110011011;
   19673: result <= 12'b011110011011;
   19674: result <= 12'b011110011010;
   19675: result <= 12'b011110011010;
   19676: result <= 12'b011110011010;
   19677: result <= 12'b011110011010;
   19678: result <= 12'b011110011010;
   19679: result <= 12'b011110011010;
   19680: result <= 12'b011110011010;
   19681: result <= 12'b011110011010;
   19682: result <= 12'b011110011010;
   19683: result <= 12'b011110011010;
   19684: result <= 12'b011110011010;
   19685: result <= 12'b011110011010;
   19686: result <= 12'b011110011010;
   19687: result <= 12'b011110011010;
   19688: result <= 12'b011110011010;
   19689: result <= 12'b011110011010;
   19690: result <= 12'b011110011001;
   19691: result <= 12'b011110011001;
   19692: result <= 12'b011110011001;
   19693: result <= 12'b011110011001;
   19694: result <= 12'b011110011001;
   19695: result <= 12'b011110011001;
   19696: result <= 12'b011110011001;
   19697: result <= 12'b011110011001;
   19698: result <= 12'b011110011001;
   19699: result <= 12'b011110011001;
   19700: result <= 12'b011110011001;
   19701: result <= 12'b011110011001;
   19702: result <= 12'b011110011001;
   19703: result <= 12'b011110011001;
   19704: result <= 12'b011110011001;
   19705: result <= 12'b011110011001;
   19706: result <= 12'b011110011001;
   19707: result <= 12'b011110011000;
   19708: result <= 12'b011110011000;
   19709: result <= 12'b011110011000;
   19710: result <= 12'b011110011000;
   19711: result <= 12'b011110011000;
   19712: result <= 12'b011110011000;
   19713: result <= 12'b011110011000;
   19714: result <= 12'b011110011000;
   19715: result <= 12'b011110011000;
   19716: result <= 12'b011110011000;
   19717: result <= 12'b011110011000;
   19718: result <= 12'b011110011000;
   19719: result <= 12'b011110011000;
   19720: result <= 12'b011110011000;
   19721: result <= 12'b011110011000;
   19722: result <= 12'b011110011000;
   19723: result <= 12'b011110010111;
   19724: result <= 12'b011110010111;
   19725: result <= 12'b011110010111;
   19726: result <= 12'b011110010111;
   19727: result <= 12'b011110010111;
   19728: result <= 12'b011110010111;
   19729: result <= 12'b011110010111;
   19730: result <= 12'b011110010111;
   19731: result <= 12'b011110010111;
   19732: result <= 12'b011110010111;
   19733: result <= 12'b011110010111;
   19734: result <= 12'b011110010111;
   19735: result <= 12'b011110010111;
   19736: result <= 12'b011110010111;
   19737: result <= 12'b011110010111;
   19738: result <= 12'b011110010111;
   19739: result <= 12'b011110010110;
   19740: result <= 12'b011110010110;
   19741: result <= 12'b011110010110;
   19742: result <= 12'b011110010110;
   19743: result <= 12'b011110010110;
   19744: result <= 12'b011110010110;
   19745: result <= 12'b011110010110;
   19746: result <= 12'b011110010110;
   19747: result <= 12'b011110010110;
   19748: result <= 12'b011110010110;
   19749: result <= 12'b011110010110;
   19750: result <= 12'b011110010110;
   19751: result <= 12'b011110010110;
   19752: result <= 12'b011110010110;
   19753: result <= 12'b011110010110;
   19754: result <= 12'b011110010110;
   19755: result <= 12'b011110010101;
   19756: result <= 12'b011110010101;
   19757: result <= 12'b011110010101;
   19758: result <= 12'b011110010101;
   19759: result <= 12'b011110010101;
   19760: result <= 12'b011110010101;
   19761: result <= 12'b011110010101;
   19762: result <= 12'b011110010101;
   19763: result <= 12'b011110010101;
   19764: result <= 12'b011110010101;
   19765: result <= 12'b011110010101;
   19766: result <= 12'b011110010101;
   19767: result <= 12'b011110010101;
   19768: result <= 12'b011110010101;
   19769: result <= 12'b011110010101;
   19770: result <= 12'b011110010101;
   19771: result <= 12'b011110010100;
   19772: result <= 12'b011110010100;
   19773: result <= 12'b011110010100;
   19774: result <= 12'b011110010100;
   19775: result <= 12'b011110010100;
   19776: result <= 12'b011110010100;
   19777: result <= 12'b011110010100;
   19778: result <= 12'b011110010100;
   19779: result <= 12'b011110010100;
   19780: result <= 12'b011110010100;
   19781: result <= 12'b011110010100;
   19782: result <= 12'b011110010100;
   19783: result <= 12'b011110010100;
   19784: result <= 12'b011110010100;
   19785: result <= 12'b011110010100;
   19786: result <= 12'b011110010100;
   19787: result <= 12'b011110010011;
   19788: result <= 12'b011110010011;
   19789: result <= 12'b011110010011;
   19790: result <= 12'b011110010011;
   19791: result <= 12'b011110010011;
   19792: result <= 12'b011110010011;
   19793: result <= 12'b011110010011;
   19794: result <= 12'b011110010011;
   19795: result <= 12'b011110010011;
   19796: result <= 12'b011110010011;
   19797: result <= 12'b011110010011;
   19798: result <= 12'b011110010011;
   19799: result <= 12'b011110010011;
   19800: result <= 12'b011110010011;
   19801: result <= 12'b011110010011;
   19802: result <= 12'b011110010011;
   19803: result <= 12'b011110010010;
   19804: result <= 12'b011110010010;
   19805: result <= 12'b011110010010;
   19806: result <= 12'b011110010010;
   19807: result <= 12'b011110010010;
   19808: result <= 12'b011110010010;
   19809: result <= 12'b011110010010;
   19810: result <= 12'b011110010010;
   19811: result <= 12'b011110010010;
   19812: result <= 12'b011110010010;
   19813: result <= 12'b011110010010;
   19814: result <= 12'b011110010010;
   19815: result <= 12'b011110010010;
   19816: result <= 12'b011110010010;
   19817: result <= 12'b011110010010;
   19818: result <= 12'b011110010010;
   19819: result <= 12'b011110010001;
   19820: result <= 12'b011110010001;
   19821: result <= 12'b011110010001;
   19822: result <= 12'b011110010001;
   19823: result <= 12'b011110010001;
   19824: result <= 12'b011110010001;
   19825: result <= 12'b011110010001;
   19826: result <= 12'b011110010001;
   19827: result <= 12'b011110010001;
   19828: result <= 12'b011110010001;
   19829: result <= 12'b011110010001;
   19830: result <= 12'b011110010001;
   19831: result <= 12'b011110010001;
   19832: result <= 12'b011110010001;
   19833: result <= 12'b011110010001;
   19834: result <= 12'b011110010000;
   19835: result <= 12'b011110010000;
   19836: result <= 12'b011110010000;
   19837: result <= 12'b011110010000;
   19838: result <= 12'b011110010000;
   19839: result <= 12'b011110010000;
   19840: result <= 12'b011110010000;
   19841: result <= 12'b011110010000;
   19842: result <= 12'b011110010000;
   19843: result <= 12'b011110010000;
   19844: result <= 12'b011110010000;
   19845: result <= 12'b011110010000;
   19846: result <= 12'b011110010000;
   19847: result <= 12'b011110010000;
   19848: result <= 12'b011110010000;
   19849: result <= 12'b011110010000;
   19850: result <= 12'b011110001111;
   19851: result <= 12'b011110001111;
   19852: result <= 12'b011110001111;
   19853: result <= 12'b011110001111;
   19854: result <= 12'b011110001111;
   19855: result <= 12'b011110001111;
   19856: result <= 12'b011110001111;
   19857: result <= 12'b011110001111;
   19858: result <= 12'b011110001111;
   19859: result <= 12'b011110001111;
   19860: result <= 12'b011110001111;
   19861: result <= 12'b011110001111;
   19862: result <= 12'b011110001111;
   19863: result <= 12'b011110001111;
   19864: result <= 12'b011110001111;
   19865: result <= 12'b011110001111;
   19866: result <= 12'b011110001110;
   19867: result <= 12'b011110001110;
   19868: result <= 12'b011110001110;
   19869: result <= 12'b011110001110;
   19870: result <= 12'b011110001110;
   19871: result <= 12'b011110001110;
   19872: result <= 12'b011110001110;
   19873: result <= 12'b011110001110;
   19874: result <= 12'b011110001110;
   19875: result <= 12'b011110001110;
   19876: result <= 12'b011110001110;
   19877: result <= 12'b011110001110;
   19878: result <= 12'b011110001110;
   19879: result <= 12'b011110001110;
   19880: result <= 12'b011110001110;
   19881: result <= 12'b011110001101;
   19882: result <= 12'b011110001101;
   19883: result <= 12'b011110001101;
   19884: result <= 12'b011110001101;
   19885: result <= 12'b011110001101;
   19886: result <= 12'b011110001101;
   19887: result <= 12'b011110001101;
   19888: result <= 12'b011110001101;
   19889: result <= 12'b011110001101;
   19890: result <= 12'b011110001101;
   19891: result <= 12'b011110001101;
   19892: result <= 12'b011110001101;
   19893: result <= 12'b011110001101;
   19894: result <= 12'b011110001101;
   19895: result <= 12'b011110001101;
   19896: result <= 12'b011110001100;
   19897: result <= 12'b011110001100;
   19898: result <= 12'b011110001100;
   19899: result <= 12'b011110001100;
   19900: result <= 12'b011110001100;
   19901: result <= 12'b011110001100;
   19902: result <= 12'b011110001100;
   19903: result <= 12'b011110001100;
   19904: result <= 12'b011110001100;
   19905: result <= 12'b011110001100;
   19906: result <= 12'b011110001100;
   19907: result <= 12'b011110001100;
   19908: result <= 12'b011110001100;
   19909: result <= 12'b011110001100;
   19910: result <= 12'b011110001100;
   19911: result <= 12'b011110001100;
   19912: result <= 12'b011110001011;
   19913: result <= 12'b011110001011;
   19914: result <= 12'b011110001011;
   19915: result <= 12'b011110001011;
   19916: result <= 12'b011110001011;
   19917: result <= 12'b011110001011;
   19918: result <= 12'b011110001011;
   19919: result <= 12'b011110001011;
   19920: result <= 12'b011110001011;
   19921: result <= 12'b011110001011;
   19922: result <= 12'b011110001011;
   19923: result <= 12'b011110001011;
   19924: result <= 12'b011110001011;
   19925: result <= 12'b011110001011;
   19926: result <= 12'b011110001011;
   19927: result <= 12'b011110001010;
   19928: result <= 12'b011110001010;
   19929: result <= 12'b011110001010;
   19930: result <= 12'b011110001010;
   19931: result <= 12'b011110001010;
   19932: result <= 12'b011110001010;
   19933: result <= 12'b011110001010;
   19934: result <= 12'b011110001010;
   19935: result <= 12'b011110001010;
   19936: result <= 12'b011110001010;
   19937: result <= 12'b011110001010;
   19938: result <= 12'b011110001010;
   19939: result <= 12'b011110001010;
   19940: result <= 12'b011110001010;
   19941: result <= 12'b011110001010;
   19942: result <= 12'b011110001001;
   19943: result <= 12'b011110001001;
   19944: result <= 12'b011110001001;
   19945: result <= 12'b011110001001;
   19946: result <= 12'b011110001001;
   19947: result <= 12'b011110001001;
   19948: result <= 12'b011110001001;
   19949: result <= 12'b011110001001;
   19950: result <= 12'b011110001001;
   19951: result <= 12'b011110001001;
   19952: result <= 12'b011110001001;
   19953: result <= 12'b011110001001;
   19954: result <= 12'b011110001001;
   19955: result <= 12'b011110001001;
   19956: result <= 12'b011110001001;
   19957: result <= 12'b011110001001;
   19958: result <= 12'b011110001000;
   19959: result <= 12'b011110001000;
   19960: result <= 12'b011110001000;
   19961: result <= 12'b011110001000;
   19962: result <= 12'b011110001000;
   19963: result <= 12'b011110001000;
   19964: result <= 12'b011110001000;
   19965: result <= 12'b011110001000;
   19966: result <= 12'b011110001000;
   19967: result <= 12'b011110001000;
   19968: result <= 12'b011110001000;
   19969: result <= 12'b011110001000;
   19970: result <= 12'b011110001000;
   19971: result <= 12'b011110001000;
   19972: result <= 12'b011110001000;
   19973: result <= 12'b011110000111;
   19974: result <= 12'b011110000111;
   19975: result <= 12'b011110000111;
   19976: result <= 12'b011110000111;
   19977: result <= 12'b011110000111;
   19978: result <= 12'b011110000111;
   19979: result <= 12'b011110000111;
   19980: result <= 12'b011110000111;
   19981: result <= 12'b011110000111;
   19982: result <= 12'b011110000111;
   19983: result <= 12'b011110000111;
   19984: result <= 12'b011110000111;
   19985: result <= 12'b011110000111;
   19986: result <= 12'b011110000111;
   19987: result <= 12'b011110000111;
   19988: result <= 12'b011110000110;
   19989: result <= 12'b011110000110;
   19990: result <= 12'b011110000110;
   19991: result <= 12'b011110000110;
   19992: result <= 12'b011110000110;
   19993: result <= 12'b011110000110;
   19994: result <= 12'b011110000110;
   19995: result <= 12'b011110000110;
   19996: result <= 12'b011110000110;
   19997: result <= 12'b011110000110;
   19998: result <= 12'b011110000110;
   19999: result <= 12'b011110000110;
   20000: result <= 12'b011110000110;
   20001: result <= 12'b011110000110;
   20002: result <= 12'b011110000110;
   20003: result <= 12'b011110000101;
   20004: result <= 12'b011110000101;
   20005: result <= 12'b011110000101;
   20006: result <= 12'b011110000101;
   20007: result <= 12'b011110000101;
   20008: result <= 12'b011110000101;
   20009: result <= 12'b011110000101;
   20010: result <= 12'b011110000101;
   20011: result <= 12'b011110000101;
   20012: result <= 12'b011110000101;
   20013: result <= 12'b011110000101;
   20014: result <= 12'b011110000101;
   20015: result <= 12'b011110000101;
   20016: result <= 12'b011110000101;
   20017: result <= 12'b011110000101;
   20018: result <= 12'b011110000100;
   20019: result <= 12'b011110000100;
   20020: result <= 12'b011110000100;
   20021: result <= 12'b011110000100;
   20022: result <= 12'b011110000100;
   20023: result <= 12'b011110000100;
   20024: result <= 12'b011110000100;
   20025: result <= 12'b011110000100;
   20026: result <= 12'b011110000100;
   20027: result <= 12'b011110000100;
   20028: result <= 12'b011110000100;
   20029: result <= 12'b011110000100;
   20030: result <= 12'b011110000100;
   20031: result <= 12'b011110000100;
   20032: result <= 12'b011110000100;
   20033: result <= 12'b011110000011;
   20034: result <= 12'b011110000011;
   20035: result <= 12'b011110000011;
   20036: result <= 12'b011110000011;
   20037: result <= 12'b011110000011;
   20038: result <= 12'b011110000011;
   20039: result <= 12'b011110000011;
   20040: result <= 12'b011110000011;
   20041: result <= 12'b011110000011;
   20042: result <= 12'b011110000011;
   20043: result <= 12'b011110000011;
   20044: result <= 12'b011110000011;
   20045: result <= 12'b011110000011;
   20046: result <= 12'b011110000011;
   20047: result <= 12'b011110000011;
   20048: result <= 12'b011110000010;
   20049: result <= 12'b011110000010;
   20050: result <= 12'b011110000010;
   20051: result <= 12'b011110000010;
   20052: result <= 12'b011110000010;
   20053: result <= 12'b011110000010;
   20054: result <= 12'b011110000010;
   20055: result <= 12'b011110000010;
   20056: result <= 12'b011110000010;
   20057: result <= 12'b011110000010;
   20058: result <= 12'b011110000010;
   20059: result <= 12'b011110000010;
   20060: result <= 12'b011110000010;
   20061: result <= 12'b011110000010;
   20062: result <= 12'b011110000001;
   20063: result <= 12'b011110000001;
   20064: result <= 12'b011110000001;
   20065: result <= 12'b011110000001;
   20066: result <= 12'b011110000001;
   20067: result <= 12'b011110000001;
   20068: result <= 12'b011110000001;
   20069: result <= 12'b011110000001;
   20070: result <= 12'b011110000001;
   20071: result <= 12'b011110000001;
   20072: result <= 12'b011110000001;
   20073: result <= 12'b011110000001;
   20074: result <= 12'b011110000001;
   20075: result <= 12'b011110000001;
   20076: result <= 12'b011110000001;
   20077: result <= 12'b011110000000;
   20078: result <= 12'b011110000000;
   20079: result <= 12'b011110000000;
   20080: result <= 12'b011110000000;
   20081: result <= 12'b011110000000;
   20082: result <= 12'b011110000000;
   20083: result <= 12'b011110000000;
   20084: result <= 12'b011110000000;
   20085: result <= 12'b011110000000;
   20086: result <= 12'b011110000000;
   20087: result <= 12'b011110000000;
   20088: result <= 12'b011110000000;
   20089: result <= 12'b011110000000;
   20090: result <= 12'b011110000000;
   20091: result <= 12'b011110000000;
   20092: result <= 12'b011101111111;
   20093: result <= 12'b011101111111;
   20094: result <= 12'b011101111111;
   20095: result <= 12'b011101111111;
   20096: result <= 12'b011101111111;
   20097: result <= 12'b011101111111;
   20098: result <= 12'b011101111111;
   20099: result <= 12'b011101111111;
   20100: result <= 12'b011101111111;
   20101: result <= 12'b011101111111;
   20102: result <= 12'b011101111111;
   20103: result <= 12'b011101111111;
   20104: result <= 12'b011101111111;
   20105: result <= 12'b011101111111;
   20106: result <= 12'b011101111110;
   20107: result <= 12'b011101111110;
   20108: result <= 12'b011101111110;
   20109: result <= 12'b011101111110;
   20110: result <= 12'b011101111110;
   20111: result <= 12'b011101111110;
   20112: result <= 12'b011101111110;
   20113: result <= 12'b011101111110;
   20114: result <= 12'b011101111110;
   20115: result <= 12'b011101111110;
   20116: result <= 12'b011101111110;
   20117: result <= 12'b011101111110;
   20118: result <= 12'b011101111110;
   20119: result <= 12'b011101111110;
   20120: result <= 12'b011101111110;
   20121: result <= 12'b011101111101;
   20122: result <= 12'b011101111101;
   20123: result <= 12'b011101111101;
   20124: result <= 12'b011101111101;
   20125: result <= 12'b011101111101;
   20126: result <= 12'b011101111101;
   20127: result <= 12'b011101111101;
   20128: result <= 12'b011101111101;
   20129: result <= 12'b011101111101;
   20130: result <= 12'b011101111101;
   20131: result <= 12'b011101111101;
   20132: result <= 12'b011101111101;
   20133: result <= 12'b011101111101;
   20134: result <= 12'b011101111101;
   20135: result <= 12'b011101111100;
   20136: result <= 12'b011101111100;
   20137: result <= 12'b011101111100;
   20138: result <= 12'b011101111100;
   20139: result <= 12'b011101111100;
   20140: result <= 12'b011101111100;
   20141: result <= 12'b011101111100;
   20142: result <= 12'b011101111100;
   20143: result <= 12'b011101111100;
   20144: result <= 12'b011101111100;
   20145: result <= 12'b011101111100;
   20146: result <= 12'b011101111100;
   20147: result <= 12'b011101111100;
   20148: result <= 12'b011101111100;
   20149: result <= 12'b011101111100;
   20150: result <= 12'b011101111011;
   20151: result <= 12'b011101111011;
   20152: result <= 12'b011101111011;
   20153: result <= 12'b011101111011;
   20154: result <= 12'b011101111011;
   20155: result <= 12'b011101111011;
   20156: result <= 12'b011101111011;
   20157: result <= 12'b011101111011;
   20158: result <= 12'b011101111011;
   20159: result <= 12'b011101111011;
   20160: result <= 12'b011101111011;
   20161: result <= 12'b011101111011;
   20162: result <= 12'b011101111011;
   20163: result <= 12'b011101111011;
   20164: result <= 12'b011101111010;
   20165: result <= 12'b011101111010;
   20166: result <= 12'b011101111010;
   20167: result <= 12'b011101111010;
   20168: result <= 12'b011101111010;
   20169: result <= 12'b011101111010;
   20170: result <= 12'b011101111010;
   20171: result <= 12'b011101111010;
   20172: result <= 12'b011101111010;
   20173: result <= 12'b011101111010;
   20174: result <= 12'b011101111010;
   20175: result <= 12'b011101111010;
   20176: result <= 12'b011101111010;
   20177: result <= 12'b011101111010;
   20178: result <= 12'b011101111010;
   20179: result <= 12'b011101111001;
   20180: result <= 12'b011101111001;
   20181: result <= 12'b011101111001;
   20182: result <= 12'b011101111001;
   20183: result <= 12'b011101111001;
   20184: result <= 12'b011101111001;
   20185: result <= 12'b011101111001;
   20186: result <= 12'b011101111001;
   20187: result <= 12'b011101111001;
   20188: result <= 12'b011101111001;
   20189: result <= 12'b011101111001;
   20190: result <= 12'b011101111001;
   20191: result <= 12'b011101111001;
   20192: result <= 12'b011101111001;
   20193: result <= 12'b011101111000;
   20194: result <= 12'b011101111000;
   20195: result <= 12'b011101111000;
   20196: result <= 12'b011101111000;
   20197: result <= 12'b011101111000;
   20198: result <= 12'b011101111000;
   20199: result <= 12'b011101111000;
   20200: result <= 12'b011101111000;
   20201: result <= 12'b011101111000;
   20202: result <= 12'b011101111000;
   20203: result <= 12'b011101111000;
   20204: result <= 12'b011101111000;
   20205: result <= 12'b011101111000;
   20206: result <= 12'b011101111000;
   20207: result <= 12'b011101110111;
   20208: result <= 12'b011101110111;
   20209: result <= 12'b011101110111;
   20210: result <= 12'b011101110111;
   20211: result <= 12'b011101110111;
   20212: result <= 12'b011101110111;
   20213: result <= 12'b011101110111;
   20214: result <= 12'b011101110111;
   20215: result <= 12'b011101110111;
   20216: result <= 12'b011101110111;
   20217: result <= 12'b011101110111;
   20218: result <= 12'b011101110111;
   20219: result <= 12'b011101110111;
   20220: result <= 12'b011101110111;
   20221: result <= 12'b011101110110;
   20222: result <= 12'b011101110110;
   20223: result <= 12'b011101110110;
   20224: result <= 12'b011101110110;
   20225: result <= 12'b011101110110;
   20226: result <= 12'b011101110110;
   20227: result <= 12'b011101110110;
   20228: result <= 12'b011101110110;
   20229: result <= 12'b011101110110;
   20230: result <= 12'b011101110110;
   20231: result <= 12'b011101110110;
   20232: result <= 12'b011101110110;
   20233: result <= 12'b011101110110;
   20234: result <= 12'b011101110110;
   20235: result <= 12'b011101110101;
   20236: result <= 12'b011101110101;
   20237: result <= 12'b011101110101;
   20238: result <= 12'b011101110101;
   20239: result <= 12'b011101110101;
   20240: result <= 12'b011101110101;
   20241: result <= 12'b011101110101;
   20242: result <= 12'b011101110101;
   20243: result <= 12'b011101110101;
   20244: result <= 12'b011101110101;
   20245: result <= 12'b011101110101;
   20246: result <= 12'b011101110101;
   20247: result <= 12'b011101110101;
   20248: result <= 12'b011101110101;
   20249: result <= 12'b011101110100;
   20250: result <= 12'b011101110100;
   20251: result <= 12'b011101110100;
   20252: result <= 12'b011101110100;
   20253: result <= 12'b011101110100;
   20254: result <= 12'b011101110100;
   20255: result <= 12'b011101110100;
   20256: result <= 12'b011101110100;
   20257: result <= 12'b011101110100;
   20258: result <= 12'b011101110100;
   20259: result <= 12'b011101110100;
   20260: result <= 12'b011101110100;
   20261: result <= 12'b011101110100;
   20262: result <= 12'b011101110100;
   20263: result <= 12'b011101110011;
   20264: result <= 12'b011101110011;
   20265: result <= 12'b011101110011;
   20266: result <= 12'b011101110011;
   20267: result <= 12'b011101110011;
   20268: result <= 12'b011101110011;
   20269: result <= 12'b011101110011;
   20270: result <= 12'b011101110011;
   20271: result <= 12'b011101110011;
   20272: result <= 12'b011101110011;
   20273: result <= 12'b011101110011;
   20274: result <= 12'b011101110011;
   20275: result <= 12'b011101110011;
   20276: result <= 12'b011101110011;
   20277: result <= 12'b011101110010;
   20278: result <= 12'b011101110010;
   20279: result <= 12'b011101110010;
   20280: result <= 12'b011101110010;
   20281: result <= 12'b011101110010;
   20282: result <= 12'b011101110010;
   20283: result <= 12'b011101110010;
   20284: result <= 12'b011101110010;
   20285: result <= 12'b011101110010;
   20286: result <= 12'b011101110010;
   20287: result <= 12'b011101110010;
   20288: result <= 12'b011101110010;
   20289: result <= 12'b011101110010;
   20290: result <= 12'b011101110010;
   20291: result <= 12'b011101110001;
   20292: result <= 12'b011101110001;
   20293: result <= 12'b011101110001;
   20294: result <= 12'b011101110001;
   20295: result <= 12'b011101110001;
   20296: result <= 12'b011101110001;
   20297: result <= 12'b011101110001;
   20298: result <= 12'b011101110001;
   20299: result <= 12'b011101110001;
   20300: result <= 12'b011101110001;
   20301: result <= 12'b011101110001;
   20302: result <= 12'b011101110001;
   20303: result <= 12'b011101110001;
   20304: result <= 12'b011101110001;
   20305: result <= 12'b011101110000;
   20306: result <= 12'b011101110000;
   20307: result <= 12'b011101110000;
   20308: result <= 12'b011101110000;
   20309: result <= 12'b011101110000;
   20310: result <= 12'b011101110000;
   20311: result <= 12'b011101110000;
   20312: result <= 12'b011101110000;
   20313: result <= 12'b011101110000;
   20314: result <= 12'b011101110000;
   20315: result <= 12'b011101110000;
   20316: result <= 12'b011101110000;
   20317: result <= 12'b011101110000;
   20318: result <= 12'b011101110000;
   20319: result <= 12'b011101101111;
   20320: result <= 12'b011101101111;
   20321: result <= 12'b011101101111;
   20322: result <= 12'b011101101111;
   20323: result <= 12'b011101101111;
   20324: result <= 12'b011101101111;
   20325: result <= 12'b011101101111;
   20326: result <= 12'b011101101111;
   20327: result <= 12'b011101101111;
   20328: result <= 12'b011101101111;
   20329: result <= 12'b011101101111;
   20330: result <= 12'b011101101111;
   20331: result <= 12'b011101101111;
   20332: result <= 12'b011101101111;
   20333: result <= 12'b011101101110;
   20334: result <= 12'b011101101110;
   20335: result <= 12'b011101101110;
   20336: result <= 12'b011101101110;
   20337: result <= 12'b011101101110;
   20338: result <= 12'b011101101110;
   20339: result <= 12'b011101101110;
   20340: result <= 12'b011101101110;
   20341: result <= 12'b011101101110;
   20342: result <= 12'b011101101110;
   20343: result <= 12'b011101101110;
   20344: result <= 12'b011101101110;
   20345: result <= 12'b011101101110;
   20346: result <= 12'b011101101110;
   20347: result <= 12'b011101101101;
   20348: result <= 12'b011101101101;
   20349: result <= 12'b011101101101;
   20350: result <= 12'b011101101101;
   20351: result <= 12'b011101101101;
   20352: result <= 12'b011101101101;
   20353: result <= 12'b011101101101;
   20354: result <= 12'b011101101101;
   20355: result <= 12'b011101101101;
   20356: result <= 12'b011101101101;
   20357: result <= 12'b011101101101;
   20358: result <= 12'b011101101101;
   20359: result <= 12'b011101101101;
   20360: result <= 12'b011101101100;
   20361: result <= 12'b011101101100;
   20362: result <= 12'b011101101100;
   20363: result <= 12'b011101101100;
   20364: result <= 12'b011101101100;
   20365: result <= 12'b011101101100;
   20366: result <= 12'b011101101100;
   20367: result <= 12'b011101101100;
   20368: result <= 12'b011101101100;
   20369: result <= 12'b011101101100;
   20370: result <= 12'b011101101100;
   20371: result <= 12'b011101101100;
   20372: result <= 12'b011101101100;
   20373: result <= 12'b011101101100;
   20374: result <= 12'b011101101011;
   20375: result <= 12'b011101101011;
   20376: result <= 12'b011101101011;
   20377: result <= 12'b011101101011;
   20378: result <= 12'b011101101011;
   20379: result <= 12'b011101101011;
   20380: result <= 12'b011101101011;
   20381: result <= 12'b011101101011;
   20382: result <= 12'b011101101011;
   20383: result <= 12'b011101101011;
   20384: result <= 12'b011101101011;
   20385: result <= 12'b011101101011;
   20386: result <= 12'b011101101011;
   20387: result <= 12'b011101101011;
   20388: result <= 12'b011101101010;
   20389: result <= 12'b011101101010;
   20390: result <= 12'b011101101010;
   20391: result <= 12'b011101101010;
   20392: result <= 12'b011101101010;
   20393: result <= 12'b011101101010;
   20394: result <= 12'b011101101010;
   20395: result <= 12'b011101101010;
   20396: result <= 12'b011101101010;
   20397: result <= 12'b011101101010;
   20398: result <= 12'b011101101010;
   20399: result <= 12'b011101101010;
   20400: result <= 12'b011101101010;
   20401: result <= 12'b011101101001;
   20402: result <= 12'b011101101001;
   20403: result <= 12'b011101101001;
   20404: result <= 12'b011101101001;
   20405: result <= 12'b011101101001;
   20406: result <= 12'b011101101001;
   20407: result <= 12'b011101101001;
   20408: result <= 12'b011101101001;
   20409: result <= 12'b011101101001;
   20410: result <= 12'b011101101001;
   20411: result <= 12'b011101101001;
   20412: result <= 12'b011101101001;
   20413: result <= 12'b011101101001;
   20414: result <= 12'b011101101001;
   20415: result <= 12'b011101101000;
   20416: result <= 12'b011101101000;
   20417: result <= 12'b011101101000;
   20418: result <= 12'b011101101000;
   20419: result <= 12'b011101101000;
   20420: result <= 12'b011101101000;
   20421: result <= 12'b011101101000;
   20422: result <= 12'b011101101000;
   20423: result <= 12'b011101101000;
   20424: result <= 12'b011101101000;
   20425: result <= 12'b011101101000;
   20426: result <= 12'b011101101000;
   20427: result <= 12'b011101101000;
   20428: result <= 12'b011101100111;
   20429: result <= 12'b011101100111;
   20430: result <= 12'b011101100111;
   20431: result <= 12'b011101100111;
   20432: result <= 12'b011101100111;
   20433: result <= 12'b011101100111;
   20434: result <= 12'b011101100111;
   20435: result <= 12'b011101100111;
   20436: result <= 12'b011101100111;
   20437: result <= 12'b011101100111;
   20438: result <= 12'b011101100111;
   20439: result <= 12'b011101100111;
   20440: result <= 12'b011101100111;
   20441: result <= 12'b011101100111;
   20442: result <= 12'b011101100110;
   20443: result <= 12'b011101100110;
   20444: result <= 12'b011101100110;
   20445: result <= 12'b011101100110;
   20446: result <= 12'b011101100110;
   20447: result <= 12'b011101100110;
   20448: result <= 12'b011101100110;
   20449: result <= 12'b011101100110;
   20450: result <= 12'b011101100110;
   20451: result <= 12'b011101100110;
   20452: result <= 12'b011101100110;
   20453: result <= 12'b011101100110;
   20454: result <= 12'b011101100110;
   20455: result <= 12'b011101100101;
   20456: result <= 12'b011101100101;
   20457: result <= 12'b011101100101;
   20458: result <= 12'b011101100101;
   20459: result <= 12'b011101100101;
   20460: result <= 12'b011101100101;
   20461: result <= 12'b011101100101;
   20462: result <= 12'b011101100101;
   20463: result <= 12'b011101100101;
   20464: result <= 12'b011101100101;
   20465: result <= 12'b011101100101;
   20466: result <= 12'b011101100101;
   20467: result <= 12'b011101100101;
   20468: result <= 12'b011101100101;
   20469: result <= 12'b011101100100;
   20470: result <= 12'b011101100100;
   20471: result <= 12'b011101100100;
   20472: result <= 12'b011101100100;
   20473: result <= 12'b011101100100;
   20474: result <= 12'b011101100100;
   20475: result <= 12'b011101100100;
   20476: result <= 12'b011101100100;
   20477: result <= 12'b011101100100;
   20478: result <= 12'b011101100100;
   20479: result <= 12'b011101100100;
   20480: result <= 12'b011101100100;
   20481: result <= 12'b011101100100;
   20482: result <= 12'b011101100011;
   20483: result <= 12'b011101100011;
   20484: result <= 12'b011101100011;
   20485: result <= 12'b011101100011;
   20486: result <= 12'b011101100011;
   20487: result <= 12'b011101100011;
   20488: result <= 12'b011101100011;
   20489: result <= 12'b011101100011;
   20490: result <= 12'b011101100011;
   20491: result <= 12'b011101100011;
   20492: result <= 12'b011101100011;
   20493: result <= 12'b011101100011;
   20494: result <= 12'b011101100011;
   20495: result <= 12'b011101100010;
   20496: result <= 12'b011101100010;
   20497: result <= 12'b011101100010;
   20498: result <= 12'b011101100010;
   20499: result <= 12'b011101100010;
   20500: result <= 12'b011101100010;
   20501: result <= 12'b011101100010;
   20502: result <= 12'b011101100010;
   20503: result <= 12'b011101100010;
   20504: result <= 12'b011101100010;
   20505: result <= 12'b011101100010;
   20506: result <= 12'b011101100010;
   20507: result <= 12'b011101100010;
   20508: result <= 12'b011101100001;
   20509: result <= 12'b011101100001;
   20510: result <= 12'b011101100001;
   20511: result <= 12'b011101100001;
   20512: result <= 12'b011101100001;
   20513: result <= 12'b011101100001;
   20514: result <= 12'b011101100001;
   20515: result <= 12'b011101100001;
   20516: result <= 12'b011101100001;
   20517: result <= 12'b011101100001;
   20518: result <= 12'b011101100001;
   20519: result <= 12'b011101100001;
   20520: result <= 12'b011101100001;
   20521: result <= 12'b011101100001;
   20522: result <= 12'b011101100000;
   20523: result <= 12'b011101100000;
   20524: result <= 12'b011101100000;
   20525: result <= 12'b011101100000;
   20526: result <= 12'b011101100000;
   20527: result <= 12'b011101100000;
   20528: result <= 12'b011101100000;
   20529: result <= 12'b011101100000;
   20530: result <= 12'b011101100000;
   20531: result <= 12'b011101100000;
   20532: result <= 12'b011101100000;
   20533: result <= 12'b011101100000;
   20534: result <= 12'b011101100000;
   20535: result <= 12'b011101011111;
   20536: result <= 12'b011101011111;
   20537: result <= 12'b011101011111;
   20538: result <= 12'b011101011111;
   20539: result <= 12'b011101011111;
   20540: result <= 12'b011101011111;
   20541: result <= 12'b011101011111;
   20542: result <= 12'b011101011111;
   20543: result <= 12'b011101011111;
   20544: result <= 12'b011101011111;
   20545: result <= 12'b011101011111;
   20546: result <= 12'b011101011111;
   20547: result <= 12'b011101011111;
   20548: result <= 12'b011101011110;
   20549: result <= 12'b011101011110;
   20550: result <= 12'b011101011110;
   20551: result <= 12'b011101011110;
   20552: result <= 12'b011101011110;
   20553: result <= 12'b011101011110;
   20554: result <= 12'b011101011110;
   20555: result <= 12'b011101011110;
   20556: result <= 12'b011101011110;
   20557: result <= 12'b011101011110;
   20558: result <= 12'b011101011110;
   20559: result <= 12'b011101011110;
   20560: result <= 12'b011101011110;
   20561: result <= 12'b011101011101;
   20562: result <= 12'b011101011101;
   20563: result <= 12'b011101011101;
   20564: result <= 12'b011101011101;
   20565: result <= 12'b011101011101;
   20566: result <= 12'b011101011101;
   20567: result <= 12'b011101011101;
   20568: result <= 12'b011101011101;
   20569: result <= 12'b011101011101;
   20570: result <= 12'b011101011101;
   20571: result <= 12'b011101011101;
   20572: result <= 12'b011101011101;
   20573: result <= 12'b011101011101;
   20574: result <= 12'b011101011100;
   20575: result <= 12'b011101011100;
   20576: result <= 12'b011101011100;
   20577: result <= 12'b011101011100;
   20578: result <= 12'b011101011100;
   20579: result <= 12'b011101011100;
   20580: result <= 12'b011101011100;
   20581: result <= 12'b011101011100;
   20582: result <= 12'b011101011100;
   20583: result <= 12'b011101011100;
   20584: result <= 12'b011101011100;
   20585: result <= 12'b011101011100;
   20586: result <= 12'b011101011100;
   20587: result <= 12'b011101011011;
   20588: result <= 12'b011101011011;
   20589: result <= 12'b011101011011;
   20590: result <= 12'b011101011011;
   20591: result <= 12'b011101011011;
   20592: result <= 12'b011101011011;
   20593: result <= 12'b011101011011;
   20594: result <= 12'b011101011011;
   20595: result <= 12'b011101011011;
   20596: result <= 12'b011101011011;
   20597: result <= 12'b011101011011;
   20598: result <= 12'b011101011011;
   20599: result <= 12'b011101011011;
   20600: result <= 12'b011101011010;
   20601: result <= 12'b011101011010;
   20602: result <= 12'b011101011010;
   20603: result <= 12'b011101011010;
   20604: result <= 12'b011101011010;
   20605: result <= 12'b011101011010;
   20606: result <= 12'b011101011010;
   20607: result <= 12'b011101011010;
   20608: result <= 12'b011101011010;
   20609: result <= 12'b011101011010;
   20610: result <= 12'b011101011010;
   20611: result <= 12'b011101011010;
   20612: result <= 12'b011101011010;
   20613: result <= 12'b011101011001;
   20614: result <= 12'b011101011001;
   20615: result <= 12'b011101011001;
   20616: result <= 12'b011101011001;
   20617: result <= 12'b011101011001;
   20618: result <= 12'b011101011001;
   20619: result <= 12'b011101011001;
   20620: result <= 12'b011101011001;
   20621: result <= 12'b011101011001;
   20622: result <= 12'b011101011001;
   20623: result <= 12'b011101011001;
   20624: result <= 12'b011101011001;
   20625: result <= 12'b011101011001;
   20626: result <= 12'b011101011000;
   20627: result <= 12'b011101011000;
   20628: result <= 12'b011101011000;
   20629: result <= 12'b011101011000;
   20630: result <= 12'b011101011000;
   20631: result <= 12'b011101011000;
   20632: result <= 12'b011101011000;
   20633: result <= 12'b011101011000;
   20634: result <= 12'b011101011000;
   20635: result <= 12'b011101011000;
   20636: result <= 12'b011101011000;
   20637: result <= 12'b011101011000;
   20638: result <= 12'b011101011000;
   20639: result <= 12'b011101010111;
   20640: result <= 12'b011101010111;
   20641: result <= 12'b011101010111;
   20642: result <= 12'b011101010111;
   20643: result <= 12'b011101010111;
   20644: result <= 12'b011101010111;
   20645: result <= 12'b011101010111;
   20646: result <= 12'b011101010111;
   20647: result <= 12'b011101010111;
   20648: result <= 12'b011101010111;
   20649: result <= 12'b011101010111;
   20650: result <= 12'b011101010111;
   20651: result <= 12'b011101010111;
   20652: result <= 12'b011101010110;
   20653: result <= 12'b011101010110;
   20654: result <= 12'b011101010110;
   20655: result <= 12'b011101010110;
   20656: result <= 12'b011101010110;
   20657: result <= 12'b011101010110;
   20658: result <= 12'b011101010110;
   20659: result <= 12'b011101010110;
   20660: result <= 12'b011101010110;
   20661: result <= 12'b011101010110;
   20662: result <= 12'b011101010110;
   20663: result <= 12'b011101010110;
   20664: result <= 12'b011101010101;
   20665: result <= 12'b011101010101;
   20666: result <= 12'b011101010101;
   20667: result <= 12'b011101010101;
   20668: result <= 12'b011101010101;
   20669: result <= 12'b011101010101;
   20670: result <= 12'b011101010101;
   20671: result <= 12'b011101010101;
   20672: result <= 12'b011101010101;
   20673: result <= 12'b011101010101;
   20674: result <= 12'b011101010101;
   20675: result <= 12'b011101010101;
   20676: result <= 12'b011101010101;
   20677: result <= 12'b011101010100;
   20678: result <= 12'b011101010100;
   20679: result <= 12'b011101010100;
   20680: result <= 12'b011101010100;
   20681: result <= 12'b011101010100;
   20682: result <= 12'b011101010100;
   20683: result <= 12'b011101010100;
   20684: result <= 12'b011101010100;
   20685: result <= 12'b011101010100;
   20686: result <= 12'b011101010100;
   20687: result <= 12'b011101010100;
   20688: result <= 12'b011101010100;
   20689: result <= 12'b011101010100;
   20690: result <= 12'b011101010011;
   20691: result <= 12'b011101010011;
   20692: result <= 12'b011101010011;
   20693: result <= 12'b011101010011;
   20694: result <= 12'b011101010011;
   20695: result <= 12'b011101010011;
   20696: result <= 12'b011101010011;
   20697: result <= 12'b011101010011;
   20698: result <= 12'b011101010011;
   20699: result <= 12'b011101010011;
   20700: result <= 12'b011101010011;
   20701: result <= 12'b011101010011;
   20702: result <= 12'b011101010010;
   20703: result <= 12'b011101010010;
   20704: result <= 12'b011101010010;
   20705: result <= 12'b011101010010;
   20706: result <= 12'b011101010010;
   20707: result <= 12'b011101010010;
   20708: result <= 12'b011101010010;
   20709: result <= 12'b011101010010;
   20710: result <= 12'b011101010010;
   20711: result <= 12'b011101010010;
   20712: result <= 12'b011101010010;
   20713: result <= 12'b011101010010;
   20714: result <= 12'b011101010010;
   20715: result <= 12'b011101010001;
   20716: result <= 12'b011101010001;
   20717: result <= 12'b011101010001;
   20718: result <= 12'b011101010001;
   20719: result <= 12'b011101010001;
   20720: result <= 12'b011101010001;
   20721: result <= 12'b011101010001;
   20722: result <= 12'b011101010001;
   20723: result <= 12'b011101010001;
   20724: result <= 12'b011101010001;
   20725: result <= 12'b011101010001;
   20726: result <= 12'b011101010001;
   20727: result <= 12'b011101010001;
   20728: result <= 12'b011101010000;
   20729: result <= 12'b011101010000;
   20730: result <= 12'b011101010000;
   20731: result <= 12'b011101010000;
   20732: result <= 12'b011101010000;
   20733: result <= 12'b011101010000;
   20734: result <= 12'b011101010000;
   20735: result <= 12'b011101010000;
   20736: result <= 12'b011101010000;
   20737: result <= 12'b011101010000;
   20738: result <= 12'b011101010000;
   20739: result <= 12'b011101010000;
   20740: result <= 12'b011101001111;
   20741: result <= 12'b011101001111;
   20742: result <= 12'b011101001111;
   20743: result <= 12'b011101001111;
   20744: result <= 12'b011101001111;
   20745: result <= 12'b011101001111;
   20746: result <= 12'b011101001111;
   20747: result <= 12'b011101001111;
   20748: result <= 12'b011101001111;
   20749: result <= 12'b011101001111;
   20750: result <= 12'b011101001111;
   20751: result <= 12'b011101001111;
   20752: result <= 12'b011101001111;
   20753: result <= 12'b011101001110;
   20754: result <= 12'b011101001110;
   20755: result <= 12'b011101001110;
   20756: result <= 12'b011101001110;
   20757: result <= 12'b011101001110;
   20758: result <= 12'b011101001110;
   20759: result <= 12'b011101001110;
   20760: result <= 12'b011101001110;
   20761: result <= 12'b011101001110;
   20762: result <= 12'b011101001110;
   20763: result <= 12'b011101001110;
   20764: result <= 12'b011101001110;
   20765: result <= 12'b011101001101;
   20766: result <= 12'b011101001101;
   20767: result <= 12'b011101001101;
   20768: result <= 12'b011101001101;
   20769: result <= 12'b011101001101;
   20770: result <= 12'b011101001101;
   20771: result <= 12'b011101001101;
   20772: result <= 12'b011101001101;
   20773: result <= 12'b011101001101;
   20774: result <= 12'b011101001101;
   20775: result <= 12'b011101001101;
   20776: result <= 12'b011101001101;
   20777: result <= 12'b011101001101;
   20778: result <= 12'b011101001100;
   20779: result <= 12'b011101001100;
   20780: result <= 12'b011101001100;
   20781: result <= 12'b011101001100;
   20782: result <= 12'b011101001100;
   20783: result <= 12'b011101001100;
   20784: result <= 12'b011101001100;
   20785: result <= 12'b011101001100;
   20786: result <= 12'b011101001100;
   20787: result <= 12'b011101001100;
   20788: result <= 12'b011101001100;
   20789: result <= 12'b011101001100;
   20790: result <= 12'b011101001011;
   20791: result <= 12'b011101001011;
   20792: result <= 12'b011101001011;
   20793: result <= 12'b011101001011;
   20794: result <= 12'b011101001011;
   20795: result <= 12'b011101001011;
   20796: result <= 12'b011101001011;
   20797: result <= 12'b011101001011;
   20798: result <= 12'b011101001011;
   20799: result <= 12'b011101001011;
   20800: result <= 12'b011101001011;
   20801: result <= 12'b011101001011;
   20802: result <= 12'b011101001011;
   20803: result <= 12'b011101001010;
   20804: result <= 12'b011101001010;
   20805: result <= 12'b011101001010;
   20806: result <= 12'b011101001010;
   20807: result <= 12'b011101001010;
   20808: result <= 12'b011101001010;
   20809: result <= 12'b011101001010;
   20810: result <= 12'b011101001010;
   20811: result <= 12'b011101001010;
   20812: result <= 12'b011101001010;
   20813: result <= 12'b011101001010;
   20814: result <= 12'b011101001010;
   20815: result <= 12'b011101001001;
   20816: result <= 12'b011101001001;
   20817: result <= 12'b011101001001;
   20818: result <= 12'b011101001001;
   20819: result <= 12'b011101001001;
   20820: result <= 12'b011101001001;
   20821: result <= 12'b011101001001;
   20822: result <= 12'b011101001001;
   20823: result <= 12'b011101001001;
   20824: result <= 12'b011101001001;
   20825: result <= 12'b011101001001;
   20826: result <= 12'b011101001001;
   20827: result <= 12'b011101001000;
   20828: result <= 12'b011101001000;
   20829: result <= 12'b011101001000;
   20830: result <= 12'b011101001000;
   20831: result <= 12'b011101001000;
   20832: result <= 12'b011101001000;
   20833: result <= 12'b011101001000;
   20834: result <= 12'b011101001000;
   20835: result <= 12'b011101001000;
   20836: result <= 12'b011101001000;
   20837: result <= 12'b011101001000;
   20838: result <= 12'b011101001000;
   20839: result <= 12'b011101001000;
   20840: result <= 12'b011101000111;
   20841: result <= 12'b011101000111;
   20842: result <= 12'b011101000111;
   20843: result <= 12'b011101000111;
   20844: result <= 12'b011101000111;
   20845: result <= 12'b011101000111;
   20846: result <= 12'b011101000111;
   20847: result <= 12'b011101000111;
   20848: result <= 12'b011101000111;
   20849: result <= 12'b011101000111;
   20850: result <= 12'b011101000111;
   20851: result <= 12'b011101000111;
   20852: result <= 12'b011101000110;
   20853: result <= 12'b011101000110;
   20854: result <= 12'b011101000110;
   20855: result <= 12'b011101000110;
   20856: result <= 12'b011101000110;
   20857: result <= 12'b011101000110;
   20858: result <= 12'b011101000110;
   20859: result <= 12'b011101000110;
   20860: result <= 12'b011101000110;
   20861: result <= 12'b011101000110;
   20862: result <= 12'b011101000110;
   20863: result <= 12'b011101000110;
   20864: result <= 12'b011101000101;
   20865: result <= 12'b011101000101;
   20866: result <= 12'b011101000101;
   20867: result <= 12'b011101000101;
   20868: result <= 12'b011101000101;
   20869: result <= 12'b011101000101;
   20870: result <= 12'b011101000101;
   20871: result <= 12'b011101000101;
   20872: result <= 12'b011101000101;
   20873: result <= 12'b011101000101;
   20874: result <= 12'b011101000101;
   20875: result <= 12'b011101000101;
   20876: result <= 12'b011101000100;
   20877: result <= 12'b011101000100;
   20878: result <= 12'b011101000100;
   20879: result <= 12'b011101000100;
   20880: result <= 12'b011101000100;
   20881: result <= 12'b011101000100;
   20882: result <= 12'b011101000100;
   20883: result <= 12'b011101000100;
   20884: result <= 12'b011101000100;
   20885: result <= 12'b011101000100;
   20886: result <= 12'b011101000100;
   20887: result <= 12'b011101000100;
   20888: result <= 12'b011101000100;
   20889: result <= 12'b011101000011;
   20890: result <= 12'b011101000011;
   20891: result <= 12'b011101000011;
   20892: result <= 12'b011101000011;
   20893: result <= 12'b011101000011;
   20894: result <= 12'b011101000011;
   20895: result <= 12'b011101000011;
   20896: result <= 12'b011101000011;
   20897: result <= 12'b011101000011;
   20898: result <= 12'b011101000011;
   20899: result <= 12'b011101000011;
   20900: result <= 12'b011101000011;
   20901: result <= 12'b011101000010;
   20902: result <= 12'b011101000010;
   20903: result <= 12'b011101000010;
   20904: result <= 12'b011101000010;
   20905: result <= 12'b011101000010;
   20906: result <= 12'b011101000010;
   20907: result <= 12'b011101000010;
   20908: result <= 12'b011101000010;
   20909: result <= 12'b011101000010;
   20910: result <= 12'b011101000010;
   20911: result <= 12'b011101000010;
   20912: result <= 12'b011101000010;
   20913: result <= 12'b011101000001;
   20914: result <= 12'b011101000001;
   20915: result <= 12'b011101000001;
   20916: result <= 12'b011101000001;
   20917: result <= 12'b011101000001;
   20918: result <= 12'b011101000001;
   20919: result <= 12'b011101000001;
   20920: result <= 12'b011101000001;
   20921: result <= 12'b011101000001;
   20922: result <= 12'b011101000001;
   20923: result <= 12'b011101000001;
   20924: result <= 12'b011101000001;
   20925: result <= 12'b011101000000;
   20926: result <= 12'b011101000000;
   20927: result <= 12'b011101000000;
   20928: result <= 12'b011101000000;
   20929: result <= 12'b011101000000;
   20930: result <= 12'b011101000000;
   20931: result <= 12'b011101000000;
   20932: result <= 12'b011101000000;
   20933: result <= 12'b011101000000;
   20934: result <= 12'b011101000000;
   20935: result <= 12'b011101000000;
   20936: result <= 12'b011101000000;
   20937: result <= 12'b011100111111;
   20938: result <= 12'b011100111111;
   20939: result <= 12'b011100111111;
   20940: result <= 12'b011100111111;
   20941: result <= 12'b011100111111;
   20942: result <= 12'b011100111111;
   20943: result <= 12'b011100111111;
   20944: result <= 12'b011100111111;
   20945: result <= 12'b011100111111;
   20946: result <= 12'b011100111111;
   20947: result <= 12'b011100111111;
   20948: result <= 12'b011100111111;
   20949: result <= 12'b011100111110;
   20950: result <= 12'b011100111110;
   20951: result <= 12'b011100111110;
   20952: result <= 12'b011100111110;
   20953: result <= 12'b011100111110;
   20954: result <= 12'b011100111110;
   20955: result <= 12'b011100111110;
   20956: result <= 12'b011100111110;
   20957: result <= 12'b011100111110;
   20958: result <= 12'b011100111110;
   20959: result <= 12'b011100111110;
   20960: result <= 12'b011100111110;
   20961: result <= 12'b011100111101;
   20962: result <= 12'b011100111101;
   20963: result <= 12'b011100111101;
   20964: result <= 12'b011100111101;
   20965: result <= 12'b011100111101;
   20966: result <= 12'b011100111101;
   20967: result <= 12'b011100111101;
   20968: result <= 12'b011100111101;
   20969: result <= 12'b011100111101;
   20970: result <= 12'b011100111101;
   20971: result <= 12'b011100111101;
   20972: result <= 12'b011100111101;
   20973: result <= 12'b011100111100;
   20974: result <= 12'b011100111100;
   20975: result <= 12'b011100111100;
   20976: result <= 12'b011100111100;
   20977: result <= 12'b011100111100;
   20978: result <= 12'b011100111100;
   20979: result <= 12'b011100111100;
   20980: result <= 12'b011100111100;
   20981: result <= 12'b011100111100;
   20982: result <= 12'b011100111100;
   20983: result <= 12'b011100111100;
   20984: result <= 12'b011100111100;
   20985: result <= 12'b011100111011;
   20986: result <= 12'b011100111011;
   20987: result <= 12'b011100111011;
   20988: result <= 12'b011100111011;
   20989: result <= 12'b011100111011;
   20990: result <= 12'b011100111011;
   20991: result <= 12'b011100111011;
   20992: result <= 12'b011100111011;
   20993: result <= 12'b011100111011;
   20994: result <= 12'b011100111011;
   20995: result <= 12'b011100111011;
   20996: result <= 12'b011100111011;
   20997: result <= 12'b011100111010;
   20998: result <= 12'b011100111010;
   20999: result <= 12'b011100111010;
   21000: result <= 12'b011100111010;
   21001: result <= 12'b011100111010;
   21002: result <= 12'b011100111010;
   21003: result <= 12'b011100111010;
   21004: result <= 12'b011100111010;
   21005: result <= 12'b011100111010;
   21006: result <= 12'b011100111010;
   21007: result <= 12'b011100111010;
   21008: result <= 12'b011100111010;
   21009: result <= 12'b011100111001;
   21010: result <= 12'b011100111001;
   21011: result <= 12'b011100111001;
   21012: result <= 12'b011100111001;
   21013: result <= 12'b011100111001;
   21014: result <= 12'b011100111001;
   21015: result <= 12'b011100111001;
   21016: result <= 12'b011100111001;
   21017: result <= 12'b011100111001;
   21018: result <= 12'b011100111001;
   21019: result <= 12'b011100111001;
   21020: result <= 12'b011100111001;
   21021: result <= 12'b011100111000;
   21022: result <= 12'b011100111000;
   21023: result <= 12'b011100111000;
   21024: result <= 12'b011100111000;
   21025: result <= 12'b011100111000;
   21026: result <= 12'b011100111000;
   21027: result <= 12'b011100111000;
   21028: result <= 12'b011100111000;
   21029: result <= 12'b011100111000;
   21030: result <= 12'b011100111000;
   21031: result <= 12'b011100111000;
   21032: result <= 12'b011100110111;
   21033: result <= 12'b011100110111;
   21034: result <= 12'b011100110111;
   21035: result <= 12'b011100110111;
   21036: result <= 12'b011100110111;
   21037: result <= 12'b011100110111;
   21038: result <= 12'b011100110111;
   21039: result <= 12'b011100110111;
   21040: result <= 12'b011100110111;
   21041: result <= 12'b011100110111;
   21042: result <= 12'b011100110111;
   21043: result <= 12'b011100110111;
   21044: result <= 12'b011100110110;
   21045: result <= 12'b011100110110;
   21046: result <= 12'b011100110110;
   21047: result <= 12'b011100110110;
   21048: result <= 12'b011100110110;
   21049: result <= 12'b011100110110;
   21050: result <= 12'b011100110110;
   21051: result <= 12'b011100110110;
   21052: result <= 12'b011100110110;
   21053: result <= 12'b011100110110;
   21054: result <= 12'b011100110110;
   21055: result <= 12'b011100110110;
   21056: result <= 12'b011100110101;
   21057: result <= 12'b011100110101;
   21058: result <= 12'b011100110101;
   21059: result <= 12'b011100110101;
   21060: result <= 12'b011100110101;
   21061: result <= 12'b011100110101;
   21062: result <= 12'b011100110101;
   21063: result <= 12'b011100110101;
   21064: result <= 12'b011100110101;
   21065: result <= 12'b011100110101;
   21066: result <= 12'b011100110101;
   21067: result <= 12'b011100110101;
   21068: result <= 12'b011100110100;
   21069: result <= 12'b011100110100;
   21070: result <= 12'b011100110100;
   21071: result <= 12'b011100110100;
   21072: result <= 12'b011100110100;
   21073: result <= 12'b011100110100;
   21074: result <= 12'b011100110100;
   21075: result <= 12'b011100110100;
   21076: result <= 12'b011100110100;
   21077: result <= 12'b011100110100;
   21078: result <= 12'b011100110100;
   21079: result <= 12'b011100110100;
   21080: result <= 12'b011100110011;
   21081: result <= 12'b011100110011;
   21082: result <= 12'b011100110011;
   21083: result <= 12'b011100110011;
   21084: result <= 12'b011100110011;
   21085: result <= 12'b011100110011;
   21086: result <= 12'b011100110011;
   21087: result <= 12'b011100110011;
   21088: result <= 12'b011100110011;
   21089: result <= 12'b011100110011;
   21090: result <= 12'b011100110011;
   21091: result <= 12'b011100110010;
   21092: result <= 12'b011100110010;
   21093: result <= 12'b011100110010;
   21094: result <= 12'b011100110010;
   21095: result <= 12'b011100110010;
   21096: result <= 12'b011100110010;
   21097: result <= 12'b011100110010;
   21098: result <= 12'b011100110010;
   21099: result <= 12'b011100110010;
   21100: result <= 12'b011100110010;
   21101: result <= 12'b011100110010;
   21102: result <= 12'b011100110010;
   21103: result <= 12'b011100110001;
   21104: result <= 12'b011100110001;
   21105: result <= 12'b011100110001;
   21106: result <= 12'b011100110001;
   21107: result <= 12'b011100110001;
   21108: result <= 12'b011100110001;
   21109: result <= 12'b011100110001;
   21110: result <= 12'b011100110001;
   21111: result <= 12'b011100110001;
   21112: result <= 12'b011100110001;
   21113: result <= 12'b011100110001;
   21114: result <= 12'b011100110001;
   21115: result <= 12'b011100110000;
   21116: result <= 12'b011100110000;
   21117: result <= 12'b011100110000;
   21118: result <= 12'b011100110000;
   21119: result <= 12'b011100110000;
   21120: result <= 12'b011100110000;
   21121: result <= 12'b011100110000;
   21122: result <= 12'b011100110000;
   21123: result <= 12'b011100110000;
   21124: result <= 12'b011100110000;
   21125: result <= 12'b011100110000;
   21126: result <= 12'b011100101111;
   21127: result <= 12'b011100101111;
   21128: result <= 12'b011100101111;
   21129: result <= 12'b011100101111;
   21130: result <= 12'b011100101111;
   21131: result <= 12'b011100101111;
   21132: result <= 12'b011100101111;
   21133: result <= 12'b011100101111;
   21134: result <= 12'b011100101111;
   21135: result <= 12'b011100101111;
   21136: result <= 12'b011100101111;
   21137: result <= 12'b011100101111;
   21138: result <= 12'b011100101110;
   21139: result <= 12'b011100101110;
   21140: result <= 12'b011100101110;
   21141: result <= 12'b011100101110;
   21142: result <= 12'b011100101110;
   21143: result <= 12'b011100101110;
   21144: result <= 12'b011100101110;
   21145: result <= 12'b011100101110;
   21146: result <= 12'b011100101110;
   21147: result <= 12'b011100101110;
   21148: result <= 12'b011100101110;
   21149: result <= 12'b011100101101;
   21150: result <= 12'b011100101101;
   21151: result <= 12'b011100101101;
   21152: result <= 12'b011100101101;
   21153: result <= 12'b011100101101;
   21154: result <= 12'b011100101101;
   21155: result <= 12'b011100101101;
   21156: result <= 12'b011100101101;
   21157: result <= 12'b011100101101;
   21158: result <= 12'b011100101101;
   21159: result <= 12'b011100101101;
   21160: result <= 12'b011100101101;
   21161: result <= 12'b011100101100;
   21162: result <= 12'b011100101100;
   21163: result <= 12'b011100101100;
   21164: result <= 12'b011100101100;
   21165: result <= 12'b011100101100;
   21166: result <= 12'b011100101100;
   21167: result <= 12'b011100101100;
   21168: result <= 12'b011100101100;
   21169: result <= 12'b011100101100;
   21170: result <= 12'b011100101100;
   21171: result <= 12'b011100101100;
   21172: result <= 12'b011100101011;
   21173: result <= 12'b011100101011;
   21174: result <= 12'b011100101011;
   21175: result <= 12'b011100101011;
   21176: result <= 12'b011100101011;
   21177: result <= 12'b011100101011;
   21178: result <= 12'b011100101011;
   21179: result <= 12'b011100101011;
   21180: result <= 12'b011100101011;
   21181: result <= 12'b011100101011;
   21182: result <= 12'b011100101011;
   21183: result <= 12'b011100101011;
   21184: result <= 12'b011100101010;
   21185: result <= 12'b011100101010;
   21186: result <= 12'b011100101010;
   21187: result <= 12'b011100101010;
   21188: result <= 12'b011100101010;
   21189: result <= 12'b011100101010;
   21190: result <= 12'b011100101010;
   21191: result <= 12'b011100101010;
   21192: result <= 12'b011100101010;
   21193: result <= 12'b011100101010;
   21194: result <= 12'b011100101010;
   21195: result <= 12'b011100101001;
   21196: result <= 12'b011100101001;
   21197: result <= 12'b011100101001;
   21198: result <= 12'b011100101001;
   21199: result <= 12'b011100101001;
   21200: result <= 12'b011100101001;
   21201: result <= 12'b011100101001;
   21202: result <= 12'b011100101001;
   21203: result <= 12'b011100101001;
   21204: result <= 12'b011100101001;
   21205: result <= 12'b011100101001;
   21206: result <= 12'b011100101001;
   21207: result <= 12'b011100101000;
   21208: result <= 12'b011100101000;
   21209: result <= 12'b011100101000;
   21210: result <= 12'b011100101000;
   21211: result <= 12'b011100101000;
   21212: result <= 12'b011100101000;
   21213: result <= 12'b011100101000;
   21214: result <= 12'b011100101000;
   21215: result <= 12'b011100101000;
   21216: result <= 12'b011100101000;
   21217: result <= 12'b011100101000;
   21218: result <= 12'b011100100111;
   21219: result <= 12'b011100100111;
   21220: result <= 12'b011100100111;
   21221: result <= 12'b011100100111;
   21222: result <= 12'b011100100111;
   21223: result <= 12'b011100100111;
   21224: result <= 12'b011100100111;
   21225: result <= 12'b011100100111;
   21226: result <= 12'b011100100111;
   21227: result <= 12'b011100100111;
   21228: result <= 12'b011100100111;
   21229: result <= 12'b011100100110;
   21230: result <= 12'b011100100110;
   21231: result <= 12'b011100100110;
   21232: result <= 12'b011100100110;
   21233: result <= 12'b011100100110;
   21234: result <= 12'b011100100110;
   21235: result <= 12'b011100100110;
   21236: result <= 12'b011100100110;
   21237: result <= 12'b011100100110;
   21238: result <= 12'b011100100110;
   21239: result <= 12'b011100100110;
   21240: result <= 12'b011100100110;
   21241: result <= 12'b011100100101;
   21242: result <= 12'b011100100101;
   21243: result <= 12'b011100100101;
   21244: result <= 12'b011100100101;
   21245: result <= 12'b011100100101;
   21246: result <= 12'b011100100101;
   21247: result <= 12'b011100100101;
   21248: result <= 12'b011100100101;
   21249: result <= 12'b011100100101;
   21250: result <= 12'b011100100101;
   21251: result <= 12'b011100100101;
   21252: result <= 12'b011100100100;
   21253: result <= 12'b011100100100;
   21254: result <= 12'b011100100100;
   21255: result <= 12'b011100100100;
   21256: result <= 12'b011100100100;
   21257: result <= 12'b011100100100;
   21258: result <= 12'b011100100100;
   21259: result <= 12'b011100100100;
   21260: result <= 12'b011100100100;
   21261: result <= 12'b011100100100;
   21262: result <= 12'b011100100100;
   21263: result <= 12'b011100100011;
   21264: result <= 12'b011100100011;
   21265: result <= 12'b011100100011;
   21266: result <= 12'b011100100011;
   21267: result <= 12'b011100100011;
   21268: result <= 12'b011100100011;
   21269: result <= 12'b011100100011;
   21270: result <= 12'b011100100011;
   21271: result <= 12'b011100100011;
   21272: result <= 12'b011100100011;
   21273: result <= 12'b011100100011;
   21274: result <= 12'b011100100011;
   21275: result <= 12'b011100100010;
   21276: result <= 12'b011100100010;
   21277: result <= 12'b011100100010;
   21278: result <= 12'b011100100010;
   21279: result <= 12'b011100100010;
   21280: result <= 12'b011100100010;
   21281: result <= 12'b011100100010;
   21282: result <= 12'b011100100010;
   21283: result <= 12'b011100100010;
   21284: result <= 12'b011100100010;
   21285: result <= 12'b011100100010;
   21286: result <= 12'b011100100001;
   21287: result <= 12'b011100100001;
   21288: result <= 12'b011100100001;
   21289: result <= 12'b011100100001;
   21290: result <= 12'b011100100001;
   21291: result <= 12'b011100100001;
   21292: result <= 12'b011100100001;
   21293: result <= 12'b011100100001;
   21294: result <= 12'b011100100001;
   21295: result <= 12'b011100100001;
   21296: result <= 12'b011100100001;
   21297: result <= 12'b011100100000;
   21298: result <= 12'b011100100000;
   21299: result <= 12'b011100100000;
   21300: result <= 12'b011100100000;
   21301: result <= 12'b011100100000;
   21302: result <= 12'b011100100000;
   21303: result <= 12'b011100100000;
   21304: result <= 12'b011100100000;
   21305: result <= 12'b011100100000;
   21306: result <= 12'b011100100000;
   21307: result <= 12'b011100100000;
   21308: result <= 12'b011100011111;
   21309: result <= 12'b011100011111;
   21310: result <= 12'b011100011111;
   21311: result <= 12'b011100011111;
   21312: result <= 12'b011100011111;
   21313: result <= 12'b011100011111;
   21314: result <= 12'b011100011111;
   21315: result <= 12'b011100011111;
   21316: result <= 12'b011100011111;
   21317: result <= 12'b011100011111;
   21318: result <= 12'b011100011111;
   21319: result <= 12'b011100011111;
   21320: result <= 12'b011100011110;
   21321: result <= 12'b011100011110;
   21322: result <= 12'b011100011110;
   21323: result <= 12'b011100011110;
   21324: result <= 12'b011100011110;
   21325: result <= 12'b011100011110;
   21326: result <= 12'b011100011110;
   21327: result <= 12'b011100011110;
   21328: result <= 12'b011100011110;
   21329: result <= 12'b011100011110;
   21330: result <= 12'b011100011110;
   21331: result <= 12'b011100011101;
   21332: result <= 12'b011100011101;
   21333: result <= 12'b011100011101;
   21334: result <= 12'b011100011101;
   21335: result <= 12'b011100011101;
   21336: result <= 12'b011100011101;
   21337: result <= 12'b011100011101;
   21338: result <= 12'b011100011101;
   21339: result <= 12'b011100011101;
   21340: result <= 12'b011100011101;
   21341: result <= 12'b011100011101;
   21342: result <= 12'b011100011100;
   21343: result <= 12'b011100011100;
   21344: result <= 12'b011100011100;
   21345: result <= 12'b011100011100;
   21346: result <= 12'b011100011100;
   21347: result <= 12'b011100011100;
   21348: result <= 12'b011100011100;
   21349: result <= 12'b011100011100;
   21350: result <= 12'b011100011100;
   21351: result <= 12'b011100011100;
   21352: result <= 12'b011100011100;
   21353: result <= 12'b011100011011;
   21354: result <= 12'b011100011011;
   21355: result <= 12'b011100011011;
   21356: result <= 12'b011100011011;
   21357: result <= 12'b011100011011;
   21358: result <= 12'b011100011011;
   21359: result <= 12'b011100011011;
   21360: result <= 12'b011100011011;
   21361: result <= 12'b011100011011;
   21362: result <= 12'b011100011011;
   21363: result <= 12'b011100011011;
   21364: result <= 12'b011100011010;
   21365: result <= 12'b011100011010;
   21366: result <= 12'b011100011010;
   21367: result <= 12'b011100011010;
   21368: result <= 12'b011100011010;
   21369: result <= 12'b011100011010;
   21370: result <= 12'b011100011010;
   21371: result <= 12'b011100011010;
   21372: result <= 12'b011100011010;
   21373: result <= 12'b011100011010;
   21374: result <= 12'b011100011010;
   21375: result <= 12'b011100011001;
   21376: result <= 12'b011100011001;
   21377: result <= 12'b011100011001;
   21378: result <= 12'b011100011001;
   21379: result <= 12'b011100011001;
   21380: result <= 12'b011100011001;
   21381: result <= 12'b011100011001;
   21382: result <= 12'b011100011001;
   21383: result <= 12'b011100011001;
   21384: result <= 12'b011100011001;
   21385: result <= 12'b011100011001;
   21386: result <= 12'b011100011000;
   21387: result <= 12'b011100011000;
   21388: result <= 12'b011100011000;
   21389: result <= 12'b011100011000;
   21390: result <= 12'b011100011000;
   21391: result <= 12'b011100011000;
   21392: result <= 12'b011100011000;
   21393: result <= 12'b011100011000;
   21394: result <= 12'b011100011000;
   21395: result <= 12'b011100011000;
   21396: result <= 12'b011100011000;
   21397: result <= 12'b011100010111;
   21398: result <= 12'b011100010111;
   21399: result <= 12'b011100010111;
   21400: result <= 12'b011100010111;
   21401: result <= 12'b011100010111;
   21402: result <= 12'b011100010111;
   21403: result <= 12'b011100010111;
   21404: result <= 12'b011100010111;
   21405: result <= 12'b011100010111;
   21406: result <= 12'b011100010111;
   21407: result <= 12'b011100010111;
   21408: result <= 12'b011100010110;
   21409: result <= 12'b011100010110;
   21410: result <= 12'b011100010110;
   21411: result <= 12'b011100010110;
   21412: result <= 12'b011100010110;
   21413: result <= 12'b011100010110;
   21414: result <= 12'b011100010110;
   21415: result <= 12'b011100010110;
   21416: result <= 12'b011100010110;
   21417: result <= 12'b011100010110;
   21418: result <= 12'b011100010110;
   21419: result <= 12'b011100010101;
   21420: result <= 12'b011100010101;
   21421: result <= 12'b011100010101;
   21422: result <= 12'b011100010101;
   21423: result <= 12'b011100010101;
   21424: result <= 12'b011100010101;
   21425: result <= 12'b011100010101;
   21426: result <= 12'b011100010101;
   21427: result <= 12'b011100010101;
   21428: result <= 12'b011100010101;
   21429: result <= 12'b011100010101;
   21430: result <= 12'b011100010100;
   21431: result <= 12'b011100010100;
   21432: result <= 12'b011100010100;
   21433: result <= 12'b011100010100;
   21434: result <= 12'b011100010100;
   21435: result <= 12'b011100010100;
   21436: result <= 12'b011100010100;
   21437: result <= 12'b011100010100;
   21438: result <= 12'b011100010100;
   21439: result <= 12'b011100010100;
   21440: result <= 12'b011100010100;
   21441: result <= 12'b011100010011;
   21442: result <= 12'b011100010011;
   21443: result <= 12'b011100010011;
   21444: result <= 12'b011100010011;
   21445: result <= 12'b011100010011;
   21446: result <= 12'b011100010011;
   21447: result <= 12'b011100010011;
   21448: result <= 12'b011100010011;
   21449: result <= 12'b011100010011;
   21450: result <= 12'b011100010011;
   21451: result <= 12'b011100010011;
   21452: result <= 12'b011100010010;
   21453: result <= 12'b011100010010;
   21454: result <= 12'b011100010010;
   21455: result <= 12'b011100010010;
   21456: result <= 12'b011100010010;
   21457: result <= 12'b011100010010;
   21458: result <= 12'b011100010010;
   21459: result <= 12'b011100010010;
   21460: result <= 12'b011100010010;
   21461: result <= 12'b011100010010;
   21462: result <= 12'b011100010010;
   21463: result <= 12'b011100010001;
   21464: result <= 12'b011100010001;
   21465: result <= 12'b011100010001;
   21466: result <= 12'b011100010001;
   21467: result <= 12'b011100010001;
   21468: result <= 12'b011100010001;
   21469: result <= 12'b011100010001;
   21470: result <= 12'b011100010001;
   21471: result <= 12'b011100010001;
   21472: result <= 12'b011100010001;
   21473: result <= 12'b011100010001;
   21474: result <= 12'b011100010000;
   21475: result <= 12'b011100010000;
   21476: result <= 12'b011100010000;
   21477: result <= 12'b011100010000;
   21478: result <= 12'b011100010000;
   21479: result <= 12'b011100010000;
   21480: result <= 12'b011100010000;
   21481: result <= 12'b011100010000;
   21482: result <= 12'b011100010000;
   21483: result <= 12'b011100010000;
   21484: result <= 12'b011100010000;
   21485: result <= 12'b011100001111;
   21486: result <= 12'b011100001111;
   21487: result <= 12'b011100001111;
   21488: result <= 12'b011100001111;
   21489: result <= 12'b011100001111;
   21490: result <= 12'b011100001111;
   21491: result <= 12'b011100001111;
   21492: result <= 12'b011100001111;
   21493: result <= 12'b011100001111;
   21494: result <= 12'b011100001111;
   21495: result <= 12'b011100001111;
   21496: result <= 12'b011100001110;
   21497: result <= 12'b011100001110;
   21498: result <= 12'b011100001110;
   21499: result <= 12'b011100001110;
   21500: result <= 12'b011100001110;
   21501: result <= 12'b011100001110;
   21502: result <= 12'b011100001110;
   21503: result <= 12'b011100001110;
   21504: result <= 12'b011100001110;
   21505: result <= 12'b011100001110;
   21506: result <= 12'b011100001101;
   21507: result <= 12'b011100001101;
   21508: result <= 12'b011100001101;
   21509: result <= 12'b011100001101;
   21510: result <= 12'b011100001101;
   21511: result <= 12'b011100001101;
   21512: result <= 12'b011100001101;
   21513: result <= 12'b011100001101;
   21514: result <= 12'b011100001101;
   21515: result <= 12'b011100001101;
   21516: result <= 12'b011100001101;
   21517: result <= 12'b011100001100;
   21518: result <= 12'b011100001100;
   21519: result <= 12'b011100001100;
   21520: result <= 12'b011100001100;
   21521: result <= 12'b011100001100;
   21522: result <= 12'b011100001100;
   21523: result <= 12'b011100001100;
   21524: result <= 12'b011100001100;
   21525: result <= 12'b011100001100;
   21526: result <= 12'b011100001100;
   21527: result <= 12'b011100001100;
   21528: result <= 12'b011100001011;
   21529: result <= 12'b011100001011;
   21530: result <= 12'b011100001011;
   21531: result <= 12'b011100001011;
   21532: result <= 12'b011100001011;
   21533: result <= 12'b011100001011;
   21534: result <= 12'b011100001011;
   21535: result <= 12'b011100001011;
   21536: result <= 12'b011100001011;
   21537: result <= 12'b011100001011;
   21538: result <= 12'b011100001011;
   21539: result <= 12'b011100001010;
   21540: result <= 12'b011100001010;
   21541: result <= 12'b011100001010;
   21542: result <= 12'b011100001010;
   21543: result <= 12'b011100001010;
   21544: result <= 12'b011100001010;
   21545: result <= 12'b011100001010;
   21546: result <= 12'b011100001010;
   21547: result <= 12'b011100001010;
   21548: result <= 12'b011100001010;
   21549: result <= 12'b011100001001;
   21550: result <= 12'b011100001001;
   21551: result <= 12'b011100001001;
   21552: result <= 12'b011100001001;
   21553: result <= 12'b011100001001;
   21554: result <= 12'b011100001001;
   21555: result <= 12'b011100001001;
   21556: result <= 12'b011100001001;
   21557: result <= 12'b011100001001;
   21558: result <= 12'b011100001001;
   21559: result <= 12'b011100001001;
   21560: result <= 12'b011100001000;
   21561: result <= 12'b011100001000;
   21562: result <= 12'b011100001000;
   21563: result <= 12'b011100001000;
   21564: result <= 12'b011100001000;
   21565: result <= 12'b011100001000;
   21566: result <= 12'b011100001000;
   21567: result <= 12'b011100001000;
   21568: result <= 12'b011100001000;
   21569: result <= 12'b011100001000;
   21570: result <= 12'b011100001000;
   21571: result <= 12'b011100000111;
   21572: result <= 12'b011100000111;
   21573: result <= 12'b011100000111;
   21574: result <= 12'b011100000111;
   21575: result <= 12'b011100000111;
   21576: result <= 12'b011100000111;
   21577: result <= 12'b011100000111;
   21578: result <= 12'b011100000111;
   21579: result <= 12'b011100000111;
   21580: result <= 12'b011100000111;
   21581: result <= 12'b011100000110;
   21582: result <= 12'b011100000110;
   21583: result <= 12'b011100000110;
   21584: result <= 12'b011100000110;
   21585: result <= 12'b011100000110;
   21586: result <= 12'b011100000110;
   21587: result <= 12'b011100000110;
   21588: result <= 12'b011100000110;
   21589: result <= 12'b011100000110;
   21590: result <= 12'b011100000110;
   21591: result <= 12'b011100000110;
   21592: result <= 12'b011100000101;
   21593: result <= 12'b011100000101;
   21594: result <= 12'b011100000101;
   21595: result <= 12'b011100000101;
   21596: result <= 12'b011100000101;
   21597: result <= 12'b011100000101;
   21598: result <= 12'b011100000101;
   21599: result <= 12'b011100000101;
   21600: result <= 12'b011100000101;
   21601: result <= 12'b011100000101;
   21602: result <= 12'b011100000101;
   21603: result <= 12'b011100000100;
   21604: result <= 12'b011100000100;
   21605: result <= 12'b011100000100;
   21606: result <= 12'b011100000100;
   21607: result <= 12'b011100000100;
   21608: result <= 12'b011100000100;
   21609: result <= 12'b011100000100;
   21610: result <= 12'b011100000100;
   21611: result <= 12'b011100000100;
   21612: result <= 12'b011100000100;
   21613: result <= 12'b011100000011;
   21614: result <= 12'b011100000011;
   21615: result <= 12'b011100000011;
   21616: result <= 12'b011100000011;
   21617: result <= 12'b011100000011;
   21618: result <= 12'b011100000011;
   21619: result <= 12'b011100000011;
   21620: result <= 12'b011100000011;
   21621: result <= 12'b011100000011;
   21622: result <= 12'b011100000011;
   21623: result <= 12'b011100000011;
   21624: result <= 12'b011100000010;
   21625: result <= 12'b011100000010;
   21626: result <= 12'b011100000010;
   21627: result <= 12'b011100000010;
   21628: result <= 12'b011100000010;
   21629: result <= 12'b011100000010;
   21630: result <= 12'b011100000010;
   21631: result <= 12'b011100000010;
   21632: result <= 12'b011100000010;
   21633: result <= 12'b011100000010;
   21634: result <= 12'b011100000010;
   21635: result <= 12'b011100000001;
   21636: result <= 12'b011100000001;
   21637: result <= 12'b011100000001;
   21638: result <= 12'b011100000001;
   21639: result <= 12'b011100000001;
   21640: result <= 12'b011100000001;
   21641: result <= 12'b011100000001;
   21642: result <= 12'b011100000001;
   21643: result <= 12'b011100000001;
   21644: result <= 12'b011100000001;
   21645: result <= 12'b011100000000;
   21646: result <= 12'b011100000000;
   21647: result <= 12'b011100000000;
   21648: result <= 12'b011100000000;
   21649: result <= 12'b011100000000;
   21650: result <= 12'b011100000000;
   21651: result <= 12'b011100000000;
   21652: result <= 12'b011100000000;
   21653: result <= 12'b011100000000;
   21654: result <= 12'b011100000000;
   21655: result <= 12'b011100000000;
   21656: result <= 12'b011011111111;
   21657: result <= 12'b011011111111;
   21658: result <= 12'b011011111111;
   21659: result <= 12'b011011111111;
   21660: result <= 12'b011011111111;
   21661: result <= 12'b011011111111;
   21662: result <= 12'b011011111111;
   21663: result <= 12'b011011111111;
   21664: result <= 12'b011011111111;
   21665: result <= 12'b011011111111;
   21666: result <= 12'b011011111110;
   21667: result <= 12'b011011111110;
   21668: result <= 12'b011011111110;
   21669: result <= 12'b011011111110;
   21670: result <= 12'b011011111110;
   21671: result <= 12'b011011111110;
   21672: result <= 12'b011011111110;
   21673: result <= 12'b011011111110;
   21674: result <= 12'b011011111110;
   21675: result <= 12'b011011111110;
   21676: result <= 12'b011011111110;
   21677: result <= 12'b011011111101;
   21678: result <= 12'b011011111101;
   21679: result <= 12'b011011111101;
   21680: result <= 12'b011011111101;
   21681: result <= 12'b011011111101;
   21682: result <= 12'b011011111101;
   21683: result <= 12'b011011111101;
   21684: result <= 12'b011011111101;
   21685: result <= 12'b011011111101;
   21686: result <= 12'b011011111101;
   21687: result <= 12'b011011111100;
   21688: result <= 12'b011011111100;
   21689: result <= 12'b011011111100;
   21690: result <= 12'b011011111100;
   21691: result <= 12'b011011111100;
   21692: result <= 12'b011011111100;
   21693: result <= 12'b011011111100;
   21694: result <= 12'b011011111100;
   21695: result <= 12'b011011111100;
   21696: result <= 12'b011011111100;
   21697: result <= 12'b011011111100;
   21698: result <= 12'b011011111011;
   21699: result <= 12'b011011111011;
   21700: result <= 12'b011011111011;
   21701: result <= 12'b011011111011;
   21702: result <= 12'b011011111011;
   21703: result <= 12'b011011111011;
   21704: result <= 12'b011011111011;
   21705: result <= 12'b011011111011;
   21706: result <= 12'b011011111011;
   21707: result <= 12'b011011111011;
   21708: result <= 12'b011011111010;
   21709: result <= 12'b011011111010;
   21710: result <= 12'b011011111010;
   21711: result <= 12'b011011111010;
   21712: result <= 12'b011011111010;
   21713: result <= 12'b011011111010;
   21714: result <= 12'b011011111010;
   21715: result <= 12'b011011111010;
   21716: result <= 12'b011011111010;
   21717: result <= 12'b011011111010;
   21718: result <= 12'b011011111001;
   21719: result <= 12'b011011111001;
   21720: result <= 12'b011011111001;
   21721: result <= 12'b011011111001;
   21722: result <= 12'b011011111001;
   21723: result <= 12'b011011111001;
   21724: result <= 12'b011011111001;
   21725: result <= 12'b011011111001;
   21726: result <= 12'b011011111001;
   21727: result <= 12'b011011111001;
   21728: result <= 12'b011011111001;
   21729: result <= 12'b011011111000;
   21730: result <= 12'b011011111000;
   21731: result <= 12'b011011111000;
   21732: result <= 12'b011011111000;
   21733: result <= 12'b011011111000;
   21734: result <= 12'b011011111000;
   21735: result <= 12'b011011111000;
   21736: result <= 12'b011011111000;
   21737: result <= 12'b011011111000;
   21738: result <= 12'b011011111000;
   21739: result <= 12'b011011110111;
   21740: result <= 12'b011011110111;
   21741: result <= 12'b011011110111;
   21742: result <= 12'b011011110111;
   21743: result <= 12'b011011110111;
   21744: result <= 12'b011011110111;
   21745: result <= 12'b011011110111;
   21746: result <= 12'b011011110111;
   21747: result <= 12'b011011110111;
   21748: result <= 12'b011011110111;
   21749: result <= 12'b011011110111;
   21750: result <= 12'b011011110110;
   21751: result <= 12'b011011110110;
   21752: result <= 12'b011011110110;
   21753: result <= 12'b011011110110;
   21754: result <= 12'b011011110110;
   21755: result <= 12'b011011110110;
   21756: result <= 12'b011011110110;
   21757: result <= 12'b011011110110;
   21758: result <= 12'b011011110110;
   21759: result <= 12'b011011110110;
   21760: result <= 12'b011011110101;
   21761: result <= 12'b011011110101;
   21762: result <= 12'b011011110101;
   21763: result <= 12'b011011110101;
   21764: result <= 12'b011011110101;
   21765: result <= 12'b011011110101;
   21766: result <= 12'b011011110101;
   21767: result <= 12'b011011110101;
   21768: result <= 12'b011011110101;
   21769: result <= 12'b011011110101;
   21770: result <= 12'b011011110100;
   21771: result <= 12'b011011110100;
   21772: result <= 12'b011011110100;
   21773: result <= 12'b011011110100;
   21774: result <= 12'b011011110100;
   21775: result <= 12'b011011110100;
   21776: result <= 12'b011011110100;
   21777: result <= 12'b011011110100;
   21778: result <= 12'b011011110100;
   21779: result <= 12'b011011110100;
   21780: result <= 12'b011011110011;
   21781: result <= 12'b011011110011;
   21782: result <= 12'b011011110011;
   21783: result <= 12'b011011110011;
   21784: result <= 12'b011011110011;
   21785: result <= 12'b011011110011;
   21786: result <= 12'b011011110011;
   21787: result <= 12'b011011110011;
   21788: result <= 12'b011011110011;
   21789: result <= 12'b011011110011;
   21790: result <= 12'b011011110011;
   21791: result <= 12'b011011110010;
   21792: result <= 12'b011011110010;
   21793: result <= 12'b011011110010;
   21794: result <= 12'b011011110010;
   21795: result <= 12'b011011110010;
   21796: result <= 12'b011011110010;
   21797: result <= 12'b011011110010;
   21798: result <= 12'b011011110010;
   21799: result <= 12'b011011110010;
   21800: result <= 12'b011011110010;
   21801: result <= 12'b011011110001;
   21802: result <= 12'b011011110001;
   21803: result <= 12'b011011110001;
   21804: result <= 12'b011011110001;
   21805: result <= 12'b011011110001;
   21806: result <= 12'b011011110001;
   21807: result <= 12'b011011110001;
   21808: result <= 12'b011011110001;
   21809: result <= 12'b011011110001;
   21810: result <= 12'b011011110001;
   21811: result <= 12'b011011110000;
   21812: result <= 12'b011011110000;
   21813: result <= 12'b011011110000;
   21814: result <= 12'b011011110000;
   21815: result <= 12'b011011110000;
   21816: result <= 12'b011011110000;
   21817: result <= 12'b011011110000;
   21818: result <= 12'b011011110000;
   21819: result <= 12'b011011110000;
   21820: result <= 12'b011011110000;
   21821: result <= 12'b011011110000;
   21822: result <= 12'b011011101111;
   21823: result <= 12'b011011101111;
   21824: result <= 12'b011011101111;
   21825: result <= 12'b011011101111;
   21826: result <= 12'b011011101111;
   21827: result <= 12'b011011101111;
   21828: result <= 12'b011011101111;
   21829: result <= 12'b011011101111;
   21830: result <= 12'b011011101111;
   21831: result <= 12'b011011101111;
   21832: result <= 12'b011011101110;
   21833: result <= 12'b011011101110;
   21834: result <= 12'b011011101110;
   21835: result <= 12'b011011101110;
   21836: result <= 12'b011011101110;
   21837: result <= 12'b011011101110;
   21838: result <= 12'b011011101110;
   21839: result <= 12'b011011101110;
   21840: result <= 12'b011011101110;
   21841: result <= 12'b011011101110;
   21842: result <= 12'b011011101101;
   21843: result <= 12'b011011101101;
   21844: result <= 12'b011011101101;
   21845: result <= 12'b011011101101;
   21846: result <= 12'b011011101101;
   21847: result <= 12'b011011101101;
   21848: result <= 12'b011011101101;
   21849: result <= 12'b011011101101;
   21850: result <= 12'b011011101101;
   21851: result <= 12'b011011101101;
   21852: result <= 12'b011011101100;
   21853: result <= 12'b011011101100;
   21854: result <= 12'b011011101100;
   21855: result <= 12'b011011101100;
   21856: result <= 12'b011011101100;
   21857: result <= 12'b011011101100;
   21858: result <= 12'b011011101100;
   21859: result <= 12'b011011101100;
   21860: result <= 12'b011011101100;
   21861: result <= 12'b011011101100;
   21862: result <= 12'b011011101011;
   21863: result <= 12'b011011101011;
   21864: result <= 12'b011011101011;
   21865: result <= 12'b011011101011;
   21866: result <= 12'b011011101011;
   21867: result <= 12'b011011101011;
   21868: result <= 12'b011011101011;
   21869: result <= 12'b011011101011;
   21870: result <= 12'b011011101011;
   21871: result <= 12'b011011101011;
   21872: result <= 12'b011011101010;
   21873: result <= 12'b011011101010;
   21874: result <= 12'b011011101010;
   21875: result <= 12'b011011101010;
   21876: result <= 12'b011011101010;
   21877: result <= 12'b011011101010;
   21878: result <= 12'b011011101010;
   21879: result <= 12'b011011101010;
   21880: result <= 12'b011011101010;
   21881: result <= 12'b011011101010;
   21882: result <= 12'b011011101010;
   21883: result <= 12'b011011101001;
   21884: result <= 12'b011011101001;
   21885: result <= 12'b011011101001;
   21886: result <= 12'b011011101001;
   21887: result <= 12'b011011101001;
   21888: result <= 12'b011011101001;
   21889: result <= 12'b011011101001;
   21890: result <= 12'b011011101001;
   21891: result <= 12'b011011101001;
   21892: result <= 12'b011011101001;
   21893: result <= 12'b011011101000;
   21894: result <= 12'b011011101000;
   21895: result <= 12'b011011101000;
   21896: result <= 12'b011011101000;
   21897: result <= 12'b011011101000;
   21898: result <= 12'b011011101000;
   21899: result <= 12'b011011101000;
   21900: result <= 12'b011011101000;
   21901: result <= 12'b011011101000;
   21902: result <= 12'b011011101000;
   21903: result <= 12'b011011100111;
   21904: result <= 12'b011011100111;
   21905: result <= 12'b011011100111;
   21906: result <= 12'b011011100111;
   21907: result <= 12'b011011100111;
   21908: result <= 12'b011011100111;
   21909: result <= 12'b011011100111;
   21910: result <= 12'b011011100111;
   21911: result <= 12'b011011100111;
   21912: result <= 12'b011011100111;
   21913: result <= 12'b011011100110;
   21914: result <= 12'b011011100110;
   21915: result <= 12'b011011100110;
   21916: result <= 12'b011011100110;
   21917: result <= 12'b011011100110;
   21918: result <= 12'b011011100110;
   21919: result <= 12'b011011100110;
   21920: result <= 12'b011011100110;
   21921: result <= 12'b011011100110;
   21922: result <= 12'b011011100110;
   21923: result <= 12'b011011100101;
   21924: result <= 12'b011011100101;
   21925: result <= 12'b011011100101;
   21926: result <= 12'b011011100101;
   21927: result <= 12'b011011100101;
   21928: result <= 12'b011011100101;
   21929: result <= 12'b011011100101;
   21930: result <= 12'b011011100101;
   21931: result <= 12'b011011100101;
   21932: result <= 12'b011011100101;
   21933: result <= 12'b011011100100;
   21934: result <= 12'b011011100100;
   21935: result <= 12'b011011100100;
   21936: result <= 12'b011011100100;
   21937: result <= 12'b011011100100;
   21938: result <= 12'b011011100100;
   21939: result <= 12'b011011100100;
   21940: result <= 12'b011011100100;
   21941: result <= 12'b011011100100;
   21942: result <= 12'b011011100100;
   21943: result <= 12'b011011100011;
   21944: result <= 12'b011011100011;
   21945: result <= 12'b011011100011;
   21946: result <= 12'b011011100011;
   21947: result <= 12'b011011100011;
   21948: result <= 12'b011011100011;
   21949: result <= 12'b011011100011;
   21950: result <= 12'b011011100011;
   21951: result <= 12'b011011100011;
   21952: result <= 12'b011011100011;
   21953: result <= 12'b011011100010;
   21954: result <= 12'b011011100010;
   21955: result <= 12'b011011100010;
   21956: result <= 12'b011011100010;
   21957: result <= 12'b011011100010;
   21958: result <= 12'b011011100010;
   21959: result <= 12'b011011100010;
   21960: result <= 12'b011011100010;
   21961: result <= 12'b011011100010;
   21962: result <= 12'b011011100010;
   21963: result <= 12'b011011100001;
   21964: result <= 12'b011011100001;
   21965: result <= 12'b011011100001;
   21966: result <= 12'b011011100001;
   21967: result <= 12'b011011100001;
   21968: result <= 12'b011011100001;
   21969: result <= 12'b011011100001;
   21970: result <= 12'b011011100001;
   21971: result <= 12'b011011100001;
   21972: result <= 12'b011011100001;
   21973: result <= 12'b011011100000;
   21974: result <= 12'b011011100000;
   21975: result <= 12'b011011100000;
   21976: result <= 12'b011011100000;
   21977: result <= 12'b011011100000;
   21978: result <= 12'b011011100000;
   21979: result <= 12'b011011100000;
   21980: result <= 12'b011011100000;
   21981: result <= 12'b011011100000;
   21982: result <= 12'b011011100000;
   21983: result <= 12'b011011011111;
   21984: result <= 12'b011011011111;
   21985: result <= 12'b011011011111;
   21986: result <= 12'b011011011111;
   21987: result <= 12'b011011011111;
   21988: result <= 12'b011011011111;
   21989: result <= 12'b011011011111;
   21990: result <= 12'b011011011111;
   21991: result <= 12'b011011011111;
   21992: result <= 12'b011011011111;
   21993: result <= 12'b011011011110;
   21994: result <= 12'b011011011110;
   21995: result <= 12'b011011011110;
   21996: result <= 12'b011011011110;
   21997: result <= 12'b011011011110;
   21998: result <= 12'b011011011110;
   21999: result <= 12'b011011011110;
   22000: result <= 12'b011011011110;
   22001: result <= 12'b011011011110;
   22002: result <= 12'b011011011110;
   22003: result <= 12'b011011011101;
   22004: result <= 12'b011011011101;
   22005: result <= 12'b011011011101;
   22006: result <= 12'b011011011101;
   22007: result <= 12'b011011011101;
   22008: result <= 12'b011011011101;
   22009: result <= 12'b011011011101;
   22010: result <= 12'b011011011101;
   22011: result <= 12'b011011011101;
   22012: result <= 12'b011011011101;
   22013: result <= 12'b011011011100;
   22014: result <= 12'b011011011100;
   22015: result <= 12'b011011011100;
   22016: result <= 12'b011011011100;
   22017: result <= 12'b011011011100;
   22018: result <= 12'b011011011100;
   22019: result <= 12'b011011011100;
   22020: result <= 12'b011011011100;
   22021: result <= 12'b011011011100;
   22022: result <= 12'b011011011100;
   22023: result <= 12'b011011011011;
   22024: result <= 12'b011011011011;
   22025: result <= 12'b011011011011;
   22026: result <= 12'b011011011011;
   22027: result <= 12'b011011011011;
   22028: result <= 12'b011011011011;
   22029: result <= 12'b011011011011;
   22030: result <= 12'b011011011011;
   22031: result <= 12'b011011011011;
   22032: result <= 12'b011011011011;
   22033: result <= 12'b011011011010;
   22034: result <= 12'b011011011010;
   22035: result <= 12'b011011011010;
   22036: result <= 12'b011011011010;
   22037: result <= 12'b011011011010;
   22038: result <= 12'b011011011010;
   22039: result <= 12'b011011011010;
   22040: result <= 12'b011011011010;
   22041: result <= 12'b011011011010;
   22042: result <= 12'b011011011001;
   22043: result <= 12'b011011011001;
   22044: result <= 12'b011011011001;
   22045: result <= 12'b011011011001;
   22046: result <= 12'b011011011001;
   22047: result <= 12'b011011011001;
   22048: result <= 12'b011011011001;
   22049: result <= 12'b011011011001;
   22050: result <= 12'b011011011001;
   22051: result <= 12'b011011011001;
   22052: result <= 12'b011011011000;
   22053: result <= 12'b011011011000;
   22054: result <= 12'b011011011000;
   22055: result <= 12'b011011011000;
   22056: result <= 12'b011011011000;
   22057: result <= 12'b011011011000;
   22058: result <= 12'b011011011000;
   22059: result <= 12'b011011011000;
   22060: result <= 12'b011011011000;
   22061: result <= 12'b011011011000;
   22062: result <= 12'b011011010111;
   22063: result <= 12'b011011010111;
   22064: result <= 12'b011011010111;
   22065: result <= 12'b011011010111;
   22066: result <= 12'b011011010111;
   22067: result <= 12'b011011010111;
   22068: result <= 12'b011011010111;
   22069: result <= 12'b011011010111;
   22070: result <= 12'b011011010111;
   22071: result <= 12'b011011010111;
   22072: result <= 12'b011011010110;
   22073: result <= 12'b011011010110;
   22074: result <= 12'b011011010110;
   22075: result <= 12'b011011010110;
   22076: result <= 12'b011011010110;
   22077: result <= 12'b011011010110;
   22078: result <= 12'b011011010110;
   22079: result <= 12'b011011010110;
   22080: result <= 12'b011011010110;
   22081: result <= 12'b011011010110;
   22082: result <= 12'b011011010101;
   22083: result <= 12'b011011010101;
   22084: result <= 12'b011011010101;
   22085: result <= 12'b011011010101;
   22086: result <= 12'b011011010101;
   22087: result <= 12'b011011010101;
   22088: result <= 12'b011011010101;
   22089: result <= 12'b011011010101;
   22090: result <= 12'b011011010101;
   22091: result <= 12'b011011010101;
   22092: result <= 12'b011011010100;
   22093: result <= 12'b011011010100;
   22094: result <= 12'b011011010100;
   22095: result <= 12'b011011010100;
   22096: result <= 12'b011011010100;
   22097: result <= 12'b011011010100;
   22098: result <= 12'b011011010100;
   22099: result <= 12'b011011010100;
   22100: result <= 12'b011011010100;
   22101: result <= 12'b011011010011;
   22102: result <= 12'b011011010011;
   22103: result <= 12'b011011010011;
   22104: result <= 12'b011011010011;
   22105: result <= 12'b011011010011;
   22106: result <= 12'b011011010011;
   22107: result <= 12'b011011010011;
   22108: result <= 12'b011011010011;
   22109: result <= 12'b011011010011;
   22110: result <= 12'b011011010011;
   22111: result <= 12'b011011010010;
   22112: result <= 12'b011011010010;
   22113: result <= 12'b011011010010;
   22114: result <= 12'b011011010010;
   22115: result <= 12'b011011010010;
   22116: result <= 12'b011011010010;
   22117: result <= 12'b011011010010;
   22118: result <= 12'b011011010010;
   22119: result <= 12'b011011010010;
   22120: result <= 12'b011011010010;
   22121: result <= 12'b011011010001;
   22122: result <= 12'b011011010001;
   22123: result <= 12'b011011010001;
   22124: result <= 12'b011011010001;
   22125: result <= 12'b011011010001;
   22126: result <= 12'b011011010001;
   22127: result <= 12'b011011010001;
   22128: result <= 12'b011011010001;
   22129: result <= 12'b011011010001;
   22130: result <= 12'b011011010001;
   22131: result <= 12'b011011010000;
   22132: result <= 12'b011011010000;
   22133: result <= 12'b011011010000;
   22134: result <= 12'b011011010000;
   22135: result <= 12'b011011010000;
   22136: result <= 12'b011011010000;
   22137: result <= 12'b011011010000;
   22138: result <= 12'b011011010000;
   22139: result <= 12'b011011010000;
   22140: result <= 12'b011011001111;
   22141: result <= 12'b011011001111;
   22142: result <= 12'b011011001111;
   22143: result <= 12'b011011001111;
   22144: result <= 12'b011011001111;
   22145: result <= 12'b011011001111;
   22146: result <= 12'b011011001111;
   22147: result <= 12'b011011001111;
   22148: result <= 12'b011011001111;
   22149: result <= 12'b011011001111;
   22150: result <= 12'b011011001110;
   22151: result <= 12'b011011001110;
   22152: result <= 12'b011011001110;
   22153: result <= 12'b011011001110;
   22154: result <= 12'b011011001110;
   22155: result <= 12'b011011001110;
   22156: result <= 12'b011011001110;
   22157: result <= 12'b011011001110;
   22158: result <= 12'b011011001110;
   22159: result <= 12'b011011001110;
   22160: result <= 12'b011011001101;
   22161: result <= 12'b011011001101;
   22162: result <= 12'b011011001101;
   22163: result <= 12'b011011001101;
   22164: result <= 12'b011011001101;
   22165: result <= 12'b011011001101;
   22166: result <= 12'b011011001101;
   22167: result <= 12'b011011001101;
   22168: result <= 12'b011011001101;
   22169: result <= 12'b011011001100;
   22170: result <= 12'b011011001100;
   22171: result <= 12'b011011001100;
   22172: result <= 12'b011011001100;
   22173: result <= 12'b011011001100;
   22174: result <= 12'b011011001100;
   22175: result <= 12'b011011001100;
   22176: result <= 12'b011011001100;
   22177: result <= 12'b011011001100;
   22178: result <= 12'b011011001100;
   22179: result <= 12'b011011001011;
   22180: result <= 12'b011011001011;
   22181: result <= 12'b011011001011;
   22182: result <= 12'b011011001011;
   22183: result <= 12'b011011001011;
   22184: result <= 12'b011011001011;
   22185: result <= 12'b011011001011;
   22186: result <= 12'b011011001011;
   22187: result <= 12'b011011001011;
   22188: result <= 12'b011011001011;
   22189: result <= 12'b011011001010;
   22190: result <= 12'b011011001010;
   22191: result <= 12'b011011001010;
   22192: result <= 12'b011011001010;
   22193: result <= 12'b011011001010;
   22194: result <= 12'b011011001010;
   22195: result <= 12'b011011001010;
   22196: result <= 12'b011011001010;
   22197: result <= 12'b011011001010;
   22198: result <= 12'b011011001001;
   22199: result <= 12'b011011001001;
   22200: result <= 12'b011011001001;
   22201: result <= 12'b011011001001;
   22202: result <= 12'b011011001001;
   22203: result <= 12'b011011001001;
   22204: result <= 12'b011011001001;
   22205: result <= 12'b011011001001;
   22206: result <= 12'b011011001001;
   22207: result <= 12'b011011001001;
   22208: result <= 12'b011011001000;
   22209: result <= 12'b011011001000;
   22210: result <= 12'b011011001000;
   22211: result <= 12'b011011001000;
   22212: result <= 12'b011011001000;
   22213: result <= 12'b011011001000;
   22214: result <= 12'b011011001000;
   22215: result <= 12'b011011001000;
   22216: result <= 12'b011011001000;
   22217: result <= 12'b011011001000;
   22218: result <= 12'b011011000111;
   22219: result <= 12'b011011000111;
   22220: result <= 12'b011011000111;
   22221: result <= 12'b011011000111;
   22222: result <= 12'b011011000111;
   22223: result <= 12'b011011000111;
   22224: result <= 12'b011011000111;
   22225: result <= 12'b011011000111;
   22226: result <= 12'b011011000111;
   22227: result <= 12'b011011000110;
   22228: result <= 12'b011011000110;
   22229: result <= 12'b011011000110;
   22230: result <= 12'b011011000110;
   22231: result <= 12'b011011000110;
   22232: result <= 12'b011011000110;
   22233: result <= 12'b011011000110;
   22234: result <= 12'b011011000110;
   22235: result <= 12'b011011000110;
   22236: result <= 12'b011011000110;
   22237: result <= 12'b011011000101;
   22238: result <= 12'b011011000101;
   22239: result <= 12'b011011000101;
   22240: result <= 12'b011011000101;
   22241: result <= 12'b011011000101;
   22242: result <= 12'b011011000101;
   22243: result <= 12'b011011000101;
   22244: result <= 12'b011011000101;
   22245: result <= 12'b011011000101;
   22246: result <= 12'b011011000100;
   22247: result <= 12'b011011000100;
   22248: result <= 12'b011011000100;
   22249: result <= 12'b011011000100;
   22250: result <= 12'b011011000100;
   22251: result <= 12'b011011000100;
   22252: result <= 12'b011011000100;
   22253: result <= 12'b011011000100;
   22254: result <= 12'b011011000100;
   22255: result <= 12'b011011000100;
   22256: result <= 12'b011011000011;
   22257: result <= 12'b011011000011;
   22258: result <= 12'b011011000011;
   22259: result <= 12'b011011000011;
   22260: result <= 12'b011011000011;
   22261: result <= 12'b011011000011;
   22262: result <= 12'b011011000011;
   22263: result <= 12'b011011000011;
   22264: result <= 12'b011011000011;
   22265: result <= 12'b011011000010;
   22266: result <= 12'b011011000010;
   22267: result <= 12'b011011000010;
   22268: result <= 12'b011011000010;
   22269: result <= 12'b011011000010;
   22270: result <= 12'b011011000010;
   22271: result <= 12'b011011000010;
   22272: result <= 12'b011011000010;
   22273: result <= 12'b011011000010;
   22274: result <= 12'b011011000010;
   22275: result <= 12'b011011000001;
   22276: result <= 12'b011011000001;
   22277: result <= 12'b011011000001;
   22278: result <= 12'b011011000001;
   22279: result <= 12'b011011000001;
   22280: result <= 12'b011011000001;
   22281: result <= 12'b011011000001;
   22282: result <= 12'b011011000001;
   22283: result <= 12'b011011000001;
   22284: result <= 12'b011011000000;
   22285: result <= 12'b011011000000;
   22286: result <= 12'b011011000000;
   22287: result <= 12'b011011000000;
   22288: result <= 12'b011011000000;
   22289: result <= 12'b011011000000;
   22290: result <= 12'b011011000000;
   22291: result <= 12'b011011000000;
   22292: result <= 12'b011011000000;
   22293: result <= 12'b011011000000;
   22294: result <= 12'b011010111111;
   22295: result <= 12'b011010111111;
   22296: result <= 12'b011010111111;
   22297: result <= 12'b011010111111;
   22298: result <= 12'b011010111111;
   22299: result <= 12'b011010111111;
   22300: result <= 12'b011010111111;
   22301: result <= 12'b011010111111;
   22302: result <= 12'b011010111111;
   22303: result <= 12'b011010111110;
   22304: result <= 12'b011010111110;
   22305: result <= 12'b011010111110;
   22306: result <= 12'b011010111110;
   22307: result <= 12'b011010111110;
   22308: result <= 12'b011010111110;
   22309: result <= 12'b011010111110;
   22310: result <= 12'b011010111110;
   22311: result <= 12'b011010111110;
   22312: result <= 12'b011010111110;
   22313: result <= 12'b011010111101;
   22314: result <= 12'b011010111101;
   22315: result <= 12'b011010111101;
   22316: result <= 12'b011010111101;
   22317: result <= 12'b011010111101;
   22318: result <= 12'b011010111101;
   22319: result <= 12'b011010111101;
   22320: result <= 12'b011010111101;
   22321: result <= 12'b011010111101;
   22322: result <= 12'b011010111100;
   22323: result <= 12'b011010111100;
   22324: result <= 12'b011010111100;
   22325: result <= 12'b011010111100;
   22326: result <= 12'b011010111100;
   22327: result <= 12'b011010111100;
   22328: result <= 12'b011010111100;
   22329: result <= 12'b011010111100;
   22330: result <= 12'b011010111100;
   22331: result <= 12'b011010111100;
   22332: result <= 12'b011010111011;
   22333: result <= 12'b011010111011;
   22334: result <= 12'b011010111011;
   22335: result <= 12'b011010111011;
   22336: result <= 12'b011010111011;
   22337: result <= 12'b011010111011;
   22338: result <= 12'b011010111011;
   22339: result <= 12'b011010111011;
   22340: result <= 12'b011010111011;
   22341: result <= 12'b011010111010;
   22342: result <= 12'b011010111010;
   22343: result <= 12'b011010111010;
   22344: result <= 12'b011010111010;
   22345: result <= 12'b011010111010;
   22346: result <= 12'b011010111010;
   22347: result <= 12'b011010111010;
   22348: result <= 12'b011010111010;
   22349: result <= 12'b011010111010;
   22350: result <= 12'b011010111010;
   22351: result <= 12'b011010111001;
   22352: result <= 12'b011010111001;
   22353: result <= 12'b011010111001;
   22354: result <= 12'b011010111001;
   22355: result <= 12'b011010111001;
   22356: result <= 12'b011010111001;
   22357: result <= 12'b011010111001;
   22358: result <= 12'b011010111001;
   22359: result <= 12'b011010111001;
   22360: result <= 12'b011010111000;
   22361: result <= 12'b011010111000;
   22362: result <= 12'b011010111000;
   22363: result <= 12'b011010111000;
   22364: result <= 12'b011010111000;
   22365: result <= 12'b011010111000;
   22366: result <= 12'b011010111000;
   22367: result <= 12'b011010111000;
   22368: result <= 12'b011010111000;
   22369: result <= 12'b011010110111;
   22370: result <= 12'b011010110111;
   22371: result <= 12'b011010110111;
   22372: result <= 12'b011010110111;
   22373: result <= 12'b011010110111;
   22374: result <= 12'b011010110111;
   22375: result <= 12'b011010110111;
   22376: result <= 12'b011010110111;
   22377: result <= 12'b011010110111;
   22378: result <= 12'b011010110111;
   22379: result <= 12'b011010110110;
   22380: result <= 12'b011010110110;
   22381: result <= 12'b011010110110;
   22382: result <= 12'b011010110110;
   22383: result <= 12'b011010110110;
   22384: result <= 12'b011010110110;
   22385: result <= 12'b011010110110;
   22386: result <= 12'b011010110110;
   22387: result <= 12'b011010110110;
   22388: result <= 12'b011010110101;
   22389: result <= 12'b011010110101;
   22390: result <= 12'b011010110101;
   22391: result <= 12'b011010110101;
   22392: result <= 12'b011010110101;
   22393: result <= 12'b011010110101;
   22394: result <= 12'b011010110101;
   22395: result <= 12'b011010110101;
   22396: result <= 12'b011010110101;
   22397: result <= 12'b011010110101;
   22398: result <= 12'b011010110100;
   22399: result <= 12'b011010110100;
   22400: result <= 12'b011010110100;
   22401: result <= 12'b011010110100;
   22402: result <= 12'b011010110100;
   22403: result <= 12'b011010110100;
   22404: result <= 12'b011010110100;
   22405: result <= 12'b011010110100;
   22406: result <= 12'b011010110100;
   22407: result <= 12'b011010110011;
   22408: result <= 12'b011010110011;
   22409: result <= 12'b011010110011;
   22410: result <= 12'b011010110011;
   22411: result <= 12'b011010110011;
   22412: result <= 12'b011010110011;
   22413: result <= 12'b011010110011;
   22414: result <= 12'b011010110011;
   22415: result <= 12'b011010110011;
   22416: result <= 12'b011010110010;
   22417: result <= 12'b011010110010;
   22418: result <= 12'b011010110010;
   22419: result <= 12'b011010110010;
   22420: result <= 12'b011010110010;
   22421: result <= 12'b011010110010;
   22422: result <= 12'b011010110010;
   22423: result <= 12'b011010110010;
   22424: result <= 12'b011010110010;
   22425: result <= 12'b011010110010;
   22426: result <= 12'b011010110001;
   22427: result <= 12'b011010110001;
   22428: result <= 12'b011010110001;
   22429: result <= 12'b011010110001;
   22430: result <= 12'b011010110001;
   22431: result <= 12'b011010110001;
   22432: result <= 12'b011010110001;
   22433: result <= 12'b011010110001;
   22434: result <= 12'b011010110001;
   22435: result <= 12'b011010110000;
   22436: result <= 12'b011010110000;
   22437: result <= 12'b011010110000;
   22438: result <= 12'b011010110000;
   22439: result <= 12'b011010110000;
   22440: result <= 12'b011010110000;
   22441: result <= 12'b011010110000;
   22442: result <= 12'b011010110000;
   22443: result <= 12'b011010110000;
   22444: result <= 12'b011010101111;
   22445: result <= 12'b011010101111;
   22446: result <= 12'b011010101111;
   22447: result <= 12'b011010101111;
   22448: result <= 12'b011010101111;
   22449: result <= 12'b011010101111;
   22450: result <= 12'b011010101111;
   22451: result <= 12'b011010101111;
   22452: result <= 12'b011010101111;
   22453: result <= 12'b011010101110;
   22454: result <= 12'b011010101110;
   22455: result <= 12'b011010101110;
   22456: result <= 12'b011010101110;
   22457: result <= 12'b011010101110;
   22458: result <= 12'b011010101110;
   22459: result <= 12'b011010101110;
   22460: result <= 12'b011010101110;
   22461: result <= 12'b011010101110;
   22462: result <= 12'b011010101110;
   22463: result <= 12'b011010101101;
   22464: result <= 12'b011010101101;
   22465: result <= 12'b011010101101;
   22466: result <= 12'b011010101101;
   22467: result <= 12'b011010101101;
   22468: result <= 12'b011010101101;
   22469: result <= 12'b011010101101;
   22470: result <= 12'b011010101101;
   22471: result <= 12'b011010101101;
   22472: result <= 12'b011010101100;
   22473: result <= 12'b011010101100;
   22474: result <= 12'b011010101100;
   22475: result <= 12'b011010101100;
   22476: result <= 12'b011010101100;
   22477: result <= 12'b011010101100;
   22478: result <= 12'b011010101100;
   22479: result <= 12'b011010101100;
   22480: result <= 12'b011010101100;
   22481: result <= 12'b011010101011;
   22482: result <= 12'b011010101011;
   22483: result <= 12'b011010101011;
   22484: result <= 12'b011010101011;
   22485: result <= 12'b011010101011;
   22486: result <= 12'b011010101011;
   22487: result <= 12'b011010101011;
   22488: result <= 12'b011010101011;
   22489: result <= 12'b011010101011;
   22490: result <= 12'b011010101010;
   22491: result <= 12'b011010101010;
   22492: result <= 12'b011010101010;
   22493: result <= 12'b011010101010;
   22494: result <= 12'b011010101010;
   22495: result <= 12'b011010101010;
   22496: result <= 12'b011010101010;
   22497: result <= 12'b011010101010;
   22498: result <= 12'b011010101010;
   22499: result <= 12'b011010101010;
   22500: result <= 12'b011010101001;
   22501: result <= 12'b011010101001;
   22502: result <= 12'b011010101001;
   22503: result <= 12'b011010101001;
   22504: result <= 12'b011010101001;
   22505: result <= 12'b011010101001;
   22506: result <= 12'b011010101001;
   22507: result <= 12'b011010101001;
   22508: result <= 12'b011010101001;
   22509: result <= 12'b011010101000;
   22510: result <= 12'b011010101000;
   22511: result <= 12'b011010101000;
   22512: result <= 12'b011010101000;
   22513: result <= 12'b011010101000;
   22514: result <= 12'b011010101000;
   22515: result <= 12'b011010101000;
   22516: result <= 12'b011010101000;
   22517: result <= 12'b011010101000;
   22518: result <= 12'b011010100111;
   22519: result <= 12'b011010100111;
   22520: result <= 12'b011010100111;
   22521: result <= 12'b011010100111;
   22522: result <= 12'b011010100111;
   22523: result <= 12'b011010100111;
   22524: result <= 12'b011010100111;
   22525: result <= 12'b011010100111;
   22526: result <= 12'b011010100111;
   22527: result <= 12'b011010100110;
   22528: result <= 12'b011010100110;
   22529: result <= 12'b011010100110;
   22530: result <= 12'b011010100110;
   22531: result <= 12'b011010100110;
   22532: result <= 12'b011010100110;
   22533: result <= 12'b011010100110;
   22534: result <= 12'b011010100110;
   22535: result <= 12'b011010100110;
   22536: result <= 12'b011010100101;
   22537: result <= 12'b011010100101;
   22538: result <= 12'b011010100101;
   22539: result <= 12'b011010100101;
   22540: result <= 12'b011010100101;
   22541: result <= 12'b011010100101;
   22542: result <= 12'b011010100101;
   22543: result <= 12'b011010100101;
   22544: result <= 12'b011010100101;
   22545: result <= 12'b011010100100;
   22546: result <= 12'b011010100100;
   22547: result <= 12'b011010100100;
   22548: result <= 12'b011010100100;
   22549: result <= 12'b011010100100;
   22550: result <= 12'b011010100100;
   22551: result <= 12'b011010100100;
   22552: result <= 12'b011010100100;
   22553: result <= 12'b011010100100;
   22554: result <= 12'b011010100100;
   22555: result <= 12'b011010100011;
   22556: result <= 12'b011010100011;
   22557: result <= 12'b011010100011;
   22558: result <= 12'b011010100011;
   22559: result <= 12'b011010100011;
   22560: result <= 12'b011010100011;
   22561: result <= 12'b011010100011;
   22562: result <= 12'b011010100011;
   22563: result <= 12'b011010100011;
   22564: result <= 12'b011010100010;
   22565: result <= 12'b011010100010;
   22566: result <= 12'b011010100010;
   22567: result <= 12'b011010100010;
   22568: result <= 12'b011010100010;
   22569: result <= 12'b011010100010;
   22570: result <= 12'b011010100010;
   22571: result <= 12'b011010100010;
   22572: result <= 12'b011010100010;
   22573: result <= 12'b011010100001;
   22574: result <= 12'b011010100001;
   22575: result <= 12'b011010100001;
   22576: result <= 12'b011010100001;
   22577: result <= 12'b011010100001;
   22578: result <= 12'b011010100001;
   22579: result <= 12'b011010100001;
   22580: result <= 12'b011010100001;
   22581: result <= 12'b011010100001;
   22582: result <= 12'b011010100000;
   22583: result <= 12'b011010100000;
   22584: result <= 12'b011010100000;
   22585: result <= 12'b011010100000;
   22586: result <= 12'b011010100000;
   22587: result <= 12'b011010100000;
   22588: result <= 12'b011010100000;
   22589: result <= 12'b011010100000;
   22590: result <= 12'b011010100000;
   22591: result <= 12'b011010011111;
   22592: result <= 12'b011010011111;
   22593: result <= 12'b011010011111;
   22594: result <= 12'b011010011111;
   22595: result <= 12'b011010011111;
   22596: result <= 12'b011010011111;
   22597: result <= 12'b011010011111;
   22598: result <= 12'b011010011111;
   22599: result <= 12'b011010011111;
   22600: result <= 12'b011010011110;
   22601: result <= 12'b011010011110;
   22602: result <= 12'b011010011110;
   22603: result <= 12'b011010011110;
   22604: result <= 12'b011010011110;
   22605: result <= 12'b011010011110;
   22606: result <= 12'b011010011110;
   22607: result <= 12'b011010011110;
   22608: result <= 12'b011010011110;
   22609: result <= 12'b011010011101;
   22610: result <= 12'b011010011101;
   22611: result <= 12'b011010011101;
   22612: result <= 12'b011010011101;
   22613: result <= 12'b011010011101;
   22614: result <= 12'b011010011101;
   22615: result <= 12'b011010011101;
   22616: result <= 12'b011010011101;
   22617: result <= 12'b011010011101;
   22618: result <= 12'b011010011100;
   22619: result <= 12'b011010011100;
   22620: result <= 12'b011010011100;
   22621: result <= 12'b011010011100;
   22622: result <= 12'b011010011100;
   22623: result <= 12'b011010011100;
   22624: result <= 12'b011010011100;
   22625: result <= 12'b011010011100;
   22626: result <= 12'b011010011100;
   22627: result <= 12'b011010011011;
   22628: result <= 12'b011010011011;
   22629: result <= 12'b011010011011;
   22630: result <= 12'b011010011011;
   22631: result <= 12'b011010011011;
   22632: result <= 12'b011010011011;
   22633: result <= 12'b011010011011;
   22634: result <= 12'b011010011011;
   22635: result <= 12'b011010011011;
   22636: result <= 12'b011010011010;
   22637: result <= 12'b011010011010;
   22638: result <= 12'b011010011010;
   22639: result <= 12'b011010011010;
   22640: result <= 12'b011010011010;
   22641: result <= 12'b011010011010;
   22642: result <= 12'b011010011010;
   22643: result <= 12'b011010011010;
   22644: result <= 12'b011010011010;
   22645: result <= 12'b011010011001;
   22646: result <= 12'b011010011001;
   22647: result <= 12'b011010011001;
   22648: result <= 12'b011010011001;
   22649: result <= 12'b011010011001;
   22650: result <= 12'b011010011001;
   22651: result <= 12'b011010011001;
   22652: result <= 12'b011010011001;
   22653: result <= 12'b011010011001;
   22654: result <= 12'b011010011000;
   22655: result <= 12'b011010011000;
   22656: result <= 12'b011010011000;
   22657: result <= 12'b011010011000;
   22658: result <= 12'b011010011000;
   22659: result <= 12'b011010011000;
   22660: result <= 12'b011010011000;
   22661: result <= 12'b011010011000;
   22662: result <= 12'b011010011000;
   22663: result <= 12'b011010010111;
   22664: result <= 12'b011010010111;
   22665: result <= 12'b011010010111;
   22666: result <= 12'b011010010111;
   22667: result <= 12'b011010010111;
   22668: result <= 12'b011010010111;
   22669: result <= 12'b011010010111;
   22670: result <= 12'b011010010111;
   22671: result <= 12'b011010010111;
   22672: result <= 12'b011010010110;
   22673: result <= 12'b011010010110;
   22674: result <= 12'b011010010110;
   22675: result <= 12'b011010010110;
   22676: result <= 12'b011010010110;
   22677: result <= 12'b011010010110;
   22678: result <= 12'b011010010110;
   22679: result <= 12'b011010010110;
   22680: result <= 12'b011010010110;
   22681: result <= 12'b011010010101;
   22682: result <= 12'b011010010101;
   22683: result <= 12'b011010010101;
   22684: result <= 12'b011010010101;
   22685: result <= 12'b011010010101;
   22686: result <= 12'b011010010101;
   22687: result <= 12'b011010010101;
   22688: result <= 12'b011010010101;
   22689: result <= 12'b011010010101;
   22690: result <= 12'b011010010100;
   22691: result <= 12'b011010010100;
   22692: result <= 12'b011010010100;
   22693: result <= 12'b011010010100;
   22694: result <= 12'b011010010100;
   22695: result <= 12'b011010010100;
   22696: result <= 12'b011010010100;
   22697: result <= 12'b011010010100;
   22698: result <= 12'b011010010100;
   22699: result <= 12'b011010010011;
   22700: result <= 12'b011010010011;
   22701: result <= 12'b011010010011;
   22702: result <= 12'b011010010011;
   22703: result <= 12'b011010010011;
   22704: result <= 12'b011010010011;
   22705: result <= 12'b011010010011;
   22706: result <= 12'b011010010011;
   22707: result <= 12'b011010010011;
   22708: result <= 12'b011010010010;
   22709: result <= 12'b011010010010;
   22710: result <= 12'b011010010010;
   22711: result <= 12'b011010010010;
   22712: result <= 12'b011010010010;
   22713: result <= 12'b011010010010;
   22714: result <= 12'b011010010010;
   22715: result <= 12'b011010010010;
   22716: result <= 12'b011010010010;
   22717: result <= 12'b011010010001;
   22718: result <= 12'b011010010001;
   22719: result <= 12'b011010010001;
   22720: result <= 12'b011010010001;
   22721: result <= 12'b011010010001;
   22722: result <= 12'b011010010001;
   22723: result <= 12'b011010010001;
   22724: result <= 12'b011010010001;
   22725: result <= 12'b011010010001;
   22726: result <= 12'b011010010000;
   22727: result <= 12'b011010010000;
   22728: result <= 12'b011010010000;
   22729: result <= 12'b011010010000;
   22730: result <= 12'b011010010000;
   22731: result <= 12'b011010010000;
   22732: result <= 12'b011010010000;
   22733: result <= 12'b011010010000;
   22734: result <= 12'b011010010000;
   22735: result <= 12'b011010001111;
   22736: result <= 12'b011010001111;
   22737: result <= 12'b011010001111;
   22738: result <= 12'b011010001111;
   22739: result <= 12'b011010001111;
   22740: result <= 12'b011010001111;
   22741: result <= 12'b011010001111;
   22742: result <= 12'b011010001111;
   22743: result <= 12'b011010001111;
   22744: result <= 12'b011010001110;
   22745: result <= 12'b011010001110;
   22746: result <= 12'b011010001110;
   22747: result <= 12'b011010001110;
   22748: result <= 12'b011010001110;
   22749: result <= 12'b011010001110;
   22750: result <= 12'b011010001110;
   22751: result <= 12'b011010001110;
   22752: result <= 12'b011010001110;
   22753: result <= 12'b011010001101;
   22754: result <= 12'b011010001101;
   22755: result <= 12'b011010001101;
   22756: result <= 12'b011010001101;
   22757: result <= 12'b011010001101;
   22758: result <= 12'b011010001101;
   22759: result <= 12'b011010001101;
   22760: result <= 12'b011010001101;
   22761: result <= 12'b011010001101;
   22762: result <= 12'b011010001100;
   22763: result <= 12'b011010001100;
   22764: result <= 12'b011010001100;
   22765: result <= 12'b011010001100;
   22766: result <= 12'b011010001100;
   22767: result <= 12'b011010001100;
   22768: result <= 12'b011010001100;
   22769: result <= 12'b011010001100;
   22770: result <= 12'b011010001011;
   22771: result <= 12'b011010001011;
   22772: result <= 12'b011010001011;
   22773: result <= 12'b011010001011;
   22774: result <= 12'b011010001011;
   22775: result <= 12'b011010001011;
   22776: result <= 12'b011010001011;
   22777: result <= 12'b011010001011;
   22778: result <= 12'b011010001011;
   22779: result <= 12'b011010001010;
   22780: result <= 12'b011010001010;
   22781: result <= 12'b011010001010;
   22782: result <= 12'b011010001010;
   22783: result <= 12'b011010001010;
   22784: result <= 12'b011010001010;
   22785: result <= 12'b011010001010;
   22786: result <= 12'b011010001010;
   22787: result <= 12'b011010001010;
   22788: result <= 12'b011010001001;
   22789: result <= 12'b011010001001;
   22790: result <= 12'b011010001001;
   22791: result <= 12'b011010001001;
   22792: result <= 12'b011010001001;
   22793: result <= 12'b011010001001;
   22794: result <= 12'b011010001001;
   22795: result <= 12'b011010001001;
   22796: result <= 12'b011010001001;
   22797: result <= 12'b011010001000;
   22798: result <= 12'b011010001000;
   22799: result <= 12'b011010001000;
   22800: result <= 12'b011010001000;
   22801: result <= 12'b011010001000;
   22802: result <= 12'b011010001000;
   22803: result <= 12'b011010001000;
   22804: result <= 12'b011010001000;
   22805: result <= 12'b011010001000;
   22806: result <= 12'b011010000111;
   22807: result <= 12'b011010000111;
   22808: result <= 12'b011010000111;
   22809: result <= 12'b011010000111;
   22810: result <= 12'b011010000111;
   22811: result <= 12'b011010000111;
   22812: result <= 12'b011010000111;
   22813: result <= 12'b011010000111;
   22814: result <= 12'b011010000111;
   22815: result <= 12'b011010000110;
   22816: result <= 12'b011010000110;
   22817: result <= 12'b011010000110;
   22818: result <= 12'b011010000110;
   22819: result <= 12'b011010000110;
   22820: result <= 12'b011010000110;
   22821: result <= 12'b011010000110;
   22822: result <= 12'b011010000110;
   22823: result <= 12'b011010000101;
   22824: result <= 12'b011010000101;
   22825: result <= 12'b011010000101;
   22826: result <= 12'b011010000101;
   22827: result <= 12'b011010000101;
   22828: result <= 12'b011010000101;
   22829: result <= 12'b011010000101;
   22830: result <= 12'b011010000101;
   22831: result <= 12'b011010000101;
   22832: result <= 12'b011010000100;
   22833: result <= 12'b011010000100;
   22834: result <= 12'b011010000100;
   22835: result <= 12'b011010000100;
   22836: result <= 12'b011010000100;
   22837: result <= 12'b011010000100;
   22838: result <= 12'b011010000100;
   22839: result <= 12'b011010000100;
   22840: result <= 12'b011010000100;
   22841: result <= 12'b011010000011;
   22842: result <= 12'b011010000011;
   22843: result <= 12'b011010000011;
   22844: result <= 12'b011010000011;
   22845: result <= 12'b011010000011;
   22846: result <= 12'b011010000011;
   22847: result <= 12'b011010000011;
   22848: result <= 12'b011010000011;
   22849: result <= 12'b011010000011;
   22850: result <= 12'b011010000010;
   22851: result <= 12'b011010000010;
   22852: result <= 12'b011010000010;
   22853: result <= 12'b011010000010;
   22854: result <= 12'b011010000010;
   22855: result <= 12'b011010000010;
   22856: result <= 12'b011010000010;
   22857: result <= 12'b011010000010;
   22858: result <= 12'b011010000010;
   22859: result <= 12'b011010000001;
   22860: result <= 12'b011010000001;
   22861: result <= 12'b011010000001;
   22862: result <= 12'b011010000001;
   22863: result <= 12'b011010000001;
   22864: result <= 12'b011010000001;
   22865: result <= 12'b011010000001;
   22866: result <= 12'b011010000001;
   22867: result <= 12'b011010000000;
   22868: result <= 12'b011010000000;
   22869: result <= 12'b011010000000;
   22870: result <= 12'b011010000000;
   22871: result <= 12'b011010000000;
   22872: result <= 12'b011010000000;
   22873: result <= 12'b011010000000;
   22874: result <= 12'b011010000000;
   22875: result <= 12'b011010000000;
   22876: result <= 12'b011001111111;
   22877: result <= 12'b011001111111;
   22878: result <= 12'b011001111111;
   22879: result <= 12'b011001111111;
   22880: result <= 12'b011001111111;
   22881: result <= 12'b011001111111;
   22882: result <= 12'b011001111111;
   22883: result <= 12'b011001111111;
   22884: result <= 12'b011001111111;
   22885: result <= 12'b011001111110;
   22886: result <= 12'b011001111110;
   22887: result <= 12'b011001111110;
   22888: result <= 12'b011001111110;
   22889: result <= 12'b011001111110;
   22890: result <= 12'b011001111110;
   22891: result <= 12'b011001111110;
   22892: result <= 12'b011001111110;
   22893: result <= 12'b011001111101;
   22894: result <= 12'b011001111101;
   22895: result <= 12'b011001111101;
   22896: result <= 12'b011001111101;
   22897: result <= 12'b011001111101;
   22898: result <= 12'b011001111101;
   22899: result <= 12'b011001111101;
   22900: result <= 12'b011001111101;
   22901: result <= 12'b011001111101;
   22902: result <= 12'b011001111100;
   22903: result <= 12'b011001111100;
   22904: result <= 12'b011001111100;
   22905: result <= 12'b011001111100;
   22906: result <= 12'b011001111100;
   22907: result <= 12'b011001111100;
   22908: result <= 12'b011001111100;
   22909: result <= 12'b011001111100;
   22910: result <= 12'b011001111100;
   22911: result <= 12'b011001111011;
   22912: result <= 12'b011001111011;
   22913: result <= 12'b011001111011;
   22914: result <= 12'b011001111011;
   22915: result <= 12'b011001111011;
   22916: result <= 12'b011001111011;
   22917: result <= 12'b011001111011;
   22918: result <= 12'b011001111011;
   22919: result <= 12'b011001111011;
   22920: result <= 12'b011001111010;
   22921: result <= 12'b011001111010;
   22922: result <= 12'b011001111010;
   22923: result <= 12'b011001111010;
   22924: result <= 12'b011001111010;
   22925: result <= 12'b011001111010;
   22926: result <= 12'b011001111010;
   22927: result <= 12'b011001111010;
   22928: result <= 12'b011001111001;
   22929: result <= 12'b011001111001;
   22930: result <= 12'b011001111001;
   22931: result <= 12'b011001111001;
   22932: result <= 12'b011001111001;
   22933: result <= 12'b011001111001;
   22934: result <= 12'b011001111001;
   22935: result <= 12'b011001111001;
   22936: result <= 12'b011001111001;
   22937: result <= 12'b011001111000;
   22938: result <= 12'b011001111000;
   22939: result <= 12'b011001111000;
   22940: result <= 12'b011001111000;
   22941: result <= 12'b011001111000;
   22942: result <= 12'b011001111000;
   22943: result <= 12'b011001111000;
   22944: result <= 12'b011001111000;
   22945: result <= 12'b011001111000;
   22946: result <= 12'b011001110111;
   22947: result <= 12'b011001110111;
   22948: result <= 12'b011001110111;
   22949: result <= 12'b011001110111;
   22950: result <= 12'b011001110111;
   22951: result <= 12'b011001110111;
   22952: result <= 12'b011001110111;
   22953: result <= 12'b011001110111;
   22954: result <= 12'b011001110110;
   22955: result <= 12'b011001110110;
   22956: result <= 12'b011001110110;
   22957: result <= 12'b011001110110;
   22958: result <= 12'b011001110110;
   22959: result <= 12'b011001110110;
   22960: result <= 12'b011001110110;
   22961: result <= 12'b011001110110;
   22962: result <= 12'b011001110110;
   22963: result <= 12'b011001110101;
   22964: result <= 12'b011001110101;
   22965: result <= 12'b011001110101;
   22966: result <= 12'b011001110101;
   22967: result <= 12'b011001110101;
   22968: result <= 12'b011001110101;
   22969: result <= 12'b011001110101;
   22970: result <= 12'b011001110101;
   22971: result <= 12'b011001110101;
   22972: result <= 12'b011001110100;
   22973: result <= 12'b011001110100;
   22974: result <= 12'b011001110100;
   22975: result <= 12'b011001110100;
   22976: result <= 12'b011001110100;
   22977: result <= 12'b011001110100;
   22978: result <= 12'b011001110100;
   22979: result <= 12'b011001110100;
   22980: result <= 12'b011001110011;
   22981: result <= 12'b011001110011;
   22982: result <= 12'b011001110011;
   22983: result <= 12'b011001110011;
   22984: result <= 12'b011001110011;
   22985: result <= 12'b011001110011;
   22986: result <= 12'b011001110011;
   22987: result <= 12'b011001110011;
   22988: result <= 12'b011001110011;
   22989: result <= 12'b011001110010;
   22990: result <= 12'b011001110010;
   22991: result <= 12'b011001110010;
   22992: result <= 12'b011001110010;
   22993: result <= 12'b011001110010;
   22994: result <= 12'b011001110010;
   22995: result <= 12'b011001110010;
   22996: result <= 12'b011001110010;
   22997: result <= 12'b011001110001;
   22998: result <= 12'b011001110001;
   22999: result <= 12'b011001110001;
   23000: result <= 12'b011001110001;
   23001: result <= 12'b011001110001;
   23002: result <= 12'b011001110001;
   23003: result <= 12'b011001110001;
   23004: result <= 12'b011001110001;
   23005: result <= 12'b011001110001;
   23006: result <= 12'b011001110000;
   23007: result <= 12'b011001110000;
   23008: result <= 12'b011001110000;
   23009: result <= 12'b011001110000;
   23010: result <= 12'b011001110000;
   23011: result <= 12'b011001110000;
   23012: result <= 12'b011001110000;
   23013: result <= 12'b011001110000;
   23014: result <= 12'b011001110000;
   23015: result <= 12'b011001101111;
   23016: result <= 12'b011001101111;
   23017: result <= 12'b011001101111;
   23018: result <= 12'b011001101111;
   23019: result <= 12'b011001101111;
   23020: result <= 12'b011001101111;
   23021: result <= 12'b011001101111;
   23022: result <= 12'b011001101111;
   23023: result <= 12'b011001101110;
   23024: result <= 12'b011001101110;
   23025: result <= 12'b011001101110;
   23026: result <= 12'b011001101110;
   23027: result <= 12'b011001101110;
   23028: result <= 12'b011001101110;
   23029: result <= 12'b011001101110;
   23030: result <= 12'b011001101110;
   23031: result <= 12'b011001101110;
   23032: result <= 12'b011001101101;
   23033: result <= 12'b011001101101;
   23034: result <= 12'b011001101101;
   23035: result <= 12'b011001101101;
   23036: result <= 12'b011001101101;
   23037: result <= 12'b011001101101;
   23038: result <= 12'b011001101101;
   23039: result <= 12'b011001101101;
   23040: result <= 12'b011001101100;
   23041: result <= 12'b011001101100;
   23042: result <= 12'b011001101100;
   23043: result <= 12'b011001101100;
   23044: result <= 12'b011001101100;
   23045: result <= 12'b011001101100;
   23046: result <= 12'b011001101100;
   23047: result <= 12'b011001101100;
   23048: result <= 12'b011001101100;
   23049: result <= 12'b011001101011;
   23050: result <= 12'b011001101011;
   23051: result <= 12'b011001101011;
   23052: result <= 12'b011001101011;
   23053: result <= 12'b011001101011;
   23054: result <= 12'b011001101011;
   23055: result <= 12'b011001101011;
   23056: result <= 12'b011001101011;
   23057: result <= 12'b011001101010;
   23058: result <= 12'b011001101010;
   23059: result <= 12'b011001101010;
   23060: result <= 12'b011001101010;
   23061: result <= 12'b011001101010;
   23062: result <= 12'b011001101010;
   23063: result <= 12'b011001101010;
   23064: result <= 12'b011001101010;
   23065: result <= 12'b011001101010;
   23066: result <= 12'b011001101001;
   23067: result <= 12'b011001101001;
   23068: result <= 12'b011001101001;
   23069: result <= 12'b011001101001;
   23070: result <= 12'b011001101001;
   23071: result <= 12'b011001101001;
   23072: result <= 12'b011001101001;
   23073: result <= 12'b011001101001;
   23074: result <= 12'b011001101000;
   23075: result <= 12'b011001101000;
   23076: result <= 12'b011001101000;
   23077: result <= 12'b011001101000;
   23078: result <= 12'b011001101000;
   23079: result <= 12'b011001101000;
   23080: result <= 12'b011001101000;
   23081: result <= 12'b011001101000;
   23082: result <= 12'b011001101000;
   23083: result <= 12'b011001100111;
   23084: result <= 12'b011001100111;
   23085: result <= 12'b011001100111;
   23086: result <= 12'b011001100111;
   23087: result <= 12'b011001100111;
   23088: result <= 12'b011001100111;
   23089: result <= 12'b011001100111;
   23090: result <= 12'b011001100111;
   23091: result <= 12'b011001100110;
   23092: result <= 12'b011001100110;
   23093: result <= 12'b011001100110;
   23094: result <= 12'b011001100110;
   23095: result <= 12'b011001100110;
   23096: result <= 12'b011001100110;
   23097: result <= 12'b011001100110;
   23098: result <= 12'b011001100110;
   23099: result <= 12'b011001100110;
   23100: result <= 12'b011001100101;
   23101: result <= 12'b011001100101;
   23102: result <= 12'b011001100101;
   23103: result <= 12'b011001100101;
   23104: result <= 12'b011001100101;
   23105: result <= 12'b011001100101;
   23106: result <= 12'b011001100101;
   23107: result <= 12'b011001100101;
   23108: result <= 12'b011001100100;
   23109: result <= 12'b011001100100;
   23110: result <= 12'b011001100100;
   23111: result <= 12'b011001100100;
   23112: result <= 12'b011001100100;
   23113: result <= 12'b011001100100;
   23114: result <= 12'b011001100100;
   23115: result <= 12'b011001100100;
   23116: result <= 12'b011001100100;
   23117: result <= 12'b011001100011;
   23118: result <= 12'b011001100011;
   23119: result <= 12'b011001100011;
   23120: result <= 12'b011001100011;
   23121: result <= 12'b011001100011;
   23122: result <= 12'b011001100011;
   23123: result <= 12'b011001100011;
   23124: result <= 12'b011001100011;
   23125: result <= 12'b011001100010;
   23126: result <= 12'b011001100010;
   23127: result <= 12'b011001100010;
   23128: result <= 12'b011001100010;
   23129: result <= 12'b011001100010;
   23130: result <= 12'b011001100010;
   23131: result <= 12'b011001100010;
   23132: result <= 12'b011001100010;
   23133: result <= 12'b011001100010;
   23134: result <= 12'b011001100001;
   23135: result <= 12'b011001100001;
   23136: result <= 12'b011001100001;
   23137: result <= 12'b011001100001;
   23138: result <= 12'b011001100001;
   23139: result <= 12'b011001100001;
   23140: result <= 12'b011001100001;
   23141: result <= 12'b011001100001;
   23142: result <= 12'b011001100000;
   23143: result <= 12'b011001100000;
   23144: result <= 12'b011001100000;
   23145: result <= 12'b011001100000;
   23146: result <= 12'b011001100000;
   23147: result <= 12'b011001100000;
   23148: result <= 12'b011001100000;
   23149: result <= 12'b011001100000;
   23150: result <= 12'b011001100000;
   23151: result <= 12'b011001011111;
   23152: result <= 12'b011001011111;
   23153: result <= 12'b011001011111;
   23154: result <= 12'b011001011111;
   23155: result <= 12'b011001011111;
   23156: result <= 12'b011001011111;
   23157: result <= 12'b011001011111;
   23158: result <= 12'b011001011111;
   23159: result <= 12'b011001011110;
   23160: result <= 12'b011001011110;
   23161: result <= 12'b011001011110;
   23162: result <= 12'b011001011110;
   23163: result <= 12'b011001011110;
   23164: result <= 12'b011001011110;
   23165: result <= 12'b011001011110;
   23166: result <= 12'b011001011110;
   23167: result <= 12'b011001011101;
   23168: result <= 12'b011001011101;
   23169: result <= 12'b011001011101;
   23170: result <= 12'b011001011101;
   23171: result <= 12'b011001011101;
   23172: result <= 12'b011001011101;
   23173: result <= 12'b011001011101;
   23174: result <= 12'b011001011101;
   23175: result <= 12'b011001011101;
   23176: result <= 12'b011001011100;
   23177: result <= 12'b011001011100;
   23178: result <= 12'b011001011100;
   23179: result <= 12'b011001011100;
   23180: result <= 12'b011001011100;
   23181: result <= 12'b011001011100;
   23182: result <= 12'b011001011100;
   23183: result <= 12'b011001011100;
   23184: result <= 12'b011001011011;
   23185: result <= 12'b011001011011;
   23186: result <= 12'b011001011011;
   23187: result <= 12'b011001011011;
   23188: result <= 12'b011001011011;
   23189: result <= 12'b011001011011;
   23190: result <= 12'b011001011011;
   23191: result <= 12'b011001011011;
   23192: result <= 12'b011001011011;
   23193: result <= 12'b011001011010;
   23194: result <= 12'b011001011010;
   23195: result <= 12'b011001011010;
   23196: result <= 12'b011001011010;
   23197: result <= 12'b011001011010;
   23198: result <= 12'b011001011010;
   23199: result <= 12'b011001011010;
   23200: result <= 12'b011001011010;
   23201: result <= 12'b011001011001;
   23202: result <= 12'b011001011001;
   23203: result <= 12'b011001011001;
   23204: result <= 12'b011001011001;
   23205: result <= 12'b011001011001;
   23206: result <= 12'b011001011001;
   23207: result <= 12'b011001011001;
   23208: result <= 12'b011001011001;
   23209: result <= 12'b011001011000;
   23210: result <= 12'b011001011000;
   23211: result <= 12'b011001011000;
   23212: result <= 12'b011001011000;
   23213: result <= 12'b011001011000;
   23214: result <= 12'b011001011000;
   23215: result <= 12'b011001011000;
   23216: result <= 12'b011001011000;
   23217: result <= 12'b011001011000;
   23218: result <= 12'b011001010111;
   23219: result <= 12'b011001010111;
   23220: result <= 12'b011001010111;
   23221: result <= 12'b011001010111;
   23222: result <= 12'b011001010111;
   23223: result <= 12'b011001010111;
   23224: result <= 12'b011001010111;
   23225: result <= 12'b011001010111;
   23226: result <= 12'b011001010110;
   23227: result <= 12'b011001010110;
   23228: result <= 12'b011001010110;
   23229: result <= 12'b011001010110;
   23230: result <= 12'b011001010110;
   23231: result <= 12'b011001010110;
   23232: result <= 12'b011001010110;
   23233: result <= 12'b011001010110;
   23234: result <= 12'b011001010101;
   23235: result <= 12'b011001010101;
   23236: result <= 12'b011001010101;
   23237: result <= 12'b011001010101;
   23238: result <= 12'b011001010101;
   23239: result <= 12'b011001010101;
   23240: result <= 12'b011001010101;
   23241: result <= 12'b011001010101;
   23242: result <= 12'b011001010101;
   23243: result <= 12'b011001010100;
   23244: result <= 12'b011001010100;
   23245: result <= 12'b011001010100;
   23246: result <= 12'b011001010100;
   23247: result <= 12'b011001010100;
   23248: result <= 12'b011001010100;
   23249: result <= 12'b011001010100;
   23250: result <= 12'b011001010100;
   23251: result <= 12'b011001010011;
   23252: result <= 12'b011001010011;
   23253: result <= 12'b011001010011;
   23254: result <= 12'b011001010011;
   23255: result <= 12'b011001010011;
   23256: result <= 12'b011001010011;
   23257: result <= 12'b011001010011;
   23258: result <= 12'b011001010011;
   23259: result <= 12'b011001010010;
   23260: result <= 12'b011001010010;
   23261: result <= 12'b011001010010;
   23262: result <= 12'b011001010010;
   23263: result <= 12'b011001010010;
   23264: result <= 12'b011001010010;
   23265: result <= 12'b011001010010;
   23266: result <= 12'b011001010010;
   23267: result <= 12'b011001010010;
   23268: result <= 12'b011001010001;
   23269: result <= 12'b011001010001;
   23270: result <= 12'b011001010001;
   23271: result <= 12'b011001010001;
   23272: result <= 12'b011001010001;
   23273: result <= 12'b011001010001;
   23274: result <= 12'b011001010001;
   23275: result <= 12'b011001010001;
   23276: result <= 12'b011001010000;
   23277: result <= 12'b011001010000;
   23278: result <= 12'b011001010000;
   23279: result <= 12'b011001010000;
   23280: result <= 12'b011001010000;
   23281: result <= 12'b011001010000;
   23282: result <= 12'b011001010000;
   23283: result <= 12'b011001010000;
   23284: result <= 12'b011001001111;
   23285: result <= 12'b011001001111;
   23286: result <= 12'b011001001111;
   23287: result <= 12'b011001001111;
   23288: result <= 12'b011001001111;
   23289: result <= 12'b011001001111;
   23290: result <= 12'b011001001111;
   23291: result <= 12'b011001001111;
   23292: result <= 12'b011001001111;
   23293: result <= 12'b011001001110;
   23294: result <= 12'b011001001110;
   23295: result <= 12'b011001001110;
   23296: result <= 12'b011001001110;
   23297: result <= 12'b011001001110;
   23298: result <= 12'b011001001110;
   23299: result <= 12'b011001001110;
   23300: result <= 12'b011001001110;
   23301: result <= 12'b011001001101;
   23302: result <= 12'b011001001101;
   23303: result <= 12'b011001001101;
   23304: result <= 12'b011001001101;
   23305: result <= 12'b011001001101;
   23306: result <= 12'b011001001101;
   23307: result <= 12'b011001001101;
   23308: result <= 12'b011001001101;
   23309: result <= 12'b011001001100;
   23310: result <= 12'b011001001100;
   23311: result <= 12'b011001001100;
   23312: result <= 12'b011001001100;
   23313: result <= 12'b011001001100;
   23314: result <= 12'b011001001100;
   23315: result <= 12'b011001001100;
   23316: result <= 12'b011001001100;
   23317: result <= 12'b011001001011;
   23318: result <= 12'b011001001011;
   23319: result <= 12'b011001001011;
   23320: result <= 12'b011001001011;
   23321: result <= 12'b011001001011;
   23322: result <= 12'b011001001011;
   23323: result <= 12'b011001001011;
   23324: result <= 12'b011001001011;
   23325: result <= 12'b011001001011;
   23326: result <= 12'b011001001010;
   23327: result <= 12'b011001001010;
   23328: result <= 12'b011001001010;
   23329: result <= 12'b011001001010;
   23330: result <= 12'b011001001010;
   23331: result <= 12'b011001001010;
   23332: result <= 12'b011001001010;
   23333: result <= 12'b011001001010;
   23334: result <= 12'b011001001001;
   23335: result <= 12'b011001001001;
   23336: result <= 12'b011001001001;
   23337: result <= 12'b011001001001;
   23338: result <= 12'b011001001001;
   23339: result <= 12'b011001001001;
   23340: result <= 12'b011001001001;
   23341: result <= 12'b011001001001;
   23342: result <= 12'b011001001000;
   23343: result <= 12'b011001001000;
   23344: result <= 12'b011001001000;
   23345: result <= 12'b011001001000;
   23346: result <= 12'b011001001000;
   23347: result <= 12'b011001001000;
   23348: result <= 12'b011001001000;
   23349: result <= 12'b011001001000;
   23350: result <= 12'b011001000111;
   23351: result <= 12'b011001000111;
   23352: result <= 12'b011001000111;
   23353: result <= 12'b011001000111;
   23354: result <= 12'b011001000111;
   23355: result <= 12'b011001000111;
   23356: result <= 12'b011001000111;
   23357: result <= 12'b011001000111;
   23358: result <= 12'b011001000111;
   23359: result <= 12'b011001000110;
   23360: result <= 12'b011001000110;
   23361: result <= 12'b011001000110;
   23362: result <= 12'b011001000110;
   23363: result <= 12'b011001000110;
   23364: result <= 12'b011001000110;
   23365: result <= 12'b011001000110;
   23366: result <= 12'b011001000110;
   23367: result <= 12'b011001000101;
   23368: result <= 12'b011001000101;
   23369: result <= 12'b011001000101;
   23370: result <= 12'b011001000101;
   23371: result <= 12'b011001000101;
   23372: result <= 12'b011001000101;
   23373: result <= 12'b011001000101;
   23374: result <= 12'b011001000101;
   23375: result <= 12'b011001000100;
   23376: result <= 12'b011001000100;
   23377: result <= 12'b011001000100;
   23378: result <= 12'b011001000100;
   23379: result <= 12'b011001000100;
   23380: result <= 12'b011001000100;
   23381: result <= 12'b011001000100;
   23382: result <= 12'b011001000100;
   23383: result <= 12'b011001000011;
   23384: result <= 12'b011001000011;
   23385: result <= 12'b011001000011;
   23386: result <= 12'b011001000011;
   23387: result <= 12'b011001000011;
   23388: result <= 12'b011001000011;
   23389: result <= 12'b011001000011;
   23390: result <= 12'b011001000011;
   23391: result <= 12'b011001000010;
   23392: result <= 12'b011001000010;
   23393: result <= 12'b011001000010;
   23394: result <= 12'b011001000010;
   23395: result <= 12'b011001000010;
   23396: result <= 12'b011001000010;
   23397: result <= 12'b011001000010;
   23398: result <= 12'b011001000010;
   23399: result <= 12'b011001000010;
   23400: result <= 12'b011001000001;
   23401: result <= 12'b011001000001;
   23402: result <= 12'b011001000001;
   23403: result <= 12'b011001000001;
   23404: result <= 12'b011001000001;
   23405: result <= 12'b011001000001;
   23406: result <= 12'b011001000001;
   23407: result <= 12'b011001000001;
   23408: result <= 12'b011001000000;
   23409: result <= 12'b011001000000;
   23410: result <= 12'b011001000000;
   23411: result <= 12'b011001000000;
   23412: result <= 12'b011001000000;
   23413: result <= 12'b011001000000;
   23414: result <= 12'b011001000000;
   23415: result <= 12'b011001000000;
   23416: result <= 12'b011000111111;
   23417: result <= 12'b011000111111;
   23418: result <= 12'b011000111111;
   23419: result <= 12'b011000111111;
   23420: result <= 12'b011000111111;
   23421: result <= 12'b011000111111;
   23422: result <= 12'b011000111111;
   23423: result <= 12'b011000111111;
   23424: result <= 12'b011000111110;
   23425: result <= 12'b011000111110;
   23426: result <= 12'b011000111110;
   23427: result <= 12'b011000111110;
   23428: result <= 12'b011000111110;
   23429: result <= 12'b011000111110;
   23430: result <= 12'b011000111110;
   23431: result <= 12'b011000111110;
   23432: result <= 12'b011000111101;
   23433: result <= 12'b011000111101;
   23434: result <= 12'b011000111101;
   23435: result <= 12'b011000111101;
   23436: result <= 12'b011000111101;
   23437: result <= 12'b011000111101;
   23438: result <= 12'b011000111101;
   23439: result <= 12'b011000111101;
   23440: result <= 12'b011000111100;
   23441: result <= 12'b011000111100;
   23442: result <= 12'b011000111100;
   23443: result <= 12'b011000111100;
   23444: result <= 12'b011000111100;
   23445: result <= 12'b011000111100;
   23446: result <= 12'b011000111100;
   23447: result <= 12'b011000111100;
   23448: result <= 12'b011000111100;
   23449: result <= 12'b011000111011;
   23450: result <= 12'b011000111011;
   23451: result <= 12'b011000111011;
   23452: result <= 12'b011000111011;
   23453: result <= 12'b011000111011;
   23454: result <= 12'b011000111011;
   23455: result <= 12'b011000111011;
   23456: result <= 12'b011000111011;
   23457: result <= 12'b011000111010;
   23458: result <= 12'b011000111010;
   23459: result <= 12'b011000111010;
   23460: result <= 12'b011000111010;
   23461: result <= 12'b011000111010;
   23462: result <= 12'b011000111010;
   23463: result <= 12'b011000111010;
   23464: result <= 12'b011000111010;
   23465: result <= 12'b011000111001;
   23466: result <= 12'b011000111001;
   23467: result <= 12'b011000111001;
   23468: result <= 12'b011000111001;
   23469: result <= 12'b011000111001;
   23470: result <= 12'b011000111001;
   23471: result <= 12'b011000111001;
   23472: result <= 12'b011000111001;
   23473: result <= 12'b011000111000;
   23474: result <= 12'b011000111000;
   23475: result <= 12'b011000111000;
   23476: result <= 12'b011000111000;
   23477: result <= 12'b011000111000;
   23478: result <= 12'b011000111000;
   23479: result <= 12'b011000111000;
   23480: result <= 12'b011000111000;
   23481: result <= 12'b011000110111;
   23482: result <= 12'b011000110111;
   23483: result <= 12'b011000110111;
   23484: result <= 12'b011000110111;
   23485: result <= 12'b011000110111;
   23486: result <= 12'b011000110111;
   23487: result <= 12'b011000110111;
   23488: result <= 12'b011000110111;
   23489: result <= 12'b011000110110;
   23490: result <= 12'b011000110110;
   23491: result <= 12'b011000110110;
   23492: result <= 12'b011000110110;
   23493: result <= 12'b011000110110;
   23494: result <= 12'b011000110110;
   23495: result <= 12'b011000110110;
   23496: result <= 12'b011000110110;
   23497: result <= 12'b011000110101;
   23498: result <= 12'b011000110101;
   23499: result <= 12'b011000110101;
   23500: result <= 12'b011000110101;
   23501: result <= 12'b011000110101;
   23502: result <= 12'b011000110101;
   23503: result <= 12'b011000110101;
   23504: result <= 12'b011000110101;
   23505: result <= 12'b011000110100;
   23506: result <= 12'b011000110100;
   23507: result <= 12'b011000110100;
   23508: result <= 12'b011000110100;
   23509: result <= 12'b011000110100;
   23510: result <= 12'b011000110100;
   23511: result <= 12'b011000110100;
   23512: result <= 12'b011000110100;
   23513: result <= 12'b011000110011;
   23514: result <= 12'b011000110011;
   23515: result <= 12'b011000110011;
   23516: result <= 12'b011000110011;
   23517: result <= 12'b011000110011;
   23518: result <= 12'b011000110011;
   23519: result <= 12'b011000110011;
   23520: result <= 12'b011000110011;
   23521: result <= 12'b011000110010;
   23522: result <= 12'b011000110010;
   23523: result <= 12'b011000110010;
   23524: result <= 12'b011000110010;
   23525: result <= 12'b011000110010;
   23526: result <= 12'b011000110010;
   23527: result <= 12'b011000110010;
   23528: result <= 12'b011000110010;
   23529: result <= 12'b011000110001;
   23530: result <= 12'b011000110001;
   23531: result <= 12'b011000110001;
   23532: result <= 12'b011000110001;
   23533: result <= 12'b011000110001;
   23534: result <= 12'b011000110001;
   23535: result <= 12'b011000110001;
   23536: result <= 12'b011000110001;
   23537: result <= 12'b011000110000;
   23538: result <= 12'b011000110000;
   23539: result <= 12'b011000110000;
   23540: result <= 12'b011000110000;
   23541: result <= 12'b011000110000;
   23542: result <= 12'b011000110000;
   23543: result <= 12'b011000110000;
   23544: result <= 12'b011000110000;
   23545: result <= 12'b011000101111;
   23546: result <= 12'b011000101111;
   23547: result <= 12'b011000101111;
   23548: result <= 12'b011000101111;
   23549: result <= 12'b011000101111;
   23550: result <= 12'b011000101111;
   23551: result <= 12'b011000101111;
   23552: result <= 12'b011000101111;
   23553: result <= 12'b011000101111;
   23554: result <= 12'b011000101110;
   23555: result <= 12'b011000101110;
   23556: result <= 12'b011000101110;
   23557: result <= 12'b011000101110;
   23558: result <= 12'b011000101110;
   23559: result <= 12'b011000101110;
   23560: result <= 12'b011000101110;
   23561: result <= 12'b011000101110;
   23562: result <= 12'b011000101101;
   23563: result <= 12'b011000101101;
   23564: result <= 12'b011000101101;
   23565: result <= 12'b011000101101;
   23566: result <= 12'b011000101101;
   23567: result <= 12'b011000101101;
   23568: result <= 12'b011000101101;
   23569: result <= 12'b011000101101;
   23570: result <= 12'b011000101100;
   23571: result <= 12'b011000101100;
   23572: result <= 12'b011000101100;
   23573: result <= 12'b011000101100;
   23574: result <= 12'b011000101100;
   23575: result <= 12'b011000101100;
   23576: result <= 12'b011000101100;
   23577: result <= 12'b011000101100;
   23578: result <= 12'b011000101011;
   23579: result <= 12'b011000101011;
   23580: result <= 12'b011000101011;
   23581: result <= 12'b011000101011;
   23582: result <= 12'b011000101011;
   23583: result <= 12'b011000101011;
   23584: result <= 12'b011000101011;
   23585: result <= 12'b011000101011;
   23586: result <= 12'b011000101010;
   23587: result <= 12'b011000101010;
   23588: result <= 12'b011000101010;
   23589: result <= 12'b011000101010;
   23590: result <= 12'b011000101010;
   23591: result <= 12'b011000101010;
   23592: result <= 12'b011000101010;
   23593: result <= 12'b011000101010;
   23594: result <= 12'b011000101001;
   23595: result <= 12'b011000101001;
   23596: result <= 12'b011000101001;
   23597: result <= 12'b011000101001;
   23598: result <= 12'b011000101001;
   23599: result <= 12'b011000101001;
   23600: result <= 12'b011000101001;
   23601: result <= 12'b011000101001;
   23602: result <= 12'b011000101000;
   23603: result <= 12'b011000101000;
   23604: result <= 12'b011000101000;
   23605: result <= 12'b011000101000;
   23606: result <= 12'b011000101000;
   23607: result <= 12'b011000101000;
   23608: result <= 12'b011000101000;
   23609: result <= 12'b011000101000;
   23610: result <= 12'b011000100111;
   23611: result <= 12'b011000100111;
   23612: result <= 12'b011000100111;
   23613: result <= 12'b011000100111;
   23614: result <= 12'b011000100111;
   23615: result <= 12'b011000100111;
   23616: result <= 12'b011000100111;
   23617: result <= 12'b011000100110;
   23618: result <= 12'b011000100110;
   23619: result <= 12'b011000100110;
   23620: result <= 12'b011000100110;
   23621: result <= 12'b011000100110;
   23622: result <= 12'b011000100110;
   23623: result <= 12'b011000100110;
   23624: result <= 12'b011000100110;
   23625: result <= 12'b011000100101;
   23626: result <= 12'b011000100101;
   23627: result <= 12'b011000100101;
   23628: result <= 12'b011000100101;
   23629: result <= 12'b011000100101;
   23630: result <= 12'b011000100101;
   23631: result <= 12'b011000100101;
   23632: result <= 12'b011000100101;
   23633: result <= 12'b011000100100;
   23634: result <= 12'b011000100100;
   23635: result <= 12'b011000100100;
   23636: result <= 12'b011000100100;
   23637: result <= 12'b011000100100;
   23638: result <= 12'b011000100100;
   23639: result <= 12'b011000100100;
   23640: result <= 12'b011000100100;
   23641: result <= 12'b011000100011;
   23642: result <= 12'b011000100011;
   23643: result <= 12'b011000100011;
   23644: result <= 12'b011000100011;
   23645: result <= 12'b011000100011;
   23646: result <= 12'b011000100011;
   23647: result <= 12'b011000100011;
   23648: result <= 12'b011000100011;
   23649: result <= 12'b011000100010;
   23650: result <= 12'b011000100010;
   23651: result <= 12'b011000100010;
   23652: result <= 12'b011000100010;
   23653: result <= 12'b011000100010;
   23654: result <= 12'b011000100010;
   23655: result <= 12'b011000100010;
   23656: result <= 12'b011000100010;
   23657: result <= 12'b011000100001;
   23658: result <= 12'b011000100001;
   23659: result <= 12'b011000100001;
   23660: result <= 12'b011000100001;
   23661: result <= 12'b011000100001;
   23662: result <= 12'b011000100001;
   23663: result <= 12'b011000100001;
   23664: result <= 12'b011000100001;
   23665: result <= 12'b011000100000;
   23666: result <= 12'b011000100000;
   23667: result <= 12'b011000100000;
   23668: result <= 12'b011000100000;
   23669: result <= 12'b011000100000;
   23670: result <= 12'b011000100000;
   23671: result <= 12'b011000100000;
   23672: result <= 12'b011000100000;
   23673: result <= 12'b011000011111;
   23674: result <= 12'b011000011111;
   23675: result <= 12'b011000011111;
   23676: result <= 12'b011000011111;
   23677: result <= 12'b011000011111;
   23678: result <= 12'b011000011111;
   23679: result <= 12'b011000011111;
   23680: result <= 12'b011000011111;
   23681: result <= 12'b011000011110;
   23682: result <= 12'b011000011110;
   23683: result <= 12'b011000011110;
   23684: result <= 12'b011000011110;
   23685: result <= 12'b011000011110;
   23686: result <= 12'b011000011110;
   23687: result <= 12'b011000011110;
   23688: result <= 12'b011000011110;
   23689: result <= 12'b011000011101;
   23690: result <= 12'b011000011101;
   23691: result <= 12'b011000011101;
   23692: result <= 12'b011000011101;
   23693: result <= 12'b011000011101;
   23694: result <= 12'b011000011101;
   23695: result <= 12'b011000011101;
   23696: result <= 12'b011000011101;
   23697: result <= 12'b011000011100;
   23698: result <= 12'b011000011100;
   23699: result <= 12'b011000011100;
   23700: result <= 12'b011000011100;
   23701: result <= 12'b011000011100;
   23702: result <= 12'b011000011100;
   23703: result <= 12'b011000011100;
   23704: result <= 12'b011000011100;
   23705: result <= 12'b011000011011;
   23706: result <= 12'b011000011011;
   23707: result <= 12'b011000011011;
   23708: result <= 12'b011000011011;
   23709: result <= 12'b011000011011;
   23710: result <= 12'b011000011011;
   23711: result <= 12'b011000011011;
   23712: result <= 12'b011000011011;
   23713: result <= 12'b011000011010;
   23714: result <= 12'b011000011010;
   23715: result <= 12'b011000011010;
   23716: result <= 12'b011000011010;
   23717: result <= 12'b011000011010;
   23718: result <= 12'b011000011010;
   23719: result <= 12'b011000011010;
   23720: result <= 12'b011000011001;
   23721: result <= 12'b011000011001;
   23722: result <= 12'b011000011001;
   23723: result <= 12'b011000011001;
   23724: result <= 12'b011000011001;
   23725: result <= 12'b011000011001;
   23726: result <= 12'b011000011001;
   23727: result <= 12'b011000011001;
   23728: result <= 12'b011000011000;
   23729: result <= 12'b011000011000;
   23730: result <= 12'b011000011000;
   23731: result <= 12'b011000011000;
   23732: result <= 12'b011000011000;
   23733: result <= 12'b011000011000;
   23734: result <= 12'b011000011000;
   23735: result <= 12'b011000011000;
   23736: result <= 12'b011000010111;
   23737: result <= 12'b011000010111;
   23738: result <= 12'b011000010111;
   23739: result <= 12'b011000010111;
   23740: result <= 12'b011000010111;
   23741: result <= 12'b011000010111;
   23742: result <= 12'b011000010111;
   23743: result <= 12'b011000010111;
   23744: result <= 12'b011000010110;
   23745: result <= 12'b011000010110;
   23746: result <= 12'b011000010110;
   23747: result <= 12'b011000010110;
   23748: result <= 12'b011000010110;
   23749: result <= 12'b011000010110;
   23750: result <= 12'b011000010110;
   23751: result <= 12'b011000010110;
   23752: result <= 12'b011000010101;
   23753: result <= 12'b011000010101;
   23754: result <= 12'b011000010101;
   23755: result <= 12'b011000010101;
   23756: result <= 12'b011000010101;
   23757: result <= 12'b011000010101;
   23758: result <= 12'b011000010101;
   23759: result <= 12'b011000010101;
   23760: result <= 12'b011000010100;
   23761: result <= 12'b011000010100;
   23762: result <= 12'b011000010100;
   23763: result <= 12'b011000010100;
   23764: result <= 12'b011000010100;
   23765: result <= 12'b011000010100;
   23766: result <= 12'b011000010100;
   23767: result <= 12'b011000010100;
   23768: result <= 12'b011000010011;
   23769: result <= 12'b011000010011;
   23770: result <= 12'b011000010011;
   23771: result <= 12'b011000010011;
   23772: result <= 12'b011000010011;
   23773: result <= 12'b011000010011;
   23774: result <= 12'b011000010011;
   23775: result <= 12'b011000010010;
   23776: result <= 12'b011000010010;
   23777: result <= 12'b011000010010;
   23778: result <= 12'b011000010010;
   23779: result <= 12'b011000010010;
   23780: result <= 12'b011000010010;
   23781: result <= 12'b011000010010;
   23782: result <= 12'b011000010010;
   23783: result <= 12'b011000010001;
   23784: result <= 12'b011000010001;
   23785: result <= 12'b011000010001;
   23786: result <= 12'b011000010001;
   23787: result <= 12'b011000010001;
   23788: result <= 12'b011000010001;
   23789: result <= 12'b011000010001;
   23790: result <= 12'b011000010001;
   23791: result <= 12'b011000010000;
   23792: result <= 12'b011000010000;
   23793: result <= 12'b011000010000;
   23794: result <= 12'b011000010000;
   23795: result <= 12'b011000010000;
   23796: result <= 12'b011000010000;
   23797: result <= 12'b011000010000;
   23798: result <= 12'b011000010000;
   23799: result <= 12'b011000001111;
   23800: result <= 12'b011000001111;
   23801: result <= 12'b011000001111;
   23802: result <= 12'b011000001111;
   23803: result <= 12'b011000001111;
   23804: result <= 12'b011000001111;
   23805: result <= 12'b011000001111;
   23806: result <= 12'b011000001111;
   23807: result <= 12'b011000001110;
   23808: result <= 12'b011000001110;
   23809: result <= 12'b011000001110;
   23810: result <= 12'b011000001110;
   23811: result <= 12'b011000001110;
   23812: result <= 12'b011000001110;
   23813: result <= 12'b011000001110;
   23814: result <= 12'b011000001101;
   23815: result <= 12'b011000001101;
   23816: result <= 12'b011000001101;
   23817: result <= 12'b011000001101;
   23818: result <= 12'b011000001101;
   23819: result <= 12'b011000001101;
   23820: result <= 12'b011000001101;
   23821: result <= 12'b011000001101;
   23822: result <= 12'b011000001100;
   23823: result <= 12'b011000001100;
   23824: result <= 12'b011000001100;
   23825: result <= 12'b011000001100;
   23826: result <= 12'b011000001100;
   23827: result <= 12'b011000001100;
   23828: result <= 12'b011000001100;
   23829: result <= 12'b011000001100;
   23830: result <= 12'b011000001011;
   23831: result <= 12'b011000001011;
   23832: result <= 12'b011000001011;
   23833: result <= 12'b011000001011;
   23834: result <= 12'b011000001011;
   23835: result <= 12'b011000001011;
   23836: result <= 12'b011000001011;
   23837: result <= 12'b011000001011;
   23838: result <= 12'b011000001010;
   23839: result <= 12'b011000001010;
   23840: result <= 12'b011000001010;
   23841: result <= 12'b011000001010;
   23842: result <= 12'b011000001010;
   23843: result <= 12'b011000001010;
   23844: result <= 12'b011000001010;
   23845: result <= 12'b011000001010;
   23846: result <= 12'b011000001001;
   23847: result <= 12'b011000001001;
   23848: result <= 12'b011000001001;
   23849: result <= 12'b011000001001;
   23850: result <= 12'b011000001001;
   23851: result <= 12'b011000001001;
   23852: result <= 12'b011000001001;
   23853: result <= 12'b011000001000;
   23854: result <= 12'b011000001000;
   23855: result <= 12'b011000001000;
   23856: result <= 12'b011000001000;
   23857: result <= 12'b011000001000;
   23858: result <= 12'b011000001000;
   23859: result <= 12'b011000001000;
   23860: result <= 12'b011000001000;
   23861: result <= 12'b011000000111;
   23862: result <= 12'b011000000111;
   23863: result <= 12'b011000000111;
   23864: result <= 12'b011000000111;
   23865: result <= 12'b011000000111;
   23866: result <= 12'b011000000111;
   23867: result <= 12'b011000000111;
   23868: result <= 12'b011000000111;
   23869: result <= 12'b011000000110;
   23870: result <= 12'b011000000110;
   23871: result <= 12'b011000000110;
   23872: result <= 12'b011000000110;
   23873: result <= 12'b011000000110;
   23874: result <= 12'b011000000110;
   23875: result <= 12'b011000000110;
   23876: result <= 12'b011000000110;
   23877: result <= 12'b011000000101;
   23878: result <= 12'b011000000101;
   23879: result <= 12'b011000000101;
   23880: result <= 12'b011000000101;
   23881: result <= 12'b011000000101;
   23882: result <= 12'b011000000101;
   23883: result <= 12'b011000000101;
   23884: result <= 12'b011000000100;
   23885: result <= 12'b011000000100;
   23886: result <= 12'b011000000100;
   23887: result <= 12'b011000000100;
   23888: result <= 12'b011000000100;
   23889: result <= 12'b011000000100;
   23890: result <= 12'b011000000100;
   23891: result <= 12'b011000000100;
   23892: result <= 12'b011000000011;
   23893: result <= 12'b011000000011;
   23894: result <= 12'b011000000011;
   23895: result <= 12'b011000000011;
   23896: result <= 12'b011000000011;
   23897: result <= 12'b011000000011;
   23898: result <= 12'b011000000011;
   23899: result <= 12'b011000000011;
   23900: result <= 12'b011000000010;
   23901: result <= 12'b011000000010;
   23902: result <= 12'b011000000010;
   23903: result <= 12'b011000000010;
   23904: result <= 12'b011000000010;
   23905: result <= 12'b011000000010;
   23906: result <= 12'b011000000010;
   23907: result <= 12'b011000000001;
   23908: result <= 12'b011000000001;
   23909: result <= 12'b011000000001;
   23910: result <= 12'b011000000001;
   23911: result <= 12'b011000000001;
   23912: result <= 12'b011000000001;
   23913: result <= 12'b011000000001;
   23914: result <= 12'b011000000001;
   23915: result <= 12'b011000000000;
   23916: result <= 12'b011000000000;
   23917: result <= 12'b011000000000;
   23918: result <= 12'b011000000000;
   23919: result <= 12'b011000000000;
   23920: result <= 12'b011000000000;
   23921: result <= 12'b011000000000;
   23922: result <= 12'b011000000000;
   23923: result <= 12'b010111111111;
   23924: result <= 12'b010111111111;
   23925: result <= 12'b010111111111;
   23926: result <= 12'b010111111111;
   23927: result <= 12'b010111111111;
   23928: result <= 12'b010111111111;
   23929: result <= 12'b010111111111;
   23930: result <= 12'b010111111111;
   23931: result <= 12'b010111111110;
   23932: result <= 12'b010111111110;
   23933: result <= 12'b010111111110;
   23934: result <= 12'b010111111110;
   23935: result <= 12'b010111111110;
   23936: result <= 12'b010111111110;
   23937: result <= 12'b010111111110;
   23938: result <= 12'b010111111101;
   23939: result <= 12'b010111111101;
   23940: result <= 12'b010111111101;
   23941: result <= 12'b010111111101;
   23942: result <= 12'b010111111101;
   23943: result <= 12'b010111111101;
   23944: result <= 12'b010111111101;
   23945: result <= 12'b010111111101;
   23946: result <= 12'b010111111100;
   23947: result <= 12'b010111111100;
   23948: result <= 12'b010111111100;
   23949: result <= 12'b010111111100;
   23950: result <= 12'b010111111100;
   23951: result <= 12'b010111111100;
   23952: result <= 12'b010111111100;
   23953: result <= 12'b010111111100;
   23954: result <= 12'b010111111011;
   23955: result <= 12'b010111111011;
   23956: result <= 12'b010111111011;
   23957: result <= 12'b010111111011;
   23958: result <= 12'b010111111011;
   23959: result <= 12'b010111111011;
   23960: result <= 12'b010111111011;
   23961: result <= 12'b010111111010;
   23962: result <= 12'b010111111010;
   23963: result <= 12'b010111111010;
   23964: result <= 12'b010111111010;
   23965: result <= 12'b010111111010;
   23966: result <= 12'b010111111010;
   23967: result <= 12'b010111111010;
   23968: result <= 12'b010111111010;
   23969: result <= 12'b010111111001;
   23970: result <= 12'b010111111001;
   23971: result <= 12'b010111111001;
   23972: result <= 12'b010111111001;
   23973: result <= 12'b010111111001;
   23974: result <= 12'b010111111001;
   23975: result <= 12'b010111111001;
   23976: result <= 12'b010111111001;
   23977: result <= 12'b010111111000;
   23978: result <= 12'b010111111000;
   23979: result <= 12'b010111111000;
   23980: result <= 12'b010111111000;
   23981: result <= 12'b010111111000;
   23982: result <= 12'b010111111000;
   23983: result <= 12'b010111111000;
   23984: result <= 12'b010111110111;
   23985: result <= 12'b010111110111;
   23986: result <= 12'b010111110111;
   23987: result <= 12'b010111110111;
   23988: result <= 12'b010111110111;
   23989: result <= 12'b010111110111;
   23990: result <= 12'b010111110111;
   23991: result <= 12'b010111110111;
   23992: result <= 12'b010111110110;
   23993: result <= 12'b010111110110;
   23994: result <= 12'b010111110110;
   23995: result <= 12'b010111110110;
   23996: result <= 12'b010111110110;
   23997: result <= 12'b010111110110;
   23998: result <= 12'b010111110110;
   23999: result <= 12'b010111110110;
   24000: result <= 12'b010111110101;
   24001: result <= 12'b010111110101;
   24002: result <= 12'b010111110101;
   24003: result <= 12'b010111110101;
   24004: result <= 12'b010111110101;
   24005: result <= 12'b010111110101;
   24006: result <= 12'b010111110101;
   24007: result <= 12'b010111110100;
   24008: result <= 12'b010111110100;
   24009: result <= 12'b010111110100;
   24010: result <= 12'b010111110100;
   24011: result <= 12'b010111110100;
   24012: result <= 12'b010111110100;
   24013: result <= 12'b010111110100;
   24014: result <= 12'b010111110100;
   24015: result <= 12'b010111110011;
   24016: result <= 12'b010111110011;
   24017: result <= 12'b010111110011;
   24018: result <= 12'b010111110011;
   24019: result <= 12'b010111110011;
   24020: result <= 12'b010111110011;
   24021: result <= 12'b010111110011;
   24022: result <= 12'b010111110010;
   24023: result <= 12'b010111110010;
   24024: result <= 12'b010111110010;
   24025: result <= 12'b010111110010;
   24026: result <= 12'b010111110010;
   24027: result <= 12'b010111110010;
   24028: result <= 12'b010111110010;
   24029: result <= 12'b010111110010;
   24030: result <= 12'b010111110001;
   24031: result <= 12'b010111110001;
   24032: result <= 12'b010111110001;
   24033: result <= 12'b010111110001;
   24034: result <= 12'b010111110001;
   24035: result <= 12'b010111110001;
   24036: result <= 12'b010111110001;
   24037: result <= 12'b010111110001;
   24038: result <= 12'b010111110000;
   24039: result <= 12'b010111110000;
   24040: result <= 12'b010111110000;
   24041: result <= 12'b010111110000;
   24042: result <= 12'b010111110000;
   24043: result <= 12'b010111110000;
   24044: result <= 12'b010111110000;
   24045: result <= 12'b010111101111;
   24046: result <= 12'b010111101111;
   24047: result <= 12'b010111101111;
   24048: result <= 12'b010111101111;
   24049: result <= 12'b010111101111;
   24050: result <= 12'b010111101111;
   24051: result <= 12'b010111101111;
   24052: result <= 12'b010111101111;
   24053: result <= 12'b010111101110;
   24054: result <= 12'b010111101110;
   24055: result <= 12'b010111101110;
   24056: result <= 12'b010111101110;
   24057: result <= 12'b010111101110;
   24058: result <= 12'b010111101110;
   24059: result <= 12'b010111101110;
   24060: result <= 12'b010111101101;
   24061: result <= 12'b010111101101;
   24062: result <= 12'b010111101101;
   24063: result <= 12'b010111101101;
   24064: result <= 12'b010111101101;
   24065: result <= 12'b010111101101;
   24066: result <= 12'b010111101101;
   24067: result <= 12'b010111101101;
   24068: result <= 12'b010111101100;
   24069: result <= 12'b010111101100;
   24070: result <= 12'b010111101100;
   24071: result <= 12'b010111101100;
   24072: result <= 12'b010111101100;
   24073: result <= 12'b010111101100;
   24074: result <= 12'b010111101100;
   24075: result <= 12'b010111101100;
   24076: result <= 12'b010111101011;
   24077: result <= 12'b010111101011;
   24078: result <= 12'b010111101011;
   24079: result <= 12'b010111101011;
   24080: result <= 12'b010111101011;
   24081: result <= 12'b010111101011;
   24082: result <= 12'b010111101011;
   24083: result <= 12'b010111101010;
   24084: result <= 12'b010111101010;
   24085: result <= 12'b010111101010;
   24086: result <= 12'b010111101010;
   24087: result <= 12'b010111101010;
   24088: result <= 12'b010111101010;
   24089: result <= 12'b010111101010;
   24090: result <= 12'b010111101010;
   24091: result <= 12'b010111101001;
   24092: result <= 12'b010111101001;
   24093: result <= 12'b010111101001;
   24094: result <= 12'b010111101001;
   24095: result <= 12'b010111101001;
   24096: result <= 12'b010111101001;
   24097: result <= 12'b010111101001;
   24098: result <= 12'b010111101000;
   24099: result <= 12'b010111101000;
   24100: result <= 12'b010111101000;
   24101: result <= 12'b010111101000;
   24102: result <= 12'b010111101000;
   24103: result <= 12'b010111101000;
   24104: result <= 12'b010111101000;
   24105: result <= 12'b010111101000;
   24106: result <= 12'b010111100111;
   24107: result <= 12'b010111100111;
   24108: result <= 12'b010111100111;
   24109: result <= 12'b010111100111;
   24110: result <= 12'b010111100111;
   24111: result <= 12'b010111100111;
   24112: result <= 12'b010111100111;
   24113: result <= 12'b010111100110;
   24114: result <= 12'b010111100110;
   24115: result <= 12'b010111100110;
   24116: result <= 12'b010111100110;
   24117: result <= 12'b010111100110;
   24118: result <= 12'b010111100110;
   24119: result <= 12'b010111100110;
   24120: result <= 12'b010111100110;
   24121: result <= 12'b010111100101;
   24122: result <= 12'b010111100101;
   24123: result <= 12'b010111100101;
   24124: result <= 12'b010111100101;
   24125: result <= 12'b010111100101;
   24126: result <= 12'b010111100101;
   24127: result <= 12'b010111100101;
   24128: result <= 12'b010111100101;
   24129: result <= 12'b010111100100;
   24130: result <= 12'b010111100100;
   24131: result <= 12'b010111100100;
   24132: result <= 12'b010111100100;
   24133: result <= 12'b010111100100;
   24134: result <= 12'b010111100100;
   24135: result <= 12'b010111100100;
   24136: result <= 12'b010111100011;
   24137: result <= 12'b010111100011;
   24138: result <= 12'b010111100011;
   24139: result <= 12'b010111100011;
   24140: result <= 12'b010111100011;
   24141: result <= 12'b010111100011;
   24142: result <= 12'b010111100011;
   24143: result <= 12'b010111100011;
   24144: result <= 12'b010111100010;
   24145: result <= 12'b010111100010;
   24146: result <= 12'b010111100010;
   24147: result <= 12'b010111100010;
   24148: result <= 12'b010111100010;
   24149: result <= 12'b010111100010;
   24150: result <= 12'b010111100010;
   24151: result <= 12'b010111100001;
   24152: result <= 12'b010111100001;
   24153: result <= 12'b010111100001;
   24154: result <= 12'b010111100001;
   24155: result <= 12'b010111100001;
   24156: result <= 12'b010111100001;
   24157: result <= 12'b010111100001;
   24158: result <= 12'b010111100001;
   24159: result <= 12'b010111100000;
   24160: result <= 12'b010111100000;
   24161: result <= 12'b010111100000;
   24162: result <= 12'b010111100000;
   24163: result <= 12'b010111100000;
   24164: result <= 12'b010111100000;
   24165: result <= 12'b010111100000;
   24166: result <= 12'b010111011111;
   24167: result <= 12'b010111011111;
   24168: result <= 12'b010111011111;
   24169: result <= 12'b010111011111;
   24170: result <= 12'b010111011111;
   24171: result <= 12'b010111011111;
   24172: result <= 12'b010111011111;
   24173: result <= 12'b010111011111;
   24174: result <= 12'b010111011110;
   24175: result <= 12'b010111011110;
   24176: result <= 12'b010111011110;
   24177: result <= 12'b010111011110;
   24178: result <= 12'b010111011110;
   24179: result <= 12'b010111011110;
   24180: result <= 12'b010111011110;
   24181: result <= 12'b010111011101;
   24182: result <= 12'b010111011101;
   24183: result <= 12'b010111011101;
   24184: result <= 12'b010111011101;
   24185: result <= 12'b010111011101;
   24186: result <= 12'b010111011101;
   24187: result <= 12'b010111011101;
   24188: result <= 12'b010111011101;
   24189: result <= 12'b010111011100;
   24190: result <= 12'b010111011100;
   24191: result <= 12'b010111011100;
   24192: result <= 12'b010111011100;
   24193: result <= 12'b010111011100;
   24194: result <= 12'b010111011100;
   24195: result <= 12'b010111011100;
   24196: result <= 12'b010111011011;
   24197: result <= 12'b010111011011;
   24198: result <= 12'b010111011011;
   24199: result <= 12'b010111011011;
   24200: result <= 12'b010111011011;
   24201: result <= 12'b010111011011;
   24202: result <= 12'b010111011011;
   24203: result <= 12'b010111011011;
   24204: result <= 12'b010111011010;
   24205: result <= 12'b010111011010;
   24206: result <= 12'b010111011010;
   24207: result <= 12'b010111011010;
   24208: result <= 12'b010111011010;
   24209: result <= 12'b010111011010;
   24210: result <= 12'b010111011010;
   24211: result <= 12'b010111011001;
   24212: result <= 12'b010111011001;
   24213: result <= 12'b010111011001;
   24214: result <= 12'b010111011001;
   24215: result <= 12'b010111011001;
   24216: result <= 12'b010111011001;
   24217: result <= 12'b010111011001;
   24218: result <= 12'b010111011000;
   24219: result <= 12'b010111011000;
   24220: result <= 12'b010111011000;
   24221: result <= 12'b010111011000;
   24222: result <= 12'b010111011000;
   24223: result <= 12'b010111011000;
   24224: result <= 12'b010111011000;
   24225: result <= 12'b010111011000;
   24226: result <= 12'b010111010111;
   24227: result <= 12'b010111010111;
   24228: result <= 12'b010111010111;
   24229: result <= 12'b010111010111;
   24230: result <= 12'b010111010111;
   24231: result <= 12'b010111010111;
   24232: result <= 12'b010111010111;
   24233: result <= 12'b010111010110;
   24234: result <= 12'b010111010110;
   24235: result <= 12'b010111010110;
   24236: result <= 12'b010111010110;
   24237: result <= 12'b010111010110;
   24238: result <= 12'b010111010110;
   24239: result <= 12'b010111010110;
   24240: result <= 12'b010111010110;
   24241: result <= 12'b010111010101;
   24242: result <= 12'b010111010101;
   24243: result <= 12'b010111010101;
   24244: result <= 12'b010111010101;
   24245: result <= 12'b010111010101;
   24246: result <= 12'b010111010101;
   24247: result <= 12'b010111010101;
   24248: result <= 12'b010111010100;
   24249: result <= 12'b010111010100;
   24250: result <= 12'b010111010100;
   24251: result <= 12'b010111010100;
   24252: result <= 12'b010111010100;
   24253: result <= 12'b010111010100;
   24254: result <= 12'b010111010100;
   24255: result <= 12'b010111010100;
   24256: result <= 12'b010111010011;
   24257: result <= 12'b010111010011;
   24258: result <= 12'b010111010011;
   24259: result <= 12'b010111010011;
   24260: result <= 12'b010111010011;
   24261: result <= 12'b010111010011;
   24262: result <= 12'b010111010011;
   24263: result <= 12'b010111010010;
   24264: result <= 12'b010111010010;
   24265: result <= 12'b010111010010;
   24266: result <= 12'b010111010010;
   24267: result <= 12'b010111010010;
   24268: result <= 12'b010111010010;
   24269: result <= 12'b010111010010;
   24270: result <= 12'b010111010010;
   24271: result <= 12'b010111010001;
   24272: result <= 12'b010111010001;
   24273: result <= 12'b010111010001;
   24274: result <= 12'b010111010001;
   24275: result <= 12'b010111010001;
   24276: result <= 12'b010111010001;
   24277: result <= 12'b010111010001;
   24278: result <= 12'b010111010000;
   24279: result <= 12'b010111010000;
   24280: result <= 12'b010111010000;
   24281: result <= 12'b010111010000;
   24282: result <= 12'b010111010000;
   24283: result <= 12'b010111010000;
   24284: result <= 12'b010111010000;
   24285: result <= 12'b010111001111;
   24286: result <= 12'b010111001111;
   24287: result <= 12'b010111001111;
   24288: result <= 12'b010111001111;
   24289: result <= 12'b010111001111;
   24290: result <= 12'b010111001111;
   24291: result <= 12'b010111001111;
   24292: result <= 12'b010111001111;
   24293: result <= 12'b010111001110;
   24294: result <= 12'b010111001110;
   24295: result <= 12'b010111001110;
   24296: result <= 12'b010111001110;
   24297: result <= 12'b010111001110;
   24298: result <= 12'b010111001110;
   24299: result <= 12'b010111001110;
   24300: result <= 12'b010111001101;
   24301: result <= 12'b010111001101;
   24302: result <= 12'b010111001101;
   24303: result <= 12'b010111001101;
   24304: result <= 12'b010111001101;
   24305: result <= 12'b010111001101;
   24306: result <= 12'b010111001101;
   24307: result <= 12'b010111001101;
   24308: result <= 12'b010111001100;
   24309: result <= 12'b010111001100;
   24310: result <= 12'b010111001100;
   24311: result <= 12'b010111001100;
   24312: result <= 12'b010111001100;
   24313: result <= 12'b010111001100;
   24314: result <= 12'b010111001100;
   24315: result <= 12'b010111001011;
   24316: result <= 12'b010111001011;
   24317: result <= 12'b010111001011;
   24318: result <= 12'b010111001011;
   24319: result <= 12'b010111001011;
   24320: result <= 12'b010111001011;
   24321: result <= 12'b010111001011;
   24322: result <= 12'b010111001010;
   24323: result <= 12'b010111001010;
   24324: result <= 12'b010111001010;
   24325: result <= 12'b010111001010;
   24326: result <= 12'b010111001010;
   24327: result <= 12'b010111001010;
   24328: result <= 12'b010111001010;
   24329: result <= 12'b010111001010;
   24330: result <= 12'b010111001001;
   24331: result <= 12'b010111001001;
   24332: result <= 12'b010111001001;
   24333: result <= 12'b010111001001;
   24334: result <= 12'b010111001001;
   24335: result <= 12'b010111001001;
   24336: result <= 12'b010111001001;
   24337: result <= 12'b010111001000;
   24338: result <= 12'b010111001000;
   24339: result <= 12'b010111001000;
   24340: result <= 12'b010111001000;
   24341: result <= 12'b010111001000;
   24342: result <= 12'b010111001000;
   24343: result <= 12'b010111001000;
   24344: result <= 12'b010111001000;
   24345: result <= 12'b010111000111;
   24346: result <= 12'b010111000111;
   24347: result <= 12'b010111000111;
   24348: result <= 12'b010111000111;
   24349: result <= 12'b010111000111;
   24350: result <= 12'b010111000111;
   24351: result <= 12'b010111000111;
   24352: result <= 12'b010111000110;
   24353: result <= 12'b010111000110;
   24354: result <= 12'b010111000110;
   24355: result <= 12'b010111000110;
   24356: result <= 12'b010111000110;
   24357: result <= 12'b010111000110;
   24358: result <= 12'b010111000110;
   24359: result <= 12'b010111000101;
   24360: result <= 12'b010111000101;
   24361: result <= 12'b010111000101;
   24362: result <= 12'b010111000101;
   24363: result <= 12'b010111000101;
   24364: result <= 12'b010111000101;
   24365: result <= 12'b010111000101;
   24366: result <= 12'b010111000101;
   24367: result <= 12'b010111000100;
   24368: result <= 12'b010111000100;
   24369: result <= 12'b010111000100;
   24370: result <= 12'b010111000100;
   24371: result <= 12'b010111000100;
   24372: result <= 12'b010111000100;
   24373: result <= 12'b010111000100;
   24374: result <= 12'b010111000011;
   24375: result <= 12'b010111000011;
   24376: result <= 12'b010111000011;
   24377: result <= 12'b010111000011;
   24378: result <= 12'b010111000011;
   24379: result <= 12'b010111000011;
   24380: result <= 12'b010111000011;
   24381: result <= 12'b010111000010;
   24382: result <= 12'b010111000010;
   24383: result <= 12'b010111000010;
   24384: result <= 12'b010111000010;
   24385: result <= 12'b010111000010;
   24386: result <= 12'b010111000010;
   24387: result <= 12'b010111000010;
   24388: result <= 12'b010111000010;
   24389: result <= 12'b010111000001;
   24390: result <= 12'b010111000001;
   24391: result <= 12'b010111000001;
   24392: result <= 12'b010111000001;
   24393: result <= 12'b010111000001;
   24394: result <= 12'b010111000001;
   24395: result <= 12'b010111000001;
   24396: result <= 12'b010111000000;
   24397: result <= 12'b010111000000;
   24398: result <= 12'b010111000000;
   24399: result <= 12'b010111000000;
   24400: result <= 12'b010111000000;
   24401: result <= 12'b010111000000;
   24402: result <= 12'b010111000000;
   24403: result <= 12'b010110111111;
   24404: result <= 12'b010110111111;
   24405: result <= 12'b010110111111;
   24406: result <= 12'b010110111111;
   24407: result <= 12'b010110111111;
   24408: result <= 12'b010110111111;
   24409: result <= 12'b010110111111;
   24410: result <= 12'b010110111111;
   24411: result <= 12'b010110111110;
   24412: result <= 12'b010110111110;
   24413: result <= 12'b010110111110;
   24414: result <= 12'b010110111110;
   24415: result <= 12'b010110111110;
   24416: result <= 12'b010110111110;
   24417: result <= 12'b010110111110;
   24418: result <= 12'b010110111101;
   24419: result <= 12'b010110111101;
   24420: result <= 12'b010110111101;
   24421: result <= 12'b010110111101;
   24422: result <= 12'b010110111101;
   24423: result <= 12'b010110111101;
   24424: result <= 12'b010110111101;
   24425: result <= 12'b010110111100;
   24426: result <= 12'b010110111100;
   24427: result <= 12'b010110111100;
   24428: result <= 12'b010110111100;
   24429: result <= 12'b010110111100;
   24430: result <= 12'b010110111100;
   24431: result <= 12'b010110111100;
   24432: result <= 12'b010110111100;
   24433: result <= 12'b010110111011;
   24434: result <= 12'b010110111011;
   24435: result <= 12'b010110111011;
   24436: result <= 12'b010110111011;
   24437: result <= 12'b010110111011;
   24438: result <= 12'b010110111011;
   24439: result <= 12'b010110111011;
   24440: result <= 12'b010110111010;
   24441: result <= 12'b010110111010;
   24442: result <= 12'b010110111010;
   24443: result <= 12'b010110111010;
   24444: result <= 12'b010110111010;
   24445: result <= 12'b010110111010;
   24446: result <= 12'b010110111010;
   24447: result <= 12'b010110111001;
   24448: result <= 12'b010110111001;
   24449: result <= 12'b010110111001;
   24450: result <= 12'b010110111001;
   24451: result <= 12'b010110111001;
   24452: result <= 12'b010110111001;
   24453: result <= 12'b010110111001;
   24454: result <= 12'b010110111000;
   24455: result <= 12'b010110111000;
   24456: result <= 12'b010110111000;
   24457: result <= 12'b010110111000;
   24458: result <= 12'b010110111000;
   24459: result <= 12'b010110111000;
   24460: result <= 12'b010110111000;
   24461: result <= 12'b010110111000;
   24462: result <= 12'b010110110111;
   24463: result <= 12'b010110110111;
   24464: result <= 12'b010110110111;
   24465: result <= 12'b010110110111;
   24466: result <= 12'b010110110111;
   24467: result <= 12'b010110110111;
   24468: result <= 12'b010110110111;
   24469: result <= 12'b010110110110;
   24470: result <= 12'b010110110110;
   24471: result <= 12'b010110110110;
   24472: result <= 12'b010110110110;
   24473: result <= 12'b010110110110;
   24474: result <= 12'b010110110110;
   24475: result <= 12'b010110110110;
   24476: result <= 12'b010110110101;
   24477: result <= 12'b010110110101;
   24478: result <= 12'b010110110101;
   24479: result <= 12'b010110110101;
   24480: result <= 12'b010110110101;
   24481: result <= 12'b010110110101;
   24482: result <= 12'b010110110101;
   24483: result <= 12'b010110110101;
   24484: result <= 12'b010110110100;
   24485: result <= 12'b010110110100;
   24486: result <= 12'b010110110100;
   24487: result <= 12'b010110110100;
   24488: result <= 12'b010110110100;
   24489: result <= 12'b010110110100;
   24490: result <= 12'b010110110100;
   24491: result <= 12'b010110110011;
   24492: result <= 12'b010110110011;
   24493: result <= 12'b010110110011;
   24494: result <= 12'b010110110011;
   24495: result <= 12'b010110110011;
   24496: result <= 12'b010110110011;
   24497: result <= 12'b010110110011;
   24498: result <= 12'b010110110010;
   24499: result <= 12'b010110110010;
   24500: result <= 12'b010110110010;
   24501: result <= 12'b010110110010;
   24502: result <= 12'b010110110010;
   24503: result <= 12'b010110110010;
   24504: result <= 12'b010110110010;
   24505: result <= 12'b010110110001;
   24506: result <= 12'b010110110001;
   24507: result <= 12'b010110110001;
   24508: result <= 12'b010110110001;
   24509: result <= 12'b010110110001;
   24510: result <= 12'b010110110001;
   24511: result <= 12'b010110110001;
   24512: result <= 12'b010110110001;
   24513: result <= 12'b010110110000;
   24514: result <= 12'b010110110000;
   24515: result <= 12'b010110110000;
   24516: result <= 12'b010110110000;
   24517: result <= 12'b010110110000;
   24518: result <= 12'b010110110000;
   24519: result <= 12'b010110110000;
   24520: result <= 12'b010110101111;
   24521: result <= 12'b010110101111;
   24522: result <= 12'b010110101111;
   24523: result <= 12'b010110101111;
   24524: result <= 12'b010110101111;
   24525: result <= 12'b010110101111;
   24526: result <= 12'b010110101111;
   24527: result <= 12'b010110101110;
   24528: result <= 12'b010110101110;
   24529: result <= 12'b010110101110;
   24530: result <= 12'b010110101110;
   24531: result <= 12'b010110101110;
   24532: result <= 12'b010110101110;
   24533: result <= 12'b010110101110;
   24534: result <= 12'b010110101101;
   24535: result <= 12'b010110101101;
   24536: result <= 12'b010110101101;
   24537: result <= 12'b010110101101;
   24538: result <= 12'b010110101101;
   24539: result <= 12'b010110101101;
   24540: result <= 12'b010110101101;
   24541: result <= 12'b010110101101;
   24542: result <= 12'b010110101100;
   24543: result <= 12'b010110101100;
   24544: result <= 12'b010110101100;
   24545: result <= 12'b010110101100;
   24546: result <= 12'b010110101100;
   24547: result <= 12'b010110101100;
   24548: result <= 12'b010110101100;
   24549: result <= 12'b010110101011;
   24550: result <= 12'b010110101011;
   24551: result <= 12'b010110101011;
   24552: result <= 12'b010110101011;
   24553: result <= 12'b010110101011;
   24554: result <= 12'b010110101011;
   24555: result <= 12'b010110101011;
   24556: result <= 12'b010110101010;
   24557: result <= 12'b010110101010;
   24558: result <= 12'b010110101010;
   24559: result <= 12'b010110101010;
   24560: result <= 12'b010110101010;
   24561: result <= 12'b010110101010;
   24562: result <= 12'b010110101010;
   24563: result <= 12'b010110101001;
   24564: result <= 12'b010110101001;
   24565: result <= 12'b010110101001;
   24566: result <= 12'b010110101001;
   24567: result <= 12'b010110101001;
   24568: result <= 12'b010110101001;
   24569: result <= 12'b010110101001;
   24570: result <= 12'b010110101000;
   24571: result <= 12'b010110101000;
   24572: result <= 12'b010110101000;
   24573: result <= 12'b010110101000;
   24574: result <= 12'b010110101000;
   24575: result <= 12'b010110101000;
   24576: result <= 12'b010110101000;
   24577: result <= 12'b010110101000;
   24578: result <= 12'b010110100111;
   24579: result <= 12'b010110100111;
   24580: result <= 12'b010110100111;
   24581: result <= 12'b010110100111;
   24582: result <= 12'b010110100111;
   24583: result <= 12'b010110100111;
   24584: result <= 12'b010110100111;
   24585: result <= 12'b010110100110;
   24586: result <= 12'b010110100110;
   24587: result <= 12'b010110100110;
   24588: result <= 12'b010110100110;
   24589: result <= 12'b010110100110;
   24590: result <= 12'b010110100110;
   24591: result <= 12'b010110100110;
   24592: result <= 12'b010110100101;
   24593: result <= 12'b010110100101;
   24594: result <= 12'b010110100101;
   24595: result <= 12'b010110100101;
   24596: result <= 12'b010110100101;
   24597: result <= 12'b010110100101;
   24598: result <= 12'b010110100101;
   24599: result <= 12'b010110100100;
   24600: result <= 12'b010110100100;
   24601: result <= 12'b010110100100;
   24602: result <= 12'b010110100100;
   24603: result <= 12'b010110100100;
   24604: result <= 12'b010110100100;
   24605: result <= 12'b010110100100;
   24606: result <= 12'b010110100011;
   24607: result <= 12'b010110100011;
   24608: result <= 12'b010110100011;
   24609: result <= 12'b010110100011;
   24610: result <= 12'b010110100011;
   24611: result <= 12'b010110100011;
   24612: result <= 12'b010110100011;
   24613: result <= 12'b010110100011;
   24614: result <= 12'b010110100010;
   24615: result <= 12'b010110100010;
   24616: result <= 12'b010110100010;
   24617: result <= 12'b010110100010;
   24618: result <= 12'b010110100010;
   24619: result <= 12'b010110100010;
   24620: result <= 12'b010110100010;
   24621: result <= 12'b010110100001;
   24622: result <= 12'b010110100001;
   24623: result <= 12'b010110100001;
   24624: result <= 12'b010110100001;
   24625: result <= 12'b010110100001;
   24626: result <= 12'b010110100001;
   24627: result <= 12'b010110100001;
   24628: result <= 12'b010110100000;
   24629: result <= 12'b010110100000;
   24630: result <= 12'b010110100000;
   24631: result <= 12'b010110100000;
   24632: result <= 12'b010110100000;
   24633: result <= 12'b010110100000;
   24634: result <= 12'b010110100000;
   24635: result <= 12'b010110011111;
   24636: result <= 12'b010110011111;
   24637: result <= 12'b010110011111;
   24638: result <= 12'b010110011111;
   24639: result <= 12'b010110011111;
   24640: result <= 12'b010110011111;
   24641: result <= 12'b010110011111;
   24642: result <= 12'b010110011110;
   24643: result <= 12'b010110011110;
   24644: result <= 12'b010110011110;
   24645: result <= 12'b010110011110;
   24646: result <= 12'b010110011110;
   24647: result <= 12'b010110011110;
   24648: result <= 12'b010110011110;
   24649: result <= 12'b010110011101;
   24650: result <= 12'b010110011101;
   24651: result <= 12'b010110011101;
   24652: result <= 12'b010110011101;
   24653: result <= 12'b010110011101;
   24654: result <= 12'b010110011101;
   24655: result <= 12'b010110011101;
   24656: result <= 12'b010110011101;
   24657: result <= 12'b010110011100;
   24658: result <= 12'b010110011100;
   24659: result <= 12'b010110011100;
   24660: result <= 12'b010110011100;
   24661: result <= 12'b010110011100;
   24662: result <= 12'b010110011100;
   24663: result <= 12'b010110011100;
   24664: result <= 12'b010110011011;
   24665: result <= 12'b010110011011;
   24666: result <= 12'b010110011011;
   24667: result <= 12'b010110011011;
   24668: result <= 12'b010110011011;
   24669: result <= 12'b010110011011;
   24670: result <= 12'b010110011011;
   24671: result <= 12'b010110011010;
   24672: result <= 12'b010110011010;
   24673: result <= 12'b010110011010;
   24674: result <= 12'b010110011010;
   24675: result <= 12'b010110011010;
   24676: result <= 12'b010110011010;
   24677: result <= 12'b010110011010;
   24678: result <= 12'b010110011001;
   24679: result <= 12'b010110011001;
   24680: result <= 12'b010110011001;
   24681: result <= 12'b010110011001;
   24682: result <= 12'b010110011001;
   24683: result <= 12'b010110011001;
   24684: result <= 12'b010110011001;
   24685: result <= 12'b010110011000;
   24686: result <= 12'b010110011000;
   24687: result <= 12'b010110011000;
   24688: result <= 12'b010110011000;
   24689: result <= 12'b010110011000;
   24690: result <= 12'b010110011000;
   24691: result <= 12'b010110011000;
   24692: result <= 12'b010110010111;
   24693: result <= 12'b010110010111;
   24694: result <= 12'b010110010111;
   24695: result <= 12'b010110010111;
   24696: result <= 12'b010110010111;
   24697: result <= 12'b010110010111;
   24698: result <= 12'b010110010111;
   24699: result <= 12'b010110010110;
   24700: result <= 12'b010110010110;
   24701: result <= 12'b010110010110;
   24702: result <= 12'b010110010110;
   24703: result <= 12'b010110010110;
   24704: result <= 12'b010110010110;
   24705: result <= 12'b010110010110;
   24706: result <= 12'b010110010101;
   24707: result <= 12'b010110010101;
   24708: result <= 12'b010110010101;
   24709: result <= 12'b010110010101;
   24710: result <= 12'b010110010101;
   24711: result <= 12'b010110010101;
   24712: result <= 12'b010110010101;
   24713: result <= 12'b010110010101;
   24714: result <= 12'b010110010100;
   24715: result <= 12'b010110010100;
   24716: result <= 12'b010110010100;
   24717: result <= 12'b010110010100;
   24718: result <= 12'b010110010100;
   24719: result <= 12'b010110010100;
   24720: result <= 12'b010110010100;
   24721: result <= 12'b010110010011;
   24722: result <= 12'b010110010011;
   24723: result <= 12'b010110010011;
   24724: result <= 12'b010110010011;
   24725: result <= 12'b010110010011;
   24726: result <= 12'b010110010011;
   24727: result <= 12'b010110010011;
   24728: result <= 12'b010110010010;
   24729: result <= 12'b010110010010;
   24730: result <= 12'b010110010010;
   24731: result <= 12'b010110010010;
   24732: result <= 12'b010110010010;
   24733: result <= 12'b010110010010;
   24734: result <= 12'b010110010010;
   24735: result <= 12'b010110010001;
   24736: result <= 12'b010110010001;
   24737: result <= 12'b010110010001;
   24738: result <= 12'b010110010001;
   24739: result <= 12'b010110010001;
   24740: result <= 12'b010110010001;
   24741: result <= 12'b010110010001;
   24742: result <= 12'b010110010000;
   24743: result <= 12'b010110010000;
   24744: result <= 12'b010110010000;
   24745: result <= 12'b010110010000;
   24746: result <= 12'b010110010000;
   24747: result <= 12'b010110010000;
   24748: result <= 12'b010110010000;
   24749: result <= 12'b010110001111;
   24750: result <= 12'b010110001111;
   24751: result <= 12'b010110001111;
   24752: result <= 12'b010110001111;
   24753: result <= 12'b010110001111;
   24754: result <= 12'b010110001111;
   24755: result <= 12'b010110001111;
   24756: result <= 12'b010110001110;
   24757: result <= 12'b010110001110;
   24758: result <= 12'b010110001110;
   24759: result <= 12'b010110001110;
   24760: result <= 12'b010110001110;
   24761: result <= 12'b010110001110;
   24762: result <= 12'b010110001110;
   24763: result <= 12'b010110001101;
   24764: result <= 12'b010110001101;
   24765: result <= 12'b010110001101;
   24766: result <= 12'b010110001101;
   24767: result <= 12'b010110001101;
   24768: result <= 12'b010110001101;
   24769: result <= 12'b010110001101;
   24770: result <= 12'b010110001100;
   24771: result <= 12'b010110001100;
   24772: result <= 12'b010110001100;
   24773: result <= 12'b010110001100;
   24774: result <= 12'b010110001100;
   24775: result <= 12'b010110001100;
   24776: result <= 12'b010110001100;
   24777: result <= 12'b010110001011;
   24778: result <= 12'b010110001011;
   24779: result <= 12'b010110001011;
   24780: result <= 12'b010110001011;
   24781: result <= 12'b010110001011;
   24782: result <= 12'b010110001011;
   24783: result <= 12'b010110001011;
   24784: result <= 12'b010110001010;
   24785: result <= 12'b010110001010;
   24786: result <= 12'b010110001010;
   24787: result <= 12'b010110001010;
   24788: result <= 12'b010110001010;
   24789: result <= 12'b010110001010;
   24790: result <= 12'b010110001010;
   24791: result <= 12'b010110001001;
   24792: result <= 12'b010110001001;
   24793: result <= 12'b010110001001;
   24794: result <= 12'b010110001001;
   24795: result <= 12'b010110001001;
   24796: result <= 12'b010110001001;
   24797: result <= 12'b010110001001;
   24798: result <= 12'b010110001001;
   24799: result <= 12'b010110001000;
   24800: result <= 12'b010110001000;
   24801: result <= 12'b010110001000;
   24802: result <= 12'b010110001000;
   24803: result <= 12'b010110001000;
   24804: result <= 12'b010110001000;
   24805: result <= 12'b010110001000;
   24806: result <= 12'b010110000111;
   24807: result <= 12'b010110000111;
   24808: result <= 12'b010110000111;
   24809: result <= 12'b010110000111;
   24810: result <= 12'b010110000111;
   24811: result <= 12'b010110000111;
   24812: result <= 12'b010110000111;
   24813: result <= 12'b010110000110;
   24814: result <= 12'b010110000110;
   24815: result <= 12'b010110000110;
   24816: result <= 12'b010110000110;
   24817: result <= 12'b010110000110;
   24818: result <= 12'b010110000110;
   24819: result <= 12'b010110000110;
   24820: result <= 12'b010110000101;
   24821: result <= 12'b010110000101;
   24822: result <= 12'b010110000101;
   24823: result <= 12'b010110000101;
   24824: result <= 12'b010110000101;
   24825: result <= 12'b010110000101;
   24826: result <= 12'b010110000101;
   24827: result <= 12'b010110000100;
   24828: result <= 12'b010110000100;
   24829: result <= 12'b010110000100;
   24830: result <= 12'b010110000100;
   24831: result <= 12'b010110000100;
   24832: result <= 12'b010110000100;
   24833: result <= 12'b010110000100;
   24834: result <= 12'b010110000011;
   24835: result <= 12'b010110000011;
   24836: result <= 12'b010110000011;
   24837: result <= 12'b010110000011;
   24838: result <= 12'b010110000011;
   24839: result <= 12'b010110000011;
   24840: result <= 12'b010110000011;
   24841: result <= 12'b010110000010;
   24842: result <= 12'b010110000010;
   24843: result <= 12'b010110000010;
   24844: result <= 12'b010110000010;
   24845: result <= 12'b010110000010;
   24846: result <= 12'b010110000010;
   24847: result <= 12'b010110000010;
   24848: result <= 12'b010110000001;
   24849: result <= 12'b010110000001;
   24850: result <= 12'b010110000001;
   24851: result <= 12'b010110000001;
   24852: result <= 12'b010110000001;
   24853: result <= 12'b010110000001;
   24854: result <= 12'b010110000001;
   24855: result <= 12'b010110000000;
   24856: result <= 12'b010110000000;
   24857: result <= 12'b010110000000;
   24858: result <= 12'b010110000000;
   24859: result <= 12'b010110000000;
   24860: result <= 12'b010110000000;
   24861: result <= 12'b010110000000;
   24862: result <= 12'b010101111111;
   24863: result <= 12'b010101111111;
   24864: result <= 12'b010101111111;
   24865: result <= 12'b010101111111;
   24866: result <= 12'b010101111111;
   24867: result <= 12'b010101111111;
   24868: result <= 12'b010101111111;
   24869: result <= 12'b010101111110;
   24870: result <= 12'b010101111110;
   24871: result <= 12'b010101111110;
   24872: result <= 12'b010101111110;
   24873: result <= 12'b010101111110;
   24874: result <= 12'b010101111110;
   24875: result <= 12'b010101111110;
   24876: result <= 12'b010101111101;
   24877: result <= 12'b010101111101;
   24878: result <= 12'b010101111101;
   24879: result <= 12'b010101111101;
   24880: result <= 12'b010101111101;
   24881: result <= 12'b010101111101;
   24882: result <= 12'b010101111101;
   24883: result <= 12'b010101111100;
   24884: result <= 12'b010101111100;
   24885: result <= 12'b010101111100;
   24886: result <= 12'b010101111100;
   24887: result <= 12'b010101111100;
   24888: result <= 12'b010101111100;
   24889: result <= 12'b010101111100;
   24890: result <= 12'b010101111011;
   24891: result <= 12'b010101111011;
   24892: result <= 12'b010101111011;
   24893: result <= 12'b010101111011;
   24894: result <= 12'b010101111011;
   24895: result <= 12'b010101111011;
   24896: result <= 12'b010101111011;
   24897: result <= 12'b010101111010;
   24898: result <= 12'b010101111010;
   24899: result <= 12'b010101111010;
   24900: result <= 12'b010101111010;
   24901: result <= 12'b010101111010;
   24902: result <= 12'b010101111010;
   24903: result <= 12'b010101111010;
   24904: result <= 12'b010101111001;
   24905: result <= 12'b010101111001;
   24906: result <= 12'b010101111001;
   24907: result <= 12'b010101111001;
   24908: result <= 12'b010101111001;
   24909: result <= 12'b010101111001;
   24910: result <= 12'b010101111001;
   24911: result <= 12'b010101111000;
   24912: result <= 12'b010101111000;
   24913: result <= 12'b010101111000;
   24914: result <= 12'b010101111000;
   24915: result <= 12'b010101111000;
   24916: result <= 12'b010101111000;
   24917: result <= 12'b010101111000;
   24918: result <= 12'b010101110111;
   24919: result <= 12'b010101110111;
   24920: result <= 12'b010101110111;
   24921: result <= 12'b010101110111;
   24922: result <= 12'b010101110111;
   24923: result <= 12'b010101110111;
   24924: result <= 12'b010101110111;
   24925: result <= 12'b010101110110;
   24926: result <= 12'b010101110110;
   24927: result <= 12'b010101110110;
   24928: result <= 12'b010101110110;
   24929: result <= 12'b010101110110;
   24930: result <= 12'b010101110110;
   24931: result <= 12'b010101110110;
   24932: result <= 12'b010101110101;
   24933: result <= 12'b010101110101;
   24934: result <= 12'b010101110101;
   24935: result <= 12'b010101110101;
   24936: result <= 12'b010101110101;
   24937: result <= 12'b010101110101;
   24938: result <= 12'b010101110101;
   24939: result <= 12'b010101110100;
   24940: result <= 12'b010101110100;
   24941: result <= 12'b010101110100;
   24942: result <= 12'b010101110100;
   24943: result <= 12'b010101110100;
   24944: result <= 12'b010101110100;
   24945: result <= 12'b010101110100;
   24946: result <= 12'b010101110011;
   24947: result <= 12'b010101110011;
   24948: result <= 12'b010101110011;
   24949: result <= 12'b010101110011;
   24950: result <= 12'b010101110011;
   24951: result <= 12'b010101110011;
   24952: result <= 12'b010101110011;
   24953: result <= 12'b010101110010;
   24954: result <= 12'b010101110010;
   24955: result <= 12'b010101110010;
   24956: result <= 12'b010101110010;
   24957: result <= 12'b010101110010;
   24958: result <= 12'b010101110010;
   24959: result <= 12'b010101110010;
   24960: result <= 12'b010101110001;
   24961: result <= 12'b010101110001;
   24962: result <= 12'b010101110001;
   24963: result <= 12'b010101110001;
   24964: result <= 12'b010101110001;
   24965: result <= 12'b010101110001;
   24966: result <= 12'b010101110001;
   24967: result <= 12'b010101110000;
   24968: result <= 12'b010101110000;
   24969: result <= 12'b010101110000;
   24970: result <= 12'b010101110000;
   24971: result <= 12'b010101110000;
   24972: result <= 12'b010101110000;
   24973: result <= 12'b010101101111;
   24974: result <= 12'b010101101111;
   24975: result <= 12'b010101101111;
   24976: result <= 12'b010101101111;
   24977: result <= 12'b010101101111;
   24978: result <= 12'b010101101111;
   24979: result <= 12'b010101101111;
   24980: result <= 12'b010101101110;
   24981: result <= 12'b010101101110;
   24982: result <= 12'b010101101110;
   24983: result <= 12'b010101101110;
   24984: result <= 12'b010101101110;
   24985: result <= 12'b010101101110;
   24986: result <= 12'b010101101110;
   24987: result <= 12'b010101101101;
   24988: result <= 12'b010101101101;
   24989: result <= 12'b010101101101;
   24990: result <= 12'b010101101101;
   24991: result <= 12'b010101101101;
   24992: result <= 12'b010101101101;
   24993: result <= 12'b010101101101;
   24994: result <= 12'b010101101100;
   24995: result <= 12'b010101101100;
   24996: result <= 12'b010101101100;
   24997: result <= 12'b010101101100;
   24998: result <= 12'b010101101100;
   24999: result <= 12'b010101101100;
   25000: result <= 12'b010101101100;
   25001: result <= 12'b010101101011;
   25002: result <= 12'b010101101011;
   25003: result <= 12'b010101101011;
   25004: result <= 12'b010101101011;
   25005: result <= 12'b010101101011;
   25006: result <= 12'b010101101011;
   25007: result <= 12'b010101101011;
   25008: result <= 12'b010101101010;
   25009: result <= 12'b010101101010;
   25010: result <= 12'b010101101010;
   25011: result <= 12'b010101101010;
   25012: result <= 12'b010101101010;
   25013: result <= 12'b010101101010;
   25014: result <= 12'b010101101010;
   25015: result <= 12'b010101101001;
   25016: result <= 12'b010101101001;
   25017: result <= 12'b010101101001;
   25018: result <= 12'b010101101001;
   25019: result <= 12'b010101101001;
   25020: result <= 12'b010101101001;
   25021: result <= 12'b010101101001;
   25022: result <= 12'b010101101000;
   25023: result <= 12'b010101101000;
   25024: result <= 12'b010101101000;
   25025: result <= 12'b010101101000;
   25026: result <= 12'b010101101000;
   25027: result <= 12'b010101101000;
   25028: result <= 12'b010101101000;
   25029: result <= 12'b010101100111;
   25030: result <= 12'b010101100111;
   25031: result <= 12'b010101100111;
   25032: result <= 12'b010101100111;
   25033: result <= 12'b010101100111;
   25034: result <= 12'b010101100111;
   25035: result <= 12'b010101100111;
   25036: result <= 12'b010101100110;
   25037: result <= 12'b010101100110;
   25038: result <= 12'b010101100110;
   25039: result <= 12'b010101100110;
   25040: result <= 12'b010101100110;
   25041: result <= 12'b010101100110;
   25042: result <= 12'b010101100110;
   25043: result <= 12'b010101100101;
   25044: result <= 12'b010101100101;
   25045: result <= 12'b010101100101;
   25046: result <= 12'b010101100101;
   25047: result <= 12'b010101100101;
   25048: result <= 12'b010101100101;
   25049: result <= 12'b010101100101;
   25050: result <= 12'b010101100100;
   25051: result <= 12'b010101100100;
   25052: result <= 12'b010101100100;
   25053: result <= 12'b010101100100;
   25054: result <= 12'b010101100100;
   25055: result <= 12'b010101100100;
   25056: result <= 12'b010101100100;
   25057: result <= 12'b010101100011;
   25058: result <= 12'b010101100011;
   25059: result <= 12'b010101100011;
   25060: result <= 12'b010101100011;
   25061: result <= 12'b010101100011;
   25062: result <= 12'b010101100011;
   25063: result <= 12'b010101100010;
   25064: result <= 12'b010101100010;
   25065: result <= 12'b010101100010;
   25066: result <= 12'b010101100010;
   25067: result <= 12'b010101100010;
   25068: result <= 12'b010101100010;
   25069: result <= 12'b010101100010;
   25070: result <= 12'b010101100001;
   25071: result <= 12'b010101100001;
   25072: result <= 12'b010101100001;
   25073: result <= 12'b010101100001;
   25074: result <= 12'b010101100001;
   25075: result <= 12'b010101100001;
   25076: result <= 12'b010101100001;
   25077: result <= 12'b010101100000;
   25078: result <= 12'b010101100000;
   25079: result <= 12'b010101100000;
   25080: result <= 12'b010101100000;
   25081: result <= 12'b010101100000;
   25082: result <= 12'b010101100000;
   25083: result <= 12'b010101100000;
   25084: result <= 12'b010101011111;
   25085: result <= 12'b010101011111;
   25086: result <= 12'b010101011111;
   25087: result <= 12'b010101011111;
   25088: result <= 12'b010101011111;
   25089: result <= 12'b010101011111;
   25090: result <= 12'b010101011111;
   25091: result <= 12'b010101011110;
   25092: result <= 12'b010101011110;
   25093: result <= 12'b010101011110;
   25094: result <= 12'b010101011110;
   25095: result <= 12'b010101011110;
   25096: result <= 12'b010101011110;
   25097: result <= 12'b010101011110;
   25098: result <= 12'b010101011101;
   25099: result <= 12'b010101011101;
   25100: result <= 12'b010101011101;
   25101: result <= 12'b010101011101;
   25102: result <= 12'b010101011101;
   25103: result <= 12'b010101011101;
   25104: result <= 12'b010101011101;
   25105: result <= 12'b010101011100;
   25106: result <= 12'b010101011100;
   25107: result <= 12'b010101011100;
   25108: result <= 12'b010101011100;
   25109: result <= 12'b010101011100;
   25110: result <= 12'b010101011100;
   25111: result <= 12'b010101011100;
   25112: result <= 12'b010101011011;
   25113: result <= 12'b010101011011;
   25114: result <= 12'b010101011011;
   25115: result <= 12'b010101011011;
   25116: result <= 12'b010101011011;
   25117: result <= 12'b010101011011;
   25118: result <= 12'b010101011010;
   25119: result <= 12'b010101011010;
   25120: result <= 12'b010101011010;
   25121: result <= 12'b010101011010;
   25122: result <= 12'b010101011010;
   25123: result <= 12'b010101011010;
   25124: result <= 12'b010101011010;
   25125: result <= 12'b010101011001;
   25126: result <= 12'b010101011001;
   25127: result <= 12'b010101011001;
   25128: result <= 12'b010101011001;
   25129: result <= 12'b010101011001;
   25130: result <= 12'b010101011001;
   25131: result <= 12'b010101011001;
   25132: result <= 12'b010101011000;
   25133: result <= 12'b010101011000;
   25134: result <= 12'b010101011000;
   25135: result <= 12'b010101011000;
   25136: result <= 12'b010101011000;
   25137: result <= 12'b010101011000;
   25138: result <= 12'b010101011000;
   25139: result <= 12'b010101010111;
   25140: result <= 12'b010101010111;
   25141: result <= 12'b010101010111;
   25142: result <= 12'b010101010111;
   25143: result <= 12'b010101010111;
   25144: result <= 12'b010101010111;
   25145: result <= 12'b010101010111;
   25146: result <= 12'b010101010110;
   25147: result <= 12'b010101010110;
   25148: result <= 12'b010101010110;
   25149: result <= 12'b010101010110;
   25150: result <= 12'b010101010110;
   25151: result <= 12'b010101010110;
   25152: result <= 12'b010101010110;
   25153: result <= 12'b010101010101;
   25154: result <= 12'b010101010101;
   25155: result <= 12'b010101010101;
   25156: result <= 12'b010101010101;
   25157: result <= 12'b010101010101;
   25158: result <= 12'b010101010101;
   25159: result <= 12'b010101010100;
   25160: result <= 12'b010101010100;
   25161: result <= 12'b010101010100;
   25162: result <= 12'b010101010100;
   25163: result <= 12'b010101010100;
   25164: result <= 12'b010101010100;
   25165: result <= 12'b010101010100;
   25166: result <= 12'b010101010011;
   25167: result <= 12'b010101010011;
   25168: result <= 12'b010101010011;
   25169: result <= 12'b010101010011;
   25170: result <= 12'b010101010011;
   25171: result <= 12'b010101010011;
   25172: result <= 12'b010101010011;
   25173: result <= 12'b010101010010;
   25174: result <= 12'b010101010010;
   25175: result <= 12'b010101010010;
   25176: result <= 12'b010101010010;
   25177: result <= 12'b010101010010;
   25178: result <= 12'b010101010010;
   25179: result <= 12'b010101010010;
   25180: result <= 12'b010101010001;
   25181: result <= 12'b010101010001;
   25182: result <= 12'b010101010001;
   25183: result <= 12'b010101010001;
   25184: result <= 12'b010101010001;
   25185: result <= 12'b010101010001;
   25186: result <= 12'b010101010001;
   25187: result <= 12'b010101010000;
   25188: result <= 12'b010101010000;
   25189: result <= 12'b010101010000;
   25190: result <= 12'b010101010000;
   25191: result <= 12'b010101010000;
   25192: result <= 12'b010101010000;
   25193: result <= 12'b010101010000;
   25194: result <= 12'b010101001111;
   25195: result <= 12'b010101001111;
   25196: result <= 12'b010101001111;
   25197: result <= 12'b010101001111;
   25198: result <= 12'b010101001111;
   25199: result <= 12'b010101001111;
   25200: result <= 12'b010101001110;
   25201: result <= 12'b010101001110;
   25202: result <= 12'b010101001110;
   25203: result <= 12'b010101001110;
   25204: result <= 12'b010101001110;
   25205: result <= 12'b010101001110;
   25206: result <= 12'b010101001110;
   25207: result <= 12'b010101001101;
   25208: result <= 12'b010101001101;
   25209: result <= 12'b010101001101;
   25210: result <= 12'b010101001101;
   25211: result <= 12'b010101001101;
   25212: result <= 12'b010101001101;
   25213: result <= 12'b010101001101;
   25214: result <= 12'b010101001100;
   25215: result <= 12'b010101001100;
   25216: result <= 12'b010101001100;
   25217: result <= 12'b010101001100;
   25218: result <= 12'b010101001100;
   25219: result <= 12'b010101001100;
   25220: result <= 12'b010101001100;
   25221: result <= 12'b010101001011;
   25222: result <= 12'b010101001011;
   25223: result <= 12'b010101001011;
   25224: result <= 12'b010101001011;
   25225: result <= 12'b010101001011;
   25226: result <= 12'b010101001011;
   25227: result <= 12'b010101001011;
   25228: result <= 12'b010101001010;
   25229: result <= 12'b010101001010;
   25230: result <= 12'b010101001010;
   25231: result <= 12'b010101001010;
   25232: result <= 12'b010101001010;
   25233: result <= 12'b010101001010;
   25234: result <= 12'b010101001001;
   25235: result <= 12'b010101001001;
   25236: result <= 12'b010101001001;
   25237: result <= 12'b010101001001;
   25238: result <= 12'b010101001001;
   25239: result <= 12'b010101001001;
   25240: result <= 12'b010101001001;
   25241: result <= 12'b010101001000;
   25242: result <= 12'b010101001000;
   25243: result <= 12'b010101001000;
   25244: result <= 12'b010101001000;
   25245: result <= 12'b010101001000;
   25246: result <= 12'b010101001000;
   25247: result <= 12'b010101001000;
   25248: result <= 12'b010101000111;
   25249: result <= 12'b010101000111;
   25250: result <= 12'b010101000111;
   25251: result <= 12'b010101000111;
   25252: result <= 12'b010101000111;
   25253: result <= 12'b010101000111;
   25254: result <= 12'b010101000111;
   25255: result <= 12'b010101000110;
   25256: result <= 12'b010101000110;
   25257: result <= 12'b010101000110;
   25258: result <= 12'b010101000110;
   25259: result <= 12'b010101000110;
   25260: result <= 12'b010101000110;
   25261: result <= 12'b010101000101;
   25262: result <= 12'b010101000101;
   25263: result <= 12'b010101000101;
   25264: result <= 12'b010101000101;
   25265: result <= 12'b010101000101;
   25266: result <= 12'b010101000101;
   25267: result <= 12'b010101000101;
   25268: result <= 12'b010101000100;
   25269: result <= 12'b010101000100;
   25270: result <= 12'b010101000100;
   25271: result <= 12'b010101000100;
   25272: result <= 12'b010101000100;
   25273: result <= 12'b010101000100;
   25274: result <= 12'b010101000100;
   25275: result <= 12'b010101000011;
   25276: result <= 12'b010101000011;
   25277: result <= 12'b010101000011;
   25278: result <= 12'b010101000011;
   25279: result <= 12'b010101000011;
   25280: result <= 12'b010101000011;
   25281: result <= 12'b010101000011;
   25282: result <= 12'b010101000010;
   25283: result <= 12'b010101000010;
   25284: result <= 12'b010101000010;
   25285: result <= 12'b010101000010;
   25286: result <= 12'b010101000010;
   25287: result <= 12'b010101000010;
   25288: result <= 12'b010101000010;
   25289: result <= 12'b010101000001;
   25290: result <= 12'b010101000001;
   25291: result <= 12'b010101000001;
   25292: result <= 12'b010101000001;
   25293: result <= 12'b010101000001;
   25294: result <= 12'b010101000001;
   25295: result <= 12'b010101000000;
   25296: result <= 12'b010101000000;
   25297: result <= 12'b010101000000;
   25298: result <= 12'b010101000000;
   25299: result <= 12'b010101000000;
   25300: result <= 12'b010101000000;
   25301: result <= 12'b010101000000;
   25302: result <= 12'b010100111111;
   25303: result <= 12'b010100111111;
   25304: result <= 12'b010100111111;
   25305: result <= 12'b010100111111;
   25306: result <= 12'b010100111111;
   25307: result <= 12'b010100111111;
   25308: result <= 12'b010100111111;
   25309: result <= 12'b010100111110;
   25310: result <= 12'b010100111110;
   25311: result <= 12'b010100111110;
   25312: result <= 12'b010100111110;
   25313: result <= 12'b010100111110;
   25314: result <= 12'b010100111110;
   25315: result <= 12'b010100111110;
   25316: result <= 12'b010100111101;
   25317: result <= 12'b010100111101;
   25318: result <= 12'b010100111101;
   25319: result <= 12'b010100111101;
   25320: result <= 12'b010100111101;
   25321: result <= 12'b010100111101;
   25322: result <= 12'b010100111100;
   25323: result <= 12'b010100111100;
   25324: result <= 12'b010100111100;
   25325: result <= 12'b010100111100;
   25326: result <= 12'b010100111100;
   25327: result <= 12'b010100111100;
   25328: result <= 12'b010100111100;
   25329: result <= 12'b010100111011;
   25330: result <= 12'b010100111011;
   25331: result <= 12'b010100111011;
   25332: result <= 12'b010100111011;
   25333: result <= 12'b010100111011;
   25334: result <= 12'b010100111011;
   25335: result <= 12'b010100111011;
   25336: result <= 12'b010100111010;
   25337: result <= 12'b010100111010;
   25338: result <= 12'b010100111010;
   25339: result <= 12'b010100111010;
   25340: result <= 12'b010100111010;
   25341: result <= 12'b010100111010;
   25342: result <= 12'b010100111001;
   25343: result <= 12'b010100111001;
   25344: result <= 12'b010100111001;
   25345: result <= 12'b010100111001;
   25346: result <= 12'b010100111001;
   25347: result <= 12'b010100111001;
   25348: result <= 12'b010100111001;
   25349: result <= 12'b010100111000;
   25350: result <= 12'b010100111000;
   25351: result <= 12'b010100111000;
   25352: result <= 12'b010100111000;
   25353: result <= 12'b010100111000;
   25354: result <= 12'b010100111000;
   25355: result <= 12'b010100111000;
   25356: result <= 12'b010100110111;
   25357: result <= 12'b010100110111;
   25358: result <= 12'b010100110111;
   25359: result <= 12'b010100110111;
   25360: result <= 12'b010100110111;
   25361: result <= 12'b010100110111;
   25362: result <= 12'b010100110111;
   25363: result <= 12'b010100110110;
   25364: result <= 12'b010100110110;
   25365: result <= 12'b010100110110;
   25366: result <= 12'b010100110110;
   25367: result <= 12'b010100110110;
   25368: result <= 12'b010100110110;
   25369: result <= 12'b010100110101;
   25370: result <= 12'b010100110101;
   25371: result <= 12'b010100110101;
   25372: result <= 12'b010100110101;
   25373: result <= 12'b010100110101;
   25374: result <= 12'b010100110101;
   25375: result <= 12'b010100110101;
   25376: result <= 12'b010100110100;
   25377: result <= 12'b010100110100;
   25378: result <= 12'b010100110100;
   25379: result <= 12'b010100110100;
   25380: result <= 12'b010100110100;
   25381: result <= 12'b010100110100;
   25382: result <= 12'b010100110100;
   25383: result <= 12'b010100110011;
   25384: result <= 12'b010100110011;
   25385: result <= 12'b010100110011;
   25386: result <= 12'b010100110011;
   25387: result <= 12'b010100110011;
   25388: result <= 12'b010100110011;
   25389: result <= 12'b010100110010;
   25390: result <= 12'b010100110010;
   25391: result <= 12'b010100110010;
   25392: result <= 12'b010100110010;
   25393: result <= 12'b010100110010;
   25394: result <= 12'b010100110010;
   25395: result <= 12'b010100110010;
   25396: result <= 12'b010100110001;
   25397: result <= 12'b010100110001;
   25398: result <= 12'b010100110001;
   25399: result <= 12'b010100110001;
   25400: result <= 12'b010100110001;
   25401: result <= 12'b010100110001;
   25402: result <= 12'b010100110001;
   25403: result <= 12'b010100110000;
   25404: result <= 12'b010100110000;
   25405: result <= 12'b010100110000;
   25406: result <= 12'b010100110000;
   25407: result <= 12'b010100110000;
   25408: result <= 12'b010100110000;
   25409: result <= 12'b010100110000;
   25410: result <= 12'b010100101111;
   25411: result <= 12'b010100101111;
   25412: result <= 12'b010100101111;
   25413: result <= 12'b010100101111;
   25414: result <= 12'b010100101111;
   25415: result <= 12'b010100101111;
   25416: result <= 12'b010100101110;
   25417: result <= 12'b010100101110;
   25418: result <= 12'b010100101110;
   25419: result <= 12'b010100101110;
   25420: result <= 12'b010100101110;
   25421: result <= 12'b010100101110;
   25422: result <= 12'b010100101110;
   25423: result <= 12'b010100101101;
   25424: result <= 12'b010100101101;
   25425: result <= 12'b010100101101;
   25426: result <= 12'b010100101101;
   25427: result <= 12'b010100101101;
   25428: result <= 12'b010100101101;
   25429: result <= 12'b010100101101;
   25430: result <= 12'b010100101100;
   25431: result <= 12'b010100101100;
   25432: result <= 12'b010100101100;
   25433: result <= 12'b010100101100;
   25434: result <= 12'b010100101100;
   25435: result <= 12'b010100101100;
   25436: result <= 12'b010100101011;
   25437: result <= 12'b010100101011;
   25438: result <= 12'b010100101011;
   25439: result <= 12'b010100101011;
   25440: result <= 12'b010100101011;
   25441: result <= 12'b010100101011;
   25442: result <= 12'b010100101011;
   25443: result <= 12'b010100101010;
   25444: result <= 12'b010100101010;
   25445: result <= 12'b010100101010;
   25446: result <= 12'b010100101010;
   25447: result <= 12'b010100101010;
   25448: result <= 12'b010100101010;
   25449: result <= 12'b010100101010;
   25450: result <= 12'b010100101001;
   25451: result <= 12'b010100101001;
   25452: result <= 12'b010100101001;
   25453: result <= 12'b010100101001;
   25454: result <= 12'b010100101001;
   25455: result <= 12'b010100101001;
   25456: result <= 12'b010100101000;
   25457: result <= 12'b010100101000;
   25458: result <= 12'b010100101000;
   25459: result <= 12'b010100101000;
   25460: result <= 12'b010100101000;
   25461: result <= 12'b010100101000;
   25462: result <= 12'b010100101000;
   25463: result <= 12'b010100100111;
   25464: result <= 12'b010100100111;
   25465: result <= 12'b010100100111;
   25466: result <= 12'b010100100111;
   25467: result <= 12'b010100100111;
   25468: result <= 12'b010100100111;
   25469: result <= 12'b010100100111;
   25470: result <= 12'b010100100110;
   25471: result <= 12'b010100100110;
   25472: result <= 12'b010100100110;
   25473: result <= 12'b010100100110;
   25474: result <= 12'b010100100110;
   25475: result <= 12'b010100100110;
   25476: result <= 12'b010100100101;
   25477: result <= 12'b010100100101;
   25478: result <= 12'b010100100101;
   25479: result <= 12'b010100100101;
   25480: result <= 12'b010100100101;
   25481: result <= 12'b010100100101;
   25482: result <= 12'b010100100101;
   25483: result <= 12'b010100100100;
   25484: result <= 12'b010100100100;
   25485: result <= 12'b010100100100;
   25486: result <= 12'b010100100100;
   25487: result <= 12'b010100100100;
   25488: result <= 12'b010100100100;
   25489: result <= 12'b010100100100;
   25490: result <= 12'b010100100011;
   25491: result <= 12'b010100100011;
   25492: result <= 12'b010100100011;
   25493: result <= 12'b010100100011;
   25494: result <= 12'b010100100011;
   25495: result <= 12'b010100100011;
   25496: result <= 12'b010100100010;
   25497: result <= 12'b010100100010;
   25498: result <= 12'b010100100010;
   25499: result <= 12'b010100100010;
   25500: result <= 12'b010100100010;
   25501: result <= 12'b010100100010;
   25502: result <= 12'b010100100010;
   25503: result <= 12'b010100100001;
   25504: result <= 12'b010100100001;
   25505: result <= 12'b010100100001;
   25506: result <= 12'b010100100001;
   25507: result <= 12'b010100100001;
   25508: result <= 12'b010100100001;
   25509: result <= 12'b010100100000;
   25510: result <= 12'b010100100000;
   25511: result <= 12'b010100100000;
   25512: result <= 12'b010100100000;
   25513: result <= 12'b010100100000;
   25514: result <= 12'b010100100000;
   25515: result <= 12'b010100100000;
   25516: result <= 12'b010100011111;
   25517: result <= 12'b010100011111;
   25518: result <= 12'b010100011111;
   25519: result <= 12'b010100011111;
   25520: result <= 12'b010100011111;
   25521: result <= 12'b010100011111;
   25522: result <= 12'b010100011111;
   25523: result <= 12'b010100011110;
   25524: result <= 12'b010100011110;
   25525: result <= 12'b010100011110;
   25526: result <= 12'b010100011110;
   25527: result <= 12'b010100011110;
   25528: result <= 12'b010100011110;
   25529: result <= 12'b010100011101;
   25530: result <= 12'b010100011101;
   25531: result <= 12'b010100011101;
   25532: result <= 12'b010100011101;
   25533: result <= 12'b010100011101;
   25534: result <= 12'b010100011101;
   25535: result <= 12'b010100011101;
   25536: result <= 12'b010100011100;
   25537: result <= 12'b010100011100;
   25538: result <= 12'b010100011100;
   25539: result <= 12'b010100011100;
   25540: result <= 12'b010100011100;
   25541: result <= 12'b010100011100;
   25542: result <= 12'b010100011100;
   25543: result <= 12'b010100011011;
   25544: result <= 12'b010100011011;
   25545: result <= 12'b010100011011;
   25546: result <= 12'b010100011011;
   25547: result <= 12'b010100011011;
   25548: result <= 12'b010100011011;
   25549: result <= 12'b010100011010;
   25550: result <= 12'b010100011010;
   25551: result <= 12'b010100011010;
   25552: result <= 12'b010100011010;
   25553: result <= 12'b010100011010;
   25554: result <= 12'b010100011010;
   25555: result <= 12'b010100011010;
   25556: result <= 12'b010100011001;
   25557: result <= 12'b010100011001;
   25558: result <= 12'b010100011001;
   25559: result <= 12'b010100011001;
   25560: result <= 12'b010100011001;
   25561: result <= 12'b010100011001;
   25562: result <= 12'b010100011000;
   25563: result <= 12'b010100011000;
   25564: result <= 12'b010100011000;
   25565: result <= 12'b010100011000;
   25566: result <= 12'b010100011000;
   25567: result <= 12'b010100011000;
   25568: result <= 12'b010100011000;
   25569: result <= 12'b010100010111;
   25570: result <= 12'b010100010111;
   25571: result <= 12'b010100010111;
   25572: result <= 12'b010100010111;
   25573: result <= 12'b010100010111;
   25574: result <= 12'b010100010111;
   25575: result <= 12'b010100010111;
   25576: result <= 12'b010100010110;
   25577: result <= 12'b010100010110;
   25578: result <= 12'b010100010110;
   25579: result <= 12'b010100010110;
   25580: result <= 12'b010100010110;
   25581: result <= 12'b010100010110;
   25582: result <= 12'b010100010101;
   25583: result <= 12'b010100010101;
   25584: result <= 12'b010100010101;
   25585: result <= 12'b010100010101;
   25586: result <= 12'b010100010101;
   25587: result <= 12'b010100010101;
   25588: result <= 12'b010100010101;
   25589: result <= 12'b010100010100;
   25590: result <= 12'b010100010100;
   25591: result <= 12'b010100010100;
   25592: result <= 12'b010100010100;
   25593: result <= 12'b010100010100;
   25594: result <= 12'b010100010100;
   25595: result <= 12'b010100010011;
   25596: result <= 12'b010100010011;
   25597: result <= 12'b010100010011;
   25598: result <= 12'b010100010011;
   25599: result <= 12'b010100010011;
   25600: result <= 12'b010100010011;
   25601: result <= 12'b010100010011;
   25602: result <= 12'b010100010010;
   25603: result <= 12'b010100010010;
   25604: result <= 12'b010100010010;
   25605: result <= 12'b010100010010;
   25606: result <= 12'b010100010010;
   25607: result <= 12'b010100010010;
   25608: result <= 12'b010100010010;
   25609: result <= 12'b010100010001;
   25610: result <= 12'b010100010001;
   25611: result <= 12'b010100010001;
   25612: result <= 12'b010100010001;
   25613: result <= 12'b010100010001;
   25614: result <= 12'b010100010001;
   25615: result <= 12'b010100010000;
   25616: result <= 12'b010100010000;
   25617: result <= 12'b010100010000;
   25618: result <= 12'b010100010000;
   25619: result <= 12'b010100010000;
   25620: result <= 12'b010100010000;
   25621: result <= 12'b010100010000;
   25622: result <= 12'b010100001111;
   25623: result <= 12'b010100001111;
   25624: result <= 12'b010100001111;
   25625: result <= 12'b010100001111;
   25626: result <= 12'b010100001111;
   25627: result <= 12'b010100001111;
   25628: result <= 12'b010100001110;
   25629: result <= 12'b010100001110;
   25630: result <= 12'b010100001110;
   25631: result <= 12'b010100001110;
   25632: result <= 12'b010100001110;
   25633: result <= 12'b010100001110;
   25634: result <= 12'b010100001110;
   25635: result <= 12'b010100001101;
   25636: result <= 12'b010100001101;
   25637: result <= 12'b010100001101;
   25638: result <= 12'b010100001101;
   25639: result <= 12'b010100001101;
   25640: result <= 12'b010100001101;
   25641: result <= 12'b010100001101;
   25642: result <= 12'b010100001100;
   25643: result <= 12'b010100001100;
   25644: result <= 12'b010100001100;
   25645: result <= 12'b010100001100;
   25646: result <= 12'b010100001100;
   25647: result <= 12'b010100001100;
   25648: result <= 12'b010100001011;
   25649: result <= 12'b010100001011;
   25650: result <= 12'b010100001011;
   25651: result <= 12'b010100001011;
   25652: result <= 12'b010100001011;
   25653: result <= 12'b010100001011;
   25654: result <= 12'b010100001011;
   25655: result <= 12'b010100001010;
   25656: result <= 12'b010100001010;
   25657: result <= 12'b010100001010;
   25658: result <= 12'b010100001010;
   25659: result <= 12'b010100001010;
   25660: result <= 12'b010100001010;
   25661: result <= 12'b010100001001;
   25662: result <= 12'b010100001001;
   25663: result <= 12'b010100001001;
   25664: result <= 12'b010100001001;
   25665: result <= 12'b010100001001;
   25666: result <= 12'b010100001001;
   25667: result <= 12'b010100001001;
   25668: result <= 12'b010100001000;
   25669: result <= 12'b010100001000;
   25670: result <= 12'b010100001000;
   25671: result <= 12'b010100001000;
   25672: result <= 12'b010100001000;
   25673: result <= 12'b010100001000;
   25674: result <= 12'b010100000111;
   25675: result <= 12'b010100000111;
   25676: result <= 12'b010100000111;
   25677: result <= 12'b010100000111;
   25678: result <= 12'b010100000111;
   25679: result <= 12'b010100000111;
   25680: result <= 12'b010100000111;
   25681: result <= 12'b010100000110;
   25682: result <= 12'b010100000110;
   25683: result <= 12'b010100000110;
   25684: result <= 12'b010100000110;
   25685: result <= 12'b010100000110;
   25686: result <= 12'b010100000110;
   25687: result <= 12'b010100000101;
   25688: result <= 12'b010100000101;
   25689: result <= 12'b010100000101;
   25690: result <= 12'b010100000101;
   25691: result <= 12'b010100000101;
   25692: result <= 12'b010100000101;
   25693: result <= 12'b010100000101;
   25694: result <= 12'b010100000100;
   25695: result <= 12'b010100000100;
   25696: result <= 12'b010100000100;
   25697: result <= 12'b010100000100;
   25698: result <= 12'b010100000100;
   25699: result <= 12'b010100000100;
   25700: result <= 12'b010100000011;
   25701: result <= 12'b010100000011;
   25702: result <= 12'b010100000011;
   25703: result <= 12'b010100000011;
   25704: result <= 12'b010100000011;
   25705: result <= 12'b010100000011;
   25706: result <= 12'b010100000011;
   25707: result <= 12'b010100000010;
   25708: result <= 12'b010100000010;
   25709: result <= 12'b010100000010;
   25710: result <= 12'b010100000010;
   25711: result <= 12'b010100000010;
   25712: result <= 12'b010100000010;
   25713: result <= 12'b010100000010;
   25714: result <= 12'b010100000001;
   25715: result <= 12'b010100000001;
   25716: result <= 12'b010100000001;
   25717: result <= 12'b010100000001;
   25718: result <= 12'b010100000001;
   25719: result <= 12'b010100000001;
   25720: result <= 12'b010100000000;
   25721: result <= 12'b010100000000;
   25722: result <= 12'b010100000000;
   25723: result <= 12'b010100000000;
   25724: result <= 12'b010100000000;
   25725: result <= 12'b010100000000;
   25726: result <= 12'b010100000000;
   25727: result <= 12'b010011111111;
   25728: result <= 12'b010011111111;
   25729: result <= 12'b010011111111;
   25730: result <= 12'b010011111111;
   25731: result <= 12'b010011111111;
   25732: result <= 12'b010011111111;
   25733: result <= 12'b010011111110;
   25734: result <= 12'b010011111110;
   25735: result <= 12'b010011111110;
   25736: result <= 12'b010011111110;
   25737: result <= 12'b010011111110;
   25738: result <= 12'b010011111110;
   25739: result <= 12'b010011111110;
   25740: result <= 12'b010011111101;
   25741: result <= 12'b010011111101;
   25742: result <= 12'b010011111101;
   25743: result <= 12'b010011111101;
   25744: result <= 12'b010011111101;
   25745: result <= 12'b010011111101;
   25746: result <= 12'b010011111100;
   25747: result <= 12'b010011111100;
   25748: result <= 12'b010011111100;
   25749: result <= 12'b010011111100;
   25750: result <= 12'b010011111100;
   25751: result <= 12'b010011111100;
   25752: result <= 12'b010011111100;
   25753: result <= 12'b010011111011;
   25754: result <= 12'b010011111011;
   25755: result <= 12'b010011111011;
   25756: result <= 12'b010011111011;
   25757: result <= 12'b010011111011;
   25758: result <= 12'b010011111011;
   25759: result <= 12'b010011111010;
   25760: result <= 12'b010011111010;
   25761: result <= 12'b010011111010;
   25762: result <= 12'b010011111010;
   25763: result <= 12'b010011111010;
   25764: result <= 12'b010011111010;
   25765: result <= 12'b010011111010;
   25766: result <= 12'b010011111001;
   25767: result <= 12'b010011111001;
   25768: result <= 12'b010011111001;
   25769: result <= 12'b010011111001;
   25770: result <= 12'b010011111001;
   25771: result <= 12'b010011111001;
   25772: result <= 12'b010011111000;
   25773: result <= 12'b010011111000;
   25774: result <= 12'b010011111000;
   25775: result <= 12'b010011111000;
   25776: result <= 12'b010011111000;
   25777: result <= 12'b010011111000;
   25778: result <= 12'b010011111000;
   25779: result <= 12'b010011110111;
   25780: result <= 12'b010011110111;
   25781: result <= 12'b010011110111;
   25782: result <= 12'b010011110111;
   25783: result <= 12'b010011110111;
   25784: result <= 12'b010011110111;
   25785: result <= 12'b010011110110;
   25786: result <= 12'b010011110110;
   25787: result <= 12'b010011110110;
   25788: result <= 12'b010011110110;
   25789: result <= 12'b010011110110;
   25790: result <= 12'b010011110110;
   25791: result <= 12'b010011110110;
   25792: result <= 12'b010011110101;
   25793: result <= 12'b010011110101;
   25794: result <= 12'b010011110101;
   25795: result <= 12'b010011110101;
   25796: result <= 12'b010011110101;
   25797: result <= 12'b010011110101;
   25798: result <= 12'b010011110100;
   25799: result <= 12'b010011110100;
   25800: result <= 12'b010011110100;
   25801: result <= 12'b010011110100;
   25802: result <= 12'b010011110100;
   25803: result <= 12'b010011110100;
   25804: result <= 12'b010011110100;
   25805: result <= 12'b010011110011;
   25806: result <= 12'b010011110011;
   25807: result <= 12'b010011110011;
   25808: result <= 12'b010011110011;
   25809: result <= 12'b010011110011;
   25810: result <= 12'b010011110011;
   25811: result <= 12'b010011110010;
   25812: result <= 12'b010011110010;
   25813: result <= 12'b010011110010;
   25814: result <= 12'b010011110010;
   25815: result <= 12'b010011110010;
   25816: result <= 12'b010011110010;
   25817: result <= 12'b010011110010;
   25818: result <= 12'b010011110001;
   25819: result <= 12'b010011110001;
   25820: result <= 12'b010011110001;
   25821: result <= 12'b010011110001;
   25822: result <= 12'b010011110001;
   25823: result <= 12'b010011110001;
   25824: result <= 12'b010011110000;
   25825: result <= 12'b010011110000;
   25826: result <= 12'b010011110000;
   25827: result <= 12'b010011110000;
   25828: result <= 12'b010011110000;
   25829: result <= 12'b010011110000;
   25830: result <= 12'b010011110000;
   25831: result <= 12'b010011101111;
   25832: result <= 12'b010011101111;
   25833: result <= 12'b010011101111;
   25834: result <= 12'b010011101111;
   25835: result <= 12'b010011101111;
   25836: result <= 12'b010011101111;
   25837: result <= 12'b010011101110;
   25838: result <= 12'b010011101110;
   25839: result <= 12'b010011101110;
   25840: result <= 12'b010011101110;
   25841: result <= 12'b010011101110;
   25842: result <= 12'b010011101110;
   25843: result <= 12'b010011101110;
   25844: result <= 12'b010011101101;
   25845: result <= 12'b010011101101;
   25846: result <= 12'b010011101101;
   25847: result <= 12'b010011101101;
   25848: result <= 12'b010011101101;
   25849: result <= 12'b010011101101;
   25850: result <= 12'b010011101100;
   25851: result <= 12'b010011101100;
   25852: result <= 12'b010011101100;
   25853: result <= 12'b010011101100;
   25854: result <= 12'b010011101100;
   25855: result <= 12'b010011101100;
   25856: result <= 12'b010011101011;
   25857: result <= 12'b010011101011;
   25858: result <= 12'b010011101011;
   25859: result <= 12'b010011101011;
   25860: result <= 12'b010011101011;
   25861: result <= 12'b010011101011;
   25862: result <= 12'b010011101011;
   25863: result <= 12'b010011101010;
   25864: result <= 12'b010011101010;
   25865: result <= 12'b010011101010;
   25866: result <= 12'b010011101010;
   25867: result <= 12'b010011101010;
   25868: result <= 12'b010011101010;
   25869: result <= 12'b010011101001;
   25870: result <= 12'b010011101001;
   25871: result <= 12'b010011101001;
   25872: result <= 12'b010011101001;
   25873: result <= 12'b010011101001;
   25874: result <= 12'b010011101001;
   25875: result <= 12'b010011101001;
   25876: result <= 12'b010011101000;
   25877: result <= 12'b010011101000;
   25878: result <= 12'b010011101000;
   25879: result <= 12'b010011101000;
   25880: result <= 12'b010011101000;
   25881: result <= 12'b010011101000;
   25882: result <= 12'b010011100111;
   25883: result <= 12'b010011100111;
   25884: result <= 12'b010011100111;
   25885: result <= 12'b010011100111;
   25886: result <= 12'b010011100111;
   25887: result <= 12'b010011100111;
   25888: result <= 12'b010011100111;
   25889: result <= 12'b010011100110;
   25890: result <= 12'b010011100110;
   25891: result <= 12'b010011100110;
   25892: result <= 12'b010011100110;
   25893: result <= 12'b010011100110;
   25894: result <= 12'b010011100110;
   25895: result <= 12'b010011100101;
   25896: result <= 12'b010011100101;
   25897: result <= 12'b010011100101;
   25898: result <= 12'b010011100101;
   25899: result <= 12'b010011100101;
   25900: result <= 12'b010011100101;
   25901: result <= 12'b010011100101;
   25902: result <= 12'b010011100100;
   25903: result <= 12'b010011100100;
   25904: result <= 12'b010011100100;
   25905: result <= 12'b010011100100;
   25906: result <= 12'b010011100100;
   25907: result <= 12'b010011100100;
   25908: result <= 12'b010011100011;
   25909: result <= 12'b010011100011;
   25910: result <= 12'b010011100011;
   25911: result <= 12'b010011100011;
   25912: result <= 12'b010011100011;
   25913: result <= 12'b010011100011;
   25914: result <= 12'b010011100010;
   25915: result <= 12'b010011100010;
   25916: result <= 12'b010011100010;
   25917: result <= 12'b010011100010;
   25918: result <= 12'b010011100010;
   25919: result <= 12'b010011100010;
   25920: result <= 12'b010011100010;
   25921: result <= 12'b010011100001;
   25922: result <= 12'b010011100001;
   25923: result <= 12'b010011100001;
   25924: result <= 12'b010011100001;
   25925: result <= 12'b010011100001;
   25926: result <= 12'b010011100001;
   25927: result <= 12'b010011100000;
   25928: result <= 12'b010011100000;
   25929: result <= 12'b010011100000;
   25930: result <= 12'b010011100000;
   25931: result <= 12'b010011100000;
   25932: result <= 12'b010011100000;
   25933: result <= 12'b010011100000;
   25934: result <= 12'b010011011111;
   25935: result <= 12'b010011011111;
   25936: result <= 12'b010011011111;
   25937: result <= 12'b010011011111;
   25938: result <= 12'b010011011111;
   25939: result <= 12'b010011011111;
   25940: result <= 12'b010011011110;
   25941: result <= 12'b010011011110;
   25942: result <= 12'b010011011110;
   25943: result <= 12'b010011011110;
   25944: result <= 12'b010011011110;
   25945: result <= 12'b010011011110;
   25946: result <= 12'b010011011110;
   25947: result <= 12'b010011011101;
   25948: result <= 12'b010011011101;
   25949: result <= 12'b010011011101;
   25950: result <= 12'b010011011101;
   25951: result <= 12'b010011011101;
   25952: result <= 12'b010011011101;
   25953: result <= 12'b010011011100;
   25954: result <= 12'b010011011100;
   25955: result <= 12'b010011011100;
   25956: result <= 12'b010011011100;
   25957: result <= 12'b010011011100;
   25958: result <= 12'b010011011100;
   25959: result <= 12'b010011011011;
   25960: result <= 12'b010011011011;
   25961: result <= 12'b010011011011;
   25962: result <= 12'b010011011011;
   25963: result <= 12'b010011011011;
   25964: result <= 12'b010011011011;
   25965: result <= 12'b010011011011;
   25966: result <= 12'b010011011010;
   25967: result <= 12'b010011011010;
   25968: result <= 12'b010011011010;
   25969: result <= 12'b010011011010;
   25970: result <= 12'b010011011010;
   25971: result <= 12'b010011011010;
   25972: result <= 12'b010011011001;
   25973: result <= 12'b010011011001;
   25974: result <= 12'b010011011001;
   25975: result <= 12'b010011011001;
   25976: result <= 12'b010011011001;
   25977: result <= 12'b010011011001;
   25978: result <= 12'b010011011001;
   25979: result <= 12'b010011011000;
   25980: result <= 12'b010011011000;
   25981: result <= 12'b010011011000;
   25982: result <= 12'b010011011000;
   25983: result <= 12'b010011011000;
   25984: result <= 12'b010011011000;
   25985: result <= 12'b010011010111;
   25986: result <= 12'b010011010111;
   25987: result <= 12'b010011010111;
   25988: result <= 12'b010011010111;
   25989: result <= 12'b010011010111;
   25990: result <= 12'b010011010111;
   25991: result <= 12'b010011010110;
   25992: result <= 12'b010011010110;
   25993: result <= 12'b010011010110;
   25994: result <= 12'b010011010110;
   25995: result <= 12'b010011010110;
   25996: result <= 12'b010011010110;
   25997: result <= 12'b010011010110;
   25998: result <= 12'b010011010101;
   25999: result <= 12'b010011010101;
   26000: result <= 12'b010011010101;
   26001: result <= 12'b010011010101;
   26002: result <= 12'b010011010101;
   26003: result <= 12'b010011010101;
   26004: result <= 12'b010011010100;
   26005: result <= 12'b010011010100;
   26006: result <= 12'b010011010100;
   26007: result <= 12'b010011010100;
   26008: result <= 12'b010011010100;
   26009: result <= 12'b010011010100;
   26010: result <= 12'b010011010100;
   26011: result <= 12'b010011010011;
   26012: result <= 12'b010011010011;
   26013: result <= 12'b010011010011;
   26014: result <= 12'b010011010011;
   26015: result <= 12'b010011010011;
   26016: result <= 12'b010011010011;
   26017: result <= 12'b010011010010;
   26018: result <= 12'b010011010010;
   26019: result <= 12'b010011010010;
   26020: result <= 12'b010011010010;
   26021: result <= 12'b010011010010;
   26022: result <= 12'b010011010010;
   26023: result <= 12'b010011010001;
   26024: result <= 12'b010011010001;
   26025: result <= 12'b010011010001;
   26026: result <= 12'b010011010001;
   26027: result <= 12'b010011010001;
   26028: result <= 12'b010011010001;
   26029: result <= 12'b010011010001;
   26030: result <= 12'b010011010000;
   26031: result <= 12'b010011010000;
   26032: result <= 12'b010011010000;
   26033: result <= 12'b010011010000;
   26034: result <= 12'b010011010000;
   26035: result <= 12'b010011010000;
   26036: result <= 12'b010011001111;
   26037: result <= 12'b010011001111;
   26038: result <= 12'b010011001111;
   26039: result <= 12'b010011001111;
   26040: result <= 12'b010011001111;
   26041: result <= 12'b010011001111;
   26042: result <= 12'b010011001111;
   26043: result <= 12'b010011001110;
   26044: result <= 12'b010011001110;
   26045: result <= 12'b010011001110;
   26046: result <= 12'b010011001110;
   26047: result <= 12'b010011001110;
   26048: result <= 12'b010011001110;
   26049: result <= 12'b010011001101;
   26050: result <= 12'b010011001101;
   26051: result <= 12'b010011001101;
   26052: result <= 12'b010011001101;
   26053: result <= 12'b010011001101;
   26054: result <= 12'b010011001101;
   26055: result <= 12'b010011001100;
   26056: result <= 12'b010011001100;
   26057: result <= 12'b010011001100;
   26058: result <= 12'b010011001100;
   26059: result <= 12'b010011001100;
   26060: result <= 12'b010011001100;
   26061: result <= 12'b010011001100;
   26062: result <= 12'b010011001011;
   26063: result <= 12'b010011001011;
   26064: result <= 12'b010011001011;
   26065: result <= 12'b010011001011;
   26066: result <= 12'b010011001011;
   26067: result <= 12'b010011001011;
   26068: result <= 12'b010011001010;
   26069: result <= 12'b010011001010;
   26070: result <= 12'b010011001010;
   26071: result <= 12'b010011001010;
   26072: result <= 12'b010011001010;
   26073: result <= 12'b010011001010;
   26074: result <= 12'b010011001001;
   26075: result <= 12'b010011001001;
   26076: result <= 12'b010011001001;
   26077: result <= 12'b010011001001;
   26078: result <= 12'b010011001001;
   26079: result <= 12'b010011001001;
   26080: result <= 12'b010011001001;
   26081: result <= 12'b010011001000;
   26082: result <= 12'b010011001000;
   26083: result <= 12'b010011001000;
   26084: result <= 12'b010011001000;
   26085: result <= 12'b010011001000;
   26086: result <= 12'b010011001000;
   26087: result <= 12'b010011000111;
   26088: result <= 12'b010011000111;
   26089: result <= 12'b010011000111;
   26090: result <= 12'b010011000111;
   26091: result <= 12'b010011000111;
   26092: result <= 12'b010011000111;
   26093: result <= 12'b010011000110;
   26094: result <= 12'b010011000110;
   26095: result <= 12'b010011000110;
   26096: result <= 12'b010011000110;
   26097: result <= 12'b010011000110;
   26098: result <= 12'b010011000110;
   26099: result <= 12'b010011000110;
   26100: result <= 12'b010011000101;
   26101: result <= 12'b010011000101;
   26102: result <= 12'b010011000101;
   26103: result <= 12'b010011000101;
   26104: result <= 12'b010011000101;
   26105: result <= 12'b010011000101;
   26106: result <= 12'b010011000100;
   26107: result <= 12'b010011000100;
   26108: result <= 12'b010011000100;
   26109: result <= 12'b010011000100;
   26110: result <= 12'b010011000100;
   26111: result <= 12'b010011000100;
   26112: result <= 12'b010011000011;
   26113: result <= 12'b010011000011;
   26114: result <= 12'b010011000011;
   26115: result <= 12'b010011000011;
   26116: result <= 12'b010011000011;
   26117: result <= 12'b010011000011;
   26118: result <= 12'b010011000011;
   26119: result <= 12'b010011000010;
   26120: result <= 12'b010011000010;
   26121: result <= 12'b010011000010;
   26122: result <= 12'b010011000010;
   26123: result <= 12'b010011000010;
   26124: result <= 12'b010011000010;
   26125: result <= 12'b010011000001;
   26126: result <= 12'b010011000001;
   26127: result <= 12'b010011000001;
   26128: result <= 12'b010011000001;
   26129: result <= 12'b010011000001;
   26130: result <= 12'b010011000001;
   26131: result <= 12'b010011000000;
   26132: result <= 12'b010011000000;
   26133: result <= 12'b010011000000;
   26134: result <= 12'b010011000000;
   26135: result <= 12'b010011000000;
   26136: result <= 12'b010011000000;
   26137: result <= 12'b010011000000;
   26138: result <= 12'b010010111111;
   26139: result <= 12'b010010111111;
   26140: result <= 12'b010010111111;
   26141: result <= 12'b010010111111;
   26142: result <= 12'b010010111111;
   26143: result <= 12'b010010111111;
   26144: result <= 12'b010010111110;
   26145: result <= 12'b010010111110;
   26146: result <= 12'b010010111110;
   26147: result <= 12'b010010111110;
   26148: result <= 12'b010010111110;
   26149: result <= 12'b010010111110;
   26150: result <= 12'b010010111101;
   26151: result <= 12'b010010111101;
   26152: result <= 12'b010010111101;
   26153: result <= 12'b010010111101;
   26154: result <= 12'b010010111101;
   26155: result <= 12'b010010111101;
   26156: result <= 12'b010010111101;
   26157: result <= 12'b010010111100;
   26158: result <= 12'b010010111100;
   26159: result <= 12'b010010111100;
   26160: result <= 12'b010010111100;
   26161: result <= 12'b010010111100;
   26162: result <= 12'b010010111100;
   26163: result <= 12'b010010111011;
   26164: result <= 12'b010010111011;
   26165: result <= 12'b010010111011;
   26166: result <= 12'b010010111011;
   26167: result <= 12'b010010111011;
   26168: result <= 12'b010010111011;
   26169: result <= 12'b010010111010;
   26170: result <= 12'b010010111010;
   26171: result <= 12'b010010111010;
   26172: result <= 12'b010010111010;
   26173: result <= 12'b010010111010;
   26174: result <= 12'b010010111010;
   26175: result <= 12'b010010111010;
   26176: result <= 12'b010010111001;
   26177: result <= 12'b010010111001;
   26178: result <= 12'b010010111001;
   26179: result <= 12'b010010111001;
   26180: result <= 12'b010010111001;
   26181: result <= 12'b010010111001;
   26182: result <= 12'b010010111000;
   26183: result <= 12'b010010111000;
   26184: result <= 12'b010010111000;
   26185: result <= 12'b010010111000;
   26186: result <= 12'b010010111000;
   26187: result <= 12'b010010111000;
   26188: result <= 12'b010010110111;
   26189: result <= 12'b010010110111;
   26190: result <= 12'b010010110111;
   26191: result <= 12'b010010110111;
   26192: result <= 12'b010010110111;
   26193: result <= 12'b010010110111;
   26194: result <= 12'b010010110111;
   26195: result <= 12'b010010110110;
   26196: result <= 12'b010010110110;
   26197: result <= 12'b010010110110;
   26198: result <= 12'b010010110110;
   26199: result <= 12'b010010110110;
   26200: result <= 12'b010010110110;
   26201: result <= 12'b010010110101;
   26202: result <= 12'b010010110101;
   26203: result <= 12'b010010110101;
   26204: result <= 12'b010010110101;
   26205: result <= 12'b010010110101;
   26206: result <= 12'b010010110101;
   26207: result <= 12'b010010110100;
   26208: result <= 12'b010010110100;
   26209: result <= 12'b010010110100;
   26210: result <= 12'b010010110100;
   26211: result <= 12'b010010110100;
   26212: result <= 12'b010010110100;
   26213: result <= 12'b010010110100;
   26214: result <= 12'b010010110011;
   26215: result <= 12'b010010110011;
   26216: result <= 12'b010010110011;
   26217: result <= 12'b010010110011;
   26218: result <= 12'b010010110011;
   26219: result <= 12'b010010110011;
   26220: result <= 12'b010010110010;
   26221: result <= 12'b010010110010;
   26222: result <= 12'b010010110010;
   26223: result <= 12'b010010110010;
   26224: result <= 12'b010010110010;
   26225: result <= 12'b010010110010;
   26226: result <= 12'b010010110001;
   26227: result <= 12'b010010110001;
   26228: result <= 12'b010010110001;
   26229: result <= 12'b010010110001;
   26230: result <= 12'b010010110001;
   26231: result <= 12'b010010110001;
   26232: result <= 12'b010010110000;
   26233: result <= 12'b010010110000;
   26234: result <= 12'b010010110000;
   26235: result <= 12'b010010110000;
   26236: result <= 12'b010010110000;
   26237: result <= 12'b010010110000;
   26238: result <= 12'b010010110000;
   26239: result <= 12'b010010101111;
   26240: result <= 12'b010010101111;
   26241: result <= 12'b010010101111;
   26242: result <= 12'b010010101111;
   26243: result <= 12'b010010101111;
   26244: result <= 12'b010010101111;
   26245: result <= 12'b010010101110;
   26246: result <= 12'b010010101110;
   26247: result <= 12'b010010101110;
   26248: result <= 12'b010010101110;
   26249: result <= 12'b010010101110;
   26250: result <= 12'b010010101110;
   26251: result <= 12'b010010101101;
   26252: result <= 12'b010010101101;
   26253: result <= 12'b010010101101;
   26254: result <= 12'b010010101101;
   26255: result <= 12'b010010101101;
   26256: result <= 12'b010010101101;
   26257: result <= 12'b010010101101;
   26258: result <= 12'b010010101100;
   26259: result <= 12'b010010101100;
   26260: result <= 12'b010010101100;
   26261: result <= 12'b010010101100;
   26262: result <= 12'b010010101100;
   26263: result <= 12'b010010101100;
   26264: result <= 12'b010010101011;
   26265: result <= 12'b010010101011;
   26266: result <= 12'b010010101011;
   26267: result <= 12'b010010101011;
   26268: result <= 12'b010010101011;
   26269: result <= 12'b010010101011;
   26270: result <= 12'b010010101010;
   26271: result <= 12'b010010101010;
   26272: result <= 12'b010010101010;
   26273: result <= 12'b010010101010;
   26274: result <= 12'b010010101010;
   26275: result <= 12'b010010101010;
   26276: result <= 12'b010010101001;
   26277: result <= 12'b010010101001;
   26278: result <= 12'b010010101001;
   26279: result <= 12'b010010101001;
   26280: result <= 12'b010010101001;
   26281: result <= 12'b010010101001;
   26282: result <= 12'b010010101001;
   26283: result <= 12'b010010101000;
   26284: result <= 12'b010010101000;
   26285: result <= 12'b010010101000;
   26286: result <= 12'b010010101000;
   26287: result <= 12'b010010101000;
   26288: result <= 12'b010010101000;
   26289: result <= 12'b010010100111;
   26290: result <= 12'b010010100111;
   26291: result <= 12'b010010100111;
   26292: result <= 12'b010010100111;
   26293: result <= 12'b010010100111;
   26294: result <= 12'b010010100111;
   26295: result <= 12'b010010100110;
   26296: result <= 12'b010010100110;
   26297: result <= 12'b010010100110;
   26298: result <= 12'b010010100110;
   26299: result <= 12'b010010100110;
   26300: result <= 12'b010010100110;
   26301: result <= 12'b010010100101;
   26302: result <= 12'b010010100101;
   26303: result <= 12'b010010100101;
   26304: result <= 12'b010010100101;
   26305: result <= 12'b010010100101;
   26306: result <= 12'b010010100101;
   26307: result <= 12'b010010100101;
   26308: result <= 12'b010010100100;
   26309: result <= 12'b010010100100;
   26310: result <= 12'b010010100100;
   26311: result <= 12'b010010100100;
   26312: result <= 12'b010010100100;
   26313: result <= 12'b010010100100;
   26314: result <= 12'b010010100011;
   26315: result <= 12'b010010100011;
   26316: result <= 12'b010010100011;
   26317: result <= 12'b010010100011;
   26318: result <= 12'b010010100011;
   26319: result <= 12'b010010100011;
   26320: result <= 12'b010010100010;
   26321: result <= 12'b010010100010;
   26322: result <= 12'b010010100010;
   26323: result <= 12'b010010100010;
   26324: result <= 12'b010010100010;
   26325: result <= 12'b010010100010;
   26326: result <= 12'b010010100001;
   26327: result <= 12'b010010100001;
   26328: result <= 12'b010010100001;
   26329: result <= 12'b010010100001;
   26330: result <= 12'b010010100001;
   26331: result <= 12'b010010100001;
   26332: result <= 12'b010010100001;
   26333: result <= 12'b010010100000;
   26334: result <= 12'b010010100000;
   26335: result <= 12'b010010100000;
   26336: result <= 12'b010010100000;
   26337: result <= 12'b010010100000;
   26338: result <= 12'b010010100000;
   26339: result <= 12'b010010011111;
   26340: result <= 12'b010010011111;
   26341: result <= 12'b010010011111;
   26342: result <= 12'b010010011111;
   26343: result <= 12'b010010011111;
   26344: result <= 12'b010010011111;
   26345: result <= 12'b010010011110;
   26346: result <= 12'b010010011110;
   26347: result <= 12'b010010011110;
   26348: result <= 12'b010010011110;
   26349: result <= 12'b010010011110;
   26350: result <= 12'b010010011110;
   26351: result <= 12'b010010011101;
   26352: result <= 12'b010010011101;
   26353: result <= 12'b010010011101;
   26354: result <= 12'b010010011101;
   26355: result <= 12'b010010011101;
   26356: result <= 12'b010010011101;
   26357: result <= 12'b010010011101;
   26358: result <= 12'b010010011100;
   26359: result <= 12'b010010011100;
   26360: result <= 12'b010010011100;
   26361: result <= 12'b010010011100;
   26362: result <= 12'b010010011100;
   26363: result <= 12'b010010011100;
   26364: result <= 12'b010010011011;
   26365: result <= 12'b010010011011;
   26366: result <= 12'b010010011011;
   26367: result <= 12'b010010011011;
   26368: result <= 12'b010010011011;
   26369: result <= 12'b010010011011;
   26370: result <= 12'b010010011010;
   26371: result <= 12'b010010011010;
   26372: result <= 12'b010010011010;
   26373: result <= 12'b010010011010;
   26374: result <= 12'b010010011010;
   26375: result <= 12'b010010011010;
   26376: result <= 12'b010010011001;
   26377: result <= 12'b010010011001;
   26378: result <= 12'b010010011001;
   26379: result <= 12'b010010011001;
   26380: result <= 12'b010010011001;
   26381: result <= 12'b010010011001;
   26382: result <= 12'b010010011001;
   26383: result <= 12'b010010011000;
   26384: result <= 12'b010010011000;
   26385: result <= 12'b010010011000;
   26386: result <= 12'b010010011000;
   26387: result <= 12'b010010011000;
   26388: result <= 12'b010010011000;
   26389: result <= 12'b010010010111;
   26390: result <= 12'b010010010111;
   26391: result <= 12'b010010010111;
   26392: result <= 12'b010010010111;
   26393: result <= 12'b010010010111;
   26394: result <= 12'b010010010111;
   26395: result <= 12'b010010010110;
   26396: result <= 12'b010010010110;
   26397: result <= 12'b010010010110;
   26398: result <= 12'b010010010110;
   26399: result <= 12'b010010010110;
   26400: result <= 12'b010010010110;
   26401: result <= 12'b010010010101;
   26402: result <= 12'b010010010101;
   26403: result <= 12'b010010010101;
   26404: result <= 12'b010010010101;
   26405: result <= 12'b010010010101;
   26406: result <= 12'b010010010101;
   26407: result <= 12'b010010010100;
   26408: result <= 12'b010010010100;
   26409: result <= 12'b010010010100;
   26410: result <= 12'b010010010100;
   26411: result <= 12'b010010010100;
   26412: result <= 12'b010010010100;
   26413: result <= 12'b010010010100;
   26414: result <= 12'b010010010011;
   26415: result <= 12'b010010010011;
   26416: result <= 12'b010010010011;
   26417: result <= 12'b010010010011;
   26418: result <= 12'b010010010011;
   26419: result <= 12'b010010010011;
   26420: result <= 12'b010010010010;
   26421: result <= 12'b010010010010;
   26422: result <= 12'b010010010010;
   26423: result <= 12'b010010010010;
   26424: result <= 12'b010010010010;
   26425: result <= 12'b010010010010;
   26426: result <= 12'b010010010001;
   26427: result <= 12'b010010010001;
   26428: result <= 12'b010010010001;
   26429: result <= 12'b010010010001;
   26430: result <= 12'b010010010001;
   26431: result <= 12'b010010010001;
   26432: result <= 12'b010010010000;
   26433: result <= 12'b010010010000;
   26434: result <= 12'b010010010000;
   26435: result <= 12'b010010010000;
   26436: result <= 12'b010010010000;
   26437: result <= 12'b010010010000;
   26438: result <= 12'b010010001111;
   26439: result <= 12'b010010001111;
   26440: result <= 12'b010010001111;
   26441: result <= 12'b010010001111;
   26442: result <= 12'b010010001111;
   26443: result <= 12'b010010001111;
   26444: result <= 12'b010010001111;
   26445: result <= 12'b010010001110;
   26446: result <= 12'b010010001110;
   26447: result <= 12'b010010001110;
   26448: result <= 12'b010010001110;
   26449: result <= 12'b010010001110;
   26450: result <= 12'b010010001110;
   26451: result <= 12'b010010001101;
   26452: result <= 12'b010010001101;
   26453: result <= 12'b010010001101;
   26454: result <= 12'b010010001101;
   26455: result <= 12'b010010001101;
   26456: result <= 12'b010010001101;
   26457: result <= 12'b010010001100;
   26458: result <= 12'b010010001100;
   26459: result <= 12'b010010001100;
   26460: result <= 12'b010010001100;
   26461: result <= 12'b010010001100;
   26462: result <= 12'b010010001100;
   26463: result <= 12'b010010001011;
   26464: result <= 12'b010010001011;
   26465: result <= 12'b010010001011;
   26466: result <= 12'b010010001011;
   26467: result <= 12'b010010001011;
   26468: result <= 12'b010010001011;
   26469: result <= 12'b010010001010;
   26470: result <= 12'b010010001010;
   26471: result <= 12'b010010001010;
   26472: result <= 12'b010010001010;
   26473: result <= 12'b010010001010;
   26474: result <= 12'b010010001010;
   26475: result <= 12'b010010001010;
   26476: result <= 12'b010010001001;
   26477: result <= 12'b010010001001;
   26478: result <= 12'b010010001001;
   26479: result <= 12'b010010001001;
   26480: result <= 12'b010010001001;
   26481: result <= 12'b010010001001;
   26482: result <= 12'b010010001000;
   26483: result <= 12'b010010001000;
   26484: result <= 12'b010010001000;
   26485: result <= 12'b010010001000;
   26486: result <= 12'b010010001000;
   26487: result <= 12'b010010001000;
   26488: result <= 12'b010010000111;
   26489: result <= 12'b010010000111;
   26490: result <= 12'b010010000111;
   26491: result <= 12'b010010000111;
   26492: result <= 12'b010010000111;
   26493: result <= 12'b010010000111;
   26494: result <= 12'b010010000110;
   26495: result <= 12'b010010000110;
   26496: result <= 12'b010010000110;
   26497: result <= 12'b010010000110;
   26498: result <= 12'b010010000110;
   26499: result <= 12'b010010000110;
   26500: result <= 12'b010010000101;
   26501: result <= 12'b010010000101;
   26502: result <= 12'b010010000101;
   26503: result <= 12'b010010000101;
   26504: result <= 12'b010010000101;
   26505: result <= 12'b010010000101;
   26506: result <= 12'b010010000100;
   26507: result <= 12'b010010000100;
   26508: result <= 12'b010010000100;
   26509: result <= 12'b010010000100;
   26510: result <= 12'b010010000100;
   26511: result <= 12'b010010000100;
   26512: result <= 12'b010010000100;
   26513: result <= 12'b010010000011;
   26514: result <= 12'b010010000011;
   26515: result <= 12'b010010000011;
   26516: result <= 12'b010010000011;
   26517: result <= 12'b010010000011;
   26518: result <= 12'b010010000011;
   26519: result <= 12'b010010000010;
   26520: result <= 12'b010010000010;
   26521: result <= 12'b010010000010;
   26522: result <= 12'b010010000010;
   26523: result <= 12'b010010000010;
   26524: result <= 12'b010010000010;
   26525: result <= 12'b010010000001;
   26526: result <= 12'b010010000001;
   26527: result <= 12'b010010000001;
   26528: result <= 12'b010010000001;
   26529: result <= 12'b010010000001;
   26530: result <= 12'b010010000001;
   26531: result <= 12'b010010000000;
   26532: result <= 12'b010010000000;
   26533: result <= 12'b010010000000;
   26534: result <= 12'b010010000000;
   26535: result <= 12'b010010000000;
   26536: result <= 12'b010010000000;
   26537: result <= 12'b010001111111;
   26538: result <= 12'b010001111111;
   26539: result <= 12'b010001111111;
   26540: result <= 12'b010001111111;
   26541: result <= 12'b010001111111;
   26542: result <= 12'b010001111111;
   26543: result <= 12'b010001111110;
   26544: result <= 12'b010001111110;
   26545: result <= 12'b010001111110;
   26546: result <= 12'b010001111110;
   26547: result <= 12'b010001111110;
   26548: result <= 12'b010001111110;
   26549: result <= 12'b010001111110;
   26550: result <= 12'b010001111101;
   26551: result <= 12'b010001111101;
   26552: result <= 12'b010001111101;
   26553: result <= 12'b010001111101;
   26554: result <= 12'b010001111101;
   26555: result <= 12'b010001111101;
   26556: result <= 12'b010001111100;
   26557: result <= 12'b010001111100;
   26558: result <= 12'b010001111100;
   26559: result <= 12'b010001111100;
   26560: result <= 12'b010001111100;
   26561: result <= 12'b010001111100;
   26562: result <= 12'b010001111011;
   26563: result <= 12'b010001111011;
   26564: result <= 12'b010001111011;
   26565: result <= 12'b010001111011;
   26566: result <= 12'b010001111011;
   26567: result <= 12'b010001111011;
   26568: result <= 12'b010001111010;
   26569: result <= 12'b010001111010;
   26570: result <= 12'b010001111010;
   26571: result <= 12'b010001111010;
   26572: result <= 12'b010001111010;
   26573: result <= 12'b010001111010;
   26574: result <= 12'b010001111001;
   26575: result <= 12'b010001111001;
   26576: result <= 12'b010001111001;
   26577: result <= 12'b010001111001;
   26578: result <= 12'b010001111001;
   26579: result <= 12'b010001111001;
   26580: result <= 12'b010001111000;
   26581: result <= 12'b010001111000;
   26582: result <= 12'b010001111000;
   26583: result <= 12'b010001111000;
   26584: result <= 12'b010001111000;
   26585: result <= 12'b010001111000;
   26586: result <= 12'b010001111000;
   26587: result <= 12'b010001110111;
   26588: result <= 12'b010001110111;
   26589: result <= 12'b010001110111;
   26590: result <= 12'b010001110111;
   26591: result <= 12'b010001110111;
   26592: result <= 12'b010001110111;
   26593: result <= 12'b010001110110;
   26594: result <= 12'b010001110110;
   26595: result <= 12'b010001110110;
   26596: result <= 12'b010001110110;
   26597: result <= 12'b010001110110;
   26598: result <= 12'b010001110110;
   26599: result <= 12'b010001110101;
   26600: result <= 12'b010001110101;
   26601: result <= 12'b010001110101;
   26602: result <= 12'b010001110101;
   26603: result <= 12'b010001110101;
   26604: result <= 12'b010001110101;
   26605: result <= 12'b010001110100;
   26606: result <= 12'b010001110100;
   26607: result <= 12'b010001110100;
   26608: result <= 12'b010001110100;
   26609: result <= 12'b010001110100;
   26610: result <= 12'b010001110100;
   26611: result <= 12'b010001110011;
   26612: result <= 12'b010001110011;
   26613: result <= 12'b010001110011;
   26614: result <= 12'b010001110011;
   26615: result <= 12'b010001110011;
   26616: result <= 12'b010001110011;
   26617: result <= 12'b010001110010;
   26618: result <= 12'b010001110010;
   26619: result <= 12'b010001110010;
   26620: result <= 12'b010001110010;
   26621: result <= 12'b010001110010;
   26622: result <= 12'b010001110010;
   26623: result <= 12'b010001110001;
   26624: result <= 12'b010001110001;
   26625: result <= 12'b010001110001;
   26626: result <= 12'b010001110001;
   26627: result <= 12'b010001110001;
   26628: result <= 12'b010001110001;
   26629: result <= 12'b010001110000;
   26630: result <= 12'b010001110000;
   26631: result <= 12'b010001110000;
   26632: result <= 12'b010001110000;
   26633: result <= 12'b010001110000;
   26634: result <= 12'b010001110000;
   26635: result <= 12'b010001110000;
   26636: result <= 12'b010001101111;
   26637: result <= 12'b010001101111;
   26638: result <= 12'b010001101111;
   26639: result <= 12'b010001101111;
   26640: result <= 12'b010001101111;
   26641: result <= 12'b010001101111;
   26642: result <= 12'b010001101110;
   26643: result <= 12'b010001101110;
   26644: result <= 12'b010001101110;
   26645: result <= 12'b010001101110;
   26646: result <= 12'b010001101110;
   26647: result <= 12'b010001101110;
   26648: result <= 12'b010001101101;
   26649: result <= 12'b010001101101;
   26650: result <= 12'b010001101101;
   26651: result <= 12'b010001101101;
   26652: result <= 12'b010001101101;
   26653: result <= 12'b010001101101;
   26654: result <= 12'b010001101100;
   26655: result <= 12'b010001101100;
   26656: result <= 12'b010001101100;
   26657: result <= 12'b010001101100;
   26658: result <= 12'b010001101100;
   26659: result <= 12'b010001101100;
   26660: result <= 12'b010001101011;
   26661: result <= 12'b010001101011;
   26662: result <= 12'b010001101011;
   26663: result <= 12'b010001101011;
   26664: result <= 12'b010001101011;
   26665: result <= 12'b010001101011;
   26666: result <= 12'b010001101010;
   26667: result <= 12'b010001101010;
   26668: result <= 12'b010001101010;
   26669: result <= 12'b010001101010;
   26670: result <= 12'b010001101010;
   26671: result <= 12'b010001101010;
   26672: result <= 12'b010001101001;
   26673: result <= 12'b010001101001;
   26674: result <= 12'b010001101001;
   26675: result <= 12'b010001101001;
   26676: result <= 12'b010001101001;
   26677: result <= 12'b010001101001;
   26678: result <= 12'b010001101000;
   26679: result <= 12'b010001101000;
   26680: result <= 12'b010001101000;
   26681: result <= 12'b010001101000;
   26682: result <= 12'b010001101000;
   26683: result <= 12'b010001101000;
   26684: result <= 12'b010001100111;
   26685: result <= 12'b010001100111;
   26686: result <= 12'b010001100111;
   26687: result <= 12'b010001100111;
   26688: result <= 12'b010001100111;
   26689: result <= 12'b010001100111;
   26690: result <= 12'b010001100111;
   26691: result <= 12'b010001100110;
   26692: result <= 12'b010001100110;
   26693: result <= 12'b010001100110;
   26694: result <= 12'b010001100110;
   26695: result <= 12'b010001100110;
   26696: result <= 12'b010001100110;
   26697: result <= 12'b010001100101;
   26698: result <= 12'b010001100101;
   26699: result <= 12'b010001100101;
   26700: result <= 12'b010001100101;
   26701: result <= 12'b010001100101;
   26702: result <= 12'b010001100101;
   26703: result <= 12'b010001100100;
   26704: result <= 12'b010001100100;
   26705: result <= 12'b010001100100;
   26706: result <= 12'b010001100100;
   26707: result <= 12'b010001100100;
   26708: result <= 12'b010001100100;
   26709: result <= 12'b010001100011;
   26710: result <= 12'b010001100011;
   26711: result <= 12'b010001100011;
   26712: result <= 12'b010001100011;
   26713: result <= 12'b010001100011;
   26714: result <= 12'b010001100011;
   26715: result <= 12'b010001100010;
   26716: result <= 12'b010001100010;
   26717: result <= 12'b010001100010;
   26718: result <= 12'b010001100010;
   26719: result <= 12'b010001100010;
   26720: result <= 12'b010001100010;
   26721: result <= 12'b010001100001;
   26722: result <= 12'b010001100001;
   26723: result <= 12'b010001100001;
   26724: result <= 12'b010001100001;
   26725: result <= 12'b010001100001;
   26726: result <= 12'b010001100001;
   26727: result <= 12'b010001100000;
   26728: result <= 12'b010001100000;
   26729: result <= 12'b010001100000;
   26730: result <= 12'b010001100000;
   26731: result <= 12'b010001100000;
   26732: result <= 12'b010001100000;
   26733: result <= 12'b010001011111;
   26734: result <= 12'b010001011111;
   26735: result <= 12'b010001011111;
   26736: result <= 12'b010001011111;
   26737: result <= 12'b010001011111;
   26738: result <= 12'b010001011111;
   26739: result <= 12'b010001011110;
   26740: result <= 12'b010001011110;
   26741: result <= 12'b010001011110;
   26742: result <= 12'b010001011110;
   26743: result <= 12'b010001011110;
   26744: result <= 12'b010001011110;
   26745: result <= 12'b010001011101;
   26746: result <= 12'b010001011101;
   26747: result <= 12'b010001011101;
   26748: result <= 12'b010001011101;
   26749: result <= 12'b010001011101;
   26750: result <= 12'b010001011101;
   26751: result <= 12'b010001011100;
   26752: result <= 12'b010001011100;
   26753: result <= 12'b010001011100;
   26754: result <= 12'b010001011100;
   26755: result <= 12'b010001011100;
   26756: result <= 12'b010001011100;
   26757: result <= 12'b010001011100;
   26758: result <= 12'b010001011011;
   26759: result <= 12'b010001011011;
   26760: result <= 12'b010001011011;
   26761: result <= 12'b010001011011;
   26762: result <= 12'b010001011011;
   26763: result <= 12'b010001011011;
   26764: result <= 12'b010001011010;
   26765: result <= 12'b010001011010;
   26766: result <= 12'b010001011010;
   26767: result <= 12'b010001011010;
   26768: result <= 12'b010001011010;
   26769: result <= 12'b010001011010;
   26770: result <= 12'b010001011001;
   26771: result <= 12'b010001011001;
   26772: result <= 12'b010001011001;
   26773: result <= 12'b010001011001;
   26774: result <= 12'b010001011001;
   26775: result <= 12'b010001011001;
   26776: result <= 12'b010001011000;
   26777: result <= 12'b010001011000;
   26778: result <= 12'b010001011000;
   26779: result <= 12'b010001011000;
   26780: result <= 12'b010001011000;
   26781: result <= 12'b010001011000;
   26782: result <= 12'b010001010111;
   26783: result <= 12'b010001010111;
   26784: result <= 12'b010001010111;
   26785: result <= 12'b010001010111;
   26786: result <= 12'b010001010111;
   26787: result <= 12'b010001010111;
   26788: result <= 12'b010001010110;
   26789: result <= 12'b010001010110;
   26790: result <= 12'b010001010110;
   26791: result <= 12'b010001010110;
   26792: result <= 12'b010001010110;
   26793: result <= 12'b010001010110;
   26794: result <= 12'b010001010101;
   26795: result <= 12'b010001010101;
   26796: result <= 12'b010001010101;
   26797: result <= 12'b010001010101;
   26798: result <= 12'b010001010101;
   26799: result <= 12'b010001010101;
   26800: result <= 12'b010001010100;
   26801: result <= 12'b010001010100;
   26802: result <= 12'b010001010100;
   26803: result <= 12'b010001010100;
   26804: result <= 12'b010001010100;
   26805: result <= 12'b010001010100;
   26806: result <= 12'b010001010011;
   26807: result <= 12'b010001010011;
   26808: result <= 12'b010001010011;
   26809: result <= 12'b010001010011;
   26810: result <= 12'b010001010011;
   26811: result <= 12'b010001010011;
   26812: result <= 12'b010001010010;
   26813: result <= 12'b010001010010;
   26814: result <= 12'b010001010010;
   26815: result <= 12'b010001010010;
   26816: result <= 12'b010001010010;
   26817: result <= 12'b010001010010;
   26818: result <= 12'b010001010001;
   26819: result <= 12'b010001010001;
   26820: result <= 12'b010001010001;
   26821: result <= 12'b010001010001;
   26822: result <= 12'b010001010001;
   26823: result <= 12'b010001010001;
   26824: result <= 12'b010001010000;
   26825: result <= 12'b010001010000;
   26826: result <= 12'b010001010000;
   26827: result <= 12'b010001010000;
   26828: result <= 12'b010001010000;
   26829: result <= 12'b010001010000;
   26830: result <= 12'b010001001111;
   26831: result <= 12'b010001001111;
   26832: result <= 12'b010001001111;
   26833: result <= 12'b010001001111;
   26834: result <= 12'b010001001111;
   26835: result <= 12'b010001001111;
   26836: result <= 12'b010001001110;
   26837: result <= 12'b010001001110;
   26838: result <= 12'b010001001110;
   26839: result <= 12'b010001001110;
   26840: result <= 12'b010001001110;
   26841: result <= 12'b010001001110;
   26842: result <= 12'b010001001101;
   26843: result <= 12'b010001001101;
   26844: result <= 12'b010001001101;
   26845: result <= 12'b010001001101;
   26846: result <= 12'b010001001101;
   26847: result <= 12'b010001001101;
   26848: result <= 12'b010001001100;
   26849: result <= 12'b010001001100;
   26850: result <= 12'b010001001100;
   26851: result <= 12'b010001001100;
   26852: result <= 12'b010001001100;
   26853: result <= 12'b010001001100;
   26854: result <= 12'b010001001011;
   26855: result <= 12'b010001001011;
   26856: result <= 12'b010001001011;
   26857: result <= 12'b010001001011;
   26858: result <= 12'b010001001011;
   26859: result <= 12'b010001001011;
   26860: result <= 12'b010001001010;
   26861: result <= 12'b010001001010;
   26862: result <= 12'b010001001010;
   26863: result <= 12'b010001001010;
   26864: result <= 12'b010001001010;
   26865: result <= 12'b010001001010;
   26866: result <= 12'b010001001001;
   26867: result <= 12'b010001001001;
   26868: result <= 12'b010001001001;
   26869: result <= 12'b010001001001;
   26870: result <= 12'b010001001001;
   26871: result <= 12'b010001001001;
   26872: result <= 12'b010001001001;
   26873: result <= 12'b010001001000;
   26874: result <= 12'b010001001000;
   26875: result <= 12'b010001001000;
   26876: result <= 12'b010001001000;
   26877: result <= 12'b010001001000;
   26878: result <= 12'b010001001000;
   26879: result <= 12'b010001000111;
   26880: result <= 12'b010001000111;
   26881: result <= 12'b010001000111;
   26882: result <= 12'b010001000111;
   26883: result <= 12'b010001000111;
   26884: result <= 12'b010001000111;
   26885: result <= 12'b010001000110;
   26886: result <= 12'b010001000110;
   26887: result <= 12'b010001000110;
   26888: result <= 12'b010001000110;
   26889: result <= 12'b010001000110;
   26890: result <= 12'b010001000110;
   26891: result <= 12'b010001000101;
   26892: result <= 12'b010001000101;
   26893: result <= 12'b010001000101;
   26894: result <= 12'b010001000101;
   26895: result <= 12'b010001000101;
   26896: result <= 12'b010001000101;
   26897: result <= 12'b010001000100;
   26898: result <= 12'b010001000100;
   26899: result <= 12'b010001000100;
   26900: result <= 12'b010001000100;
   26901: result <= 12'b010001000100;
   26902: result <= 12'b010001000100;
   26903: result <= 12'b010001000011;
   26904: result <= 12'b010001000011;
   26905: result <= 12'b010001000011;
   26906: result <= 12'b010001000011;
   26907: result <= 12'b010001000011;
   26908: result <= 12'b010001000011;
   26909: result <= 12'b010001000010;
   26910: result <= 12'b010001000010;
   26911: result <= 12'b010001000010;
   26912: result <= 12'b010001000010;
   26913: result <= 12'b010001000010;
   26914: result <= 12'b010001000010;
   26915: result <= 12'b010001000001;
   26916: result <= 12'b010001000001;
   26917: result <= 12'b010001000001;
   26918: result <= 12'b010001000001;
   26919: result <= 12'b010001000001;
   26920: result <= 12'b010001000001;
   26921: result <= 12'b010001000000;
   26922: result <= 12'b010001000000;
   26923: result <= 12'b010001000000;
   26924: result <= 12'b010001000000;
   26925: result <= 12'b010001000000;
   26926: result <= 12'b010001000000;
   26927: result <= 12'b010000111111;
   26928: result <= 12'b010000111111;
   26929: result <= 12'b010000111111;
   26930: result <= 12'b010000111111;
   26931: result <= 12'b010000111111;
   26932: result <= 12'b010000111111;
   26933: result <= 12'b010000111110;
   26934: result <= 12'b010000111110;
   26935: result <= 12'b010000111110;
   26936: result <= 12'b010000111110;
   26937: result <= 12'b010000111110;
   26938: result <= 12'b010000111110;
   26939: result <= 12'b010000111101;
   26940: result <= 12'b010000111101;
   26941: result <= 12'b010000111101;
   26942: result <= 12'b010000111101;
   26943: result <= 12'b010000111101;
   26944: result <= 12'b010000111101;
   26945: result <= 12'b010000111100;
   26946: result <= 12'b010000111100;
   26947: result <= 12'b010000111100;
   26948: result <= 12'b010000111100;
   26949: result <= 12'b010000111100;
   26950: result <= 12'b010000111100;
   26951: result <= 12'b010000111011;
   26952: result <= 12'b010000111011;
   26953: result <= 12'b010000111011;
   26954: result <= 12'b010000111011;
   26955: result <= 12'b010000111011;
   26956: result <= 12'b010000111011;
   26957: result <= 12'b010000111010;
   26958: result <= 12'b010000111010;
   26959: result <= 12'b010000111010;
   26960: result <= 12'b010000111010;
   26961: result <= 12'b010000111010;
   26962: result <= 12'b010000111010;
   26963: result <= 12'b010000111001;
   26964: result <= 12'b010000111001;
   26965: result <= 12'b010000111001;
   26966: result <= 12'b010000111001;
   26967: result <= 12'b010000111001;
   26968: result <= 12'b010000111001;
   26969: result <= 12'b010000111000;
   26970: result <= 12'b010000111000;
   26971: result <= 12'b010000111000;
   26972: result <= 12'b010000111000;
   26973: result <= 12'b010000111000;
   26974: result <= 12'b010000111000;
   26975: result <= 12'b010000110111;
   26976: result <= 12'b010000110111;
   26977: result <= 12'b010000110111;
   26978: result <= 12'b010000110111;
   26979: result <= 12'b010000110111;
   26980: result <= 12'b010000110111;
   26981: result <= 12'b010000110110;
   26982: result <= 12'b010000110110;
   26983: result <= 12'b010000110110;
   26984: result <= 12'b010000110110;
   26985: result <= 12'b010000110110;
   26986: result <= 12'b010000110110;
   26987: result <= 12'b010000110101;
   26988: result <= 12'b010000110101;
   26989: result <= 12'b010000110101;
   26990: result <= 12'b010000110101;
   26991: result <= 12'b010000110101;
   26992: result <= 12'b010000110101;
   26993: result <= 12'b010000110100;
   26994: result <= 12'b010000110100;
   26995: result <= 12'b010000110100;
   26996: result <= 12'b010000110100;
   26997: result <= 12'b010000110100;
   26998: result <= 12'b010000110100;
   26999: result <= 12'b010000110011;
   27000: result <= 12'b010000110011;
   27001: result <= 12'b010000110011;
   27002: result <= 12'b010000110011;
   27003: result <= 12'b010000110011;
   27004: result <= 12'b010000110011;
   27005: result <= 12'b010000110010;
   27006: result <= 12'b010000110010;
   27007: result <= 12'b010000110010;
   27008: result <= 12'b010000110010;
   27009: result <= 12'b010000110010;
   27010: result <= 12'b010000110010;
   27011: result <= 12'b010000110001;
   27012: result <= 12'b010000110001;
   27013: result <= 12'b010000110001;
   27014: result <= 12'b010000110001;
   27015: result <= 12'b010000110001;
   27016: result <= 12'b010000110001;
   27017: result <= 12'b010000110000;
   27018: result <= 12'b010000110000;
   27019: result <= 12'b010000110000;
   27020: result <= 12'b010000110000;
   27021: result <= 12'b010000110000;
   27022: result <= 12'b010000110000;
   27023: result <= 12'b010000101111;
   27024: result <= 12'b010000101111;
   27025: result <= 12'b010000101111;
   27026: result <= 12'b010000101111;
   27027: result <= 12'b010000101111;
   27028: result <= 12'b010000101111;
   27029: result <= 12'b010000101110;
   27030: result <= 12'b010000101110;
   27031: result <= 12'b010000101110;
   27032: result <= 12'b010000101110;
   27033: result <= 12'b010000101110;
   27034: result <= 12'b010000101110;
   27035: result <= 12'b010000101101;
   27036: result <= 12'b010000101101;
   27037: result <= 12'b010000101101;
   27038: result <= 12'b010000101101;
   27039: result <= 12'b010000101101;
   27040: result <= 12'b010000101101;
   27041: result <= 12'b010000101100;
   27042: result <= 12'b010000101100;
   27043: result <= 12'b010000101100;
   27044: result <= 12'b010000101100;
   27045: result <= 12'b010000101100;
   27046: result <= 12'b010000101100;
   27047: result <= 12'b010000101011;
   27048: result <= 12'b010000101011;
   27049: result <= 12'b010000101011;
   27050: result <= 12'b010000101011;
   27051: result <= 12'b010000101011;
   27052: result <= 12'b010000101010;
   27053: result <= 12'b010000101010;
   27054: result <= 12'b010000101010;
   27055: result <= 12'b010000101010;
   27056: result <= 12'b010000101010;
   27057: result <= 12'b010000101010;
   27058: result <= 12'b010000101001;
   27059: result <= 12'b010000101001;
   27060: result <= 12'b010000101001;
   27061: result <= 12'b010000101001;
   27062: result <= 12'b010000101001;
   27063: result <= 12'b010000101001;
   27064: result <= 12'b010000101000;
   27065: result <= 12'b010000101000;
   27066: result <= 12'b010000101000;
   27067: result <= 12'b010000101000;
   27068: result <= 12'b010000101000;
   27069: result <= 12'b010000101000;
   27070: result <= 12'b010000100111;
   27071: result <= 12'b010000100111;
   27072: result <= 12'b010000100111;
   27073: result <= 12'b010000100111;
   27074: result <= 12'b010000100111;
   27075: result <= 12'b010000100111;
   27076: result <= 12'b010000100110;
   27077: result <= 12'b010000100110;
   27078: result <= 12'b010000100110;
   27079: result <= 12'b010000100110;
   27080: result <= 12'b010000100110;
   27081: result <= 12'b010000100110;
   27082: result <= 12'b010000100101;
   27083: result <= 12'b010000100101;
   27084: result <= 12'b010000100101;
   27085: result <= 12'b010000100101;
   27086: result <= 12'b010000100101;
   27087: result <= 12'b010000100101;
   27088: result <= 12'b010000100100;
   27089: result <= 12'b010000100100;
   27090: result <= 12'b010000100100;
   27091: result <= 12'b010000100100;
   27092: result <= 12'b010000100100;
   27093: result <= 12'b010000100100;
   27094: result <= 12'b010000100011;
   27095: result <= 12'b010000100011;
   27096: result <= 12'b010000100011;
   27097: result <= 12'b010000100011;
   27098: result <= 12'b010000100011;
   27099: result <= 12'b010000100011;
   27100: result <= 12'b010000100010;
   27101: result <= 12'b010000100010;
   27102: result <= 12'b010000100010;
   27103: result <= 12'b010000100010;
   27104: result <= 12'b010000100010;
   27105: result <= 12'b010000100010;
   27106: result <= 12'b010000100001;
   27107: result <= 12'b010000100001;
   27108: result <= 12'b010000100001;
   27109: result <= 12'b010000100001;
   27110: result <= 12'b010000100001;
   27111: result <= 12'b010000100001;
   27112: result <= 12'b010000100000;
   27113: result <= 12'b010000100000;
   27114: result <= 12'b010000100000;
   27115: result <= 12'b010000100000;
   27116: result <= 12'b010000100000;
   27117: result <= 12'b010000100000;
   27118: result <= 12'b010000011111;
   27119: result <= 12'b010000011111;
   27120: result <= 12'b010000011111;
   27121: result <= 12'b010000011111;
   27122: result <= 12'b010000011111;
   27123: result <= 12'b010000011111;
   27124: result <= 12'b010000011110;
   27125: result <= 12'b010000011110;
   27126: result <= 12'b010000011110;
   27127: result <= 12'b010000011110;
   27128: result <= 12'b010000011110;
   27129: result <= 12'b010000011110;
   27130: result <= 12'b010000011101;
   27131: result <= 12'b010000011101;
   27132: result <= 12'b010000011101;
   27133: result <= 12'b010000011101;
   27134: result <= 12'b010000011101;
   27135: result <= 12'b010000011101;
   27136: result <= 12'b010000011100;
   27137: result <= 12'b010000011100;
   27138: result <= 12'b010000011100;
   27139: result <= 12'b010000011100;
   27140: result <= 12'b010000011100;
   27141: result <= 12'b010000011100;
   27142: result <= 12'b010000011011;
   27143: result <= 12'b010000011011;
   27144: result <= 12'b010000011011;
   27145: result <= 12'b010000011011;
   27146: result <= 12'b010000011011;
   27147: result <= 12'b010000011011;
   27148: result <= 12'b010000011010;
   27149: result <= 12'b010000011010;
   27150: result <= 12'b010000011010;
   27151: result <= 12'b010000011010;
   27152: result <= 12'b010000011010;
   27153: result <= 12'b010000011010;
   27154: result <= 12'b010000011001;
   27155: result <= 12'b010000011001;
   27156: result <= 12'b010000011001;
   27157: result <= 12'b010000011001;
   27158: result <= 12'b010000011001;
   27159: result <= 12'b010000011001;
   27160: result <= 12'b010000011000;
   27161: result <= 12'b010000011000;
   27162: result <= 12'b010000011000;
   27163: result <= 12'b010000011000;
   27164: result <= 12'b010000011000;
   27165: result <= 12'b010000010111;
   27166: result <= 12'b010000010111;
   27167: result <= 12'b010000010111;
   27168: result <= 12'b010000010111;
   27169: result <= 12'b010000010111;
   27170: result <= 12'b010000010111;
   27171: result <= 12'b010000010110;
   27172: result <= 12'b010000010110;
   27173: result <= 12'b010000010110;
   27174: result <= 12'b010000010110;
   27175: result <= 12'b010000010110;
   27176: result <= 12'b010000010110;
   27177: result <= 12'b010000010101;
   27178: result <= 12'b010000010101;
   27179: result <= 12'b010000010101;
   27180: result <= 12'b010000010101;
   27181: result <= 12'b010000010101;
   27182: result <= 12'b010000010101;
   27183: result <= 12'b010000010100;
   27184: result <= 12'b010000010100;
   27185: result <= 12'b010000010100;
   27186: result <= 12'b010000010100;
   27187: result <= 12'b010000010100;
   27188: result <= 12'b010000010100;
   27189: result <= 12'b010000010011;
   27190: result <= 12'b010000010011;
   27191: result <= 12'b010000010011;
   27192: result <= 12'b010000010011;
   27193: result <= 12'b010000010011;
   27194: result <= 12'b010000010011;
   27195: result <= 12'b010000010010;
   27196: result <= 12'b010000010010;
   27197: result <= 12'b010000010010;
   27198: result <= 12'b010000010010;
   27199: result <= 12'b010000010010;
   27200: result <= 12'b010000010010;
   27201: result <= 12'b010000010001;
   27202: result <= 12'b010000010001;
   27203: result <= 12'b010000010001;
   27204: result <= 12'b010000010001;
   27205: result <= 12'b010000010001;
   27206: result <= 12'b010000010001;
   27207: result <= 12'b010000010000;
   27208: result <= 12'b010000010000;
   27209: result <= 12'b010000010000;
   27210: result <= 12'b010000010000;
   27211: result <= 12'b010000010000;
   27212: result <= 12'b010000010000;
   27213: result <= 12'b010000001111;
   27214: result <= 12'b010000001111;
   27215: result <= 12'b010000001111;
   27216: result <= 12'b010000001111;
   27217: result <= 12'b010000001111;
   27218: result <= 12'b010000001111;
   27219: result <= 12'b010000001110;
   27220: result <= 12'b010000001110;
   27221: result <= 12'b010000001110;
   27222: result <= 12'b010000001110;
   27223: result <= 12'b010000001110;
   27224: result <= 12'b010000001110;
   27225: result <= 12'b010000001101;
   27226: result <= 12'b010000001101;
   27227: result <= 12'b010000001101;
   27228: result <= 12'b010000001101;
   27229: result <= 12'b010000001101;
   27230: result <= 12'b010000001101;
   27231: result <= 12'b010000001100;
   27232: result <= 12'b010000001100;
   27233: result <= 12'b010000001100;
   27234: result <= 12'b010000001100;
   27235: result <= 12'b010000001100;
   27236: result <= 12'b010000001011;
   27237: result <= 12'b010000001011;
   27238: result <= 12'b010000001011;
   27239: result <= 12'b010000001011;
   27240: result <= 12'b010000001011;
   27241: result <= 12'b010000001011;
   27242: result <= 12'b010000001010;
   27243: result <= 12'b010000001010;
   27244: result <= 12'b010000001010;
   27245: result <= 12'b010000001010;
   27246: result <= 12'b010000001010;
   27247: result <= 12'b010000001010;
   27248: result <= 12'b010000001001;
   27249: result <= 12'b010000001001;
   27250: result <= 12'b010000001001;
   27251: result <= 12'b010000001001;
   27252: result <= 12'b010000001001;
   27253: result <= 12'b010000001001;
   27254: result <= 12'b010000001000;
   27255: result <= 12'b010000001000;
   27256: result <= 12'b010000001000;
   27257: result <= 12'b010000001000;
   27258: result <= 12'b010000001000;
   27259: result <= 12'b010000001000;
   27260: result <= 12'b010000000111;
   27261: result <= 12'b010000000111;
   27262: result <= 12'b010000000111;
   27263: result <= 12'b010000000111;
   27264: result <= 12'b010000000111;
   27265: result <= 12'b010000000111;
   27266: result <= 12'b010000000110;
   27267: result <= 12'b010000000110;
   27268: result <= 12'b010000000110;
   27269: result <= 12'b010000000110;
   27270: result <= 12'b010000000110;
   27271: result <= 12'b010000000110;
   27272: result <= 12'b010000000101;
   27273: result <= 12'b010000000101;
   27274: result <= 12'b010000000101;
   27275: result <= 12'b010000000101;
   27276: result <= 12'b010000000101;
   27277: result <= 12'b010000000101;
   27278: result <= 12'b010000000100;
   27279: result <= 12'b010000000100;
   27280: result <= 12'b010000000100;
   27281: result <= 12'b010000000100;
   27282: result <= 12'b010000000100;
   27283: result <= 12'b010000000100;
   27284: result <= 12'b010000000011;
   27285: result <= 12'b010000000011;
   27286: result <= 12'b010000000011;
   27287: result <= 12'b010000000011;
   27288: result <= 12'b010000000011;
   27289: result <= 12'b010000000011;
   27290: result <= 12'b010000000010;
   27291: result <= 12'b010000000010;
   27292: result <= 12'b010000000010;
   27293: result <= 12'b010000000010;
   27294: result <= 12'b010000000010;
   27295: result <= 12'b010000000001;
   27296: result <= 12'b010000000001;
   27297: result <= 12'b010000000001;
   27298: result <= 12'b010000000001;
   27299: result <= 12'b010000000001;
   27300: result <= 12'b010000000001;
   27301: result <= 12'b010000000000;
   27302: result <= 12'b010000000000;
   27303: result <= 12'b010000000000;
   27304: result <= 12'b010000000000;
   27305: result <= 12'b010000000000;
   27306: result <= 12'b010000000000;
   27307: result <= 12'b001111111111;
   27308: result <= 12'b001111111111;
   27309: result <= 12'b001111111111;
   27310: result <= 12'b001111111111;
   27311: result <= 12'b001111111111;
   27312: result <= 12'b001111111111;
   27313: result <= 12'b001111111110;
   27314: result <= 12'b001111111110;
   27315: result <= 12'b001111111110;
   27316: result <= 12'b001111111110;
   27317: result <= 12'b001111111110;
   27318: result <= 12'b001111111110;
   27319: result <= 12'b001111111101;
   27320: result <= 12'b001111111101;
   27321: result <= 12'b001111111101;
   27322: result <= 12'b001111111101;
   27323: result <= 12'b001111111101;
   27324: result <= 12'b001111111101;
   27325: result <= 12'b001111111100;
   27326: result <= 12'b001111111100;
   27327: result <= 12'b001111111100;
   27328: result <= 12'b001111111100;
   27329: result <= 12'b001111111100;
   27330: result <= 12'b001111111100;
   27331: result <= 12'b001111111011;
   27332: result <= 12'b001111111011;
   27333: result <= 12'b001111111011;
   27334: result <= 12'b001111111011;
   27335: result <= 12'b001111111011;
   27336: result <= 12'b001111111011;
   27337: result <= 12'b001111111010;
   27338: result <= 12'b001111111010;
   27339: result <= 12'b001111111010;
   27340: result <= 12'b001111111010;
   27341: result <= 12'b001111111010;
   27342: result <= 12'b001111111001;
   27343: result <= 12'b001111111001;
   27344: result <= 12'b001111111001;
   27345: result <= 12'b001111111001;
   27346: result <= 12'b001111111001;
   27347: result <= 12'b001111111001;
   27348: result <= 12'b001111111000;
   27349: result <= 12'b001111111000;
   27350: result <= 12'b001111111000;
   27351: result <= 12'b001111111000;
   27352: result <= 12'b001111111000;
   27353: result <= 12'b001111111000;
   27354: result <= 12'b001111110111;
   27355: result <= 12'b001111110111;
   27356: result <= 12'b001111110111;
   27357: result <= 12'b001111110111;
   27358: result <= 12'b001111110111;
   27359: result <= 12'b001111110111;
   27360: result <= 12'b001111110110;
   27361: result <= 12'b001111110110;
   27362: result <= 12'b001111110110;
   27363: result <= 12'b001111110110;
   27364: result <= 12'b001111110110;
   27365: result <= 12'b001111110110;
   27366: result <= 12'b001111110101;
   27367: result <= 12'b001111110101;
   27368: result <= 12'b001111110101;
   27369: result <= 12'b001111110101;
   27370: result <= 12'b001111110101;
   27371: result <= 12'b001111110101;
   27372: result <= 12'b001111110100;
   27373: result <= 12'b001111110100;
   27374: result <= 12'b001111110100;
   27375: result <= 12'b001111110100;
   27376: result <= 12'b001111110100;
   27377: result <= 12'b001111110100;
   27378: result <= 12'b001111110011;
   27379: result <= 12'b001111110011;
   27380: result <= 12'b001111110011;
   27381: result <= 12'b001111110011;
   27382: result <= 12'b001111110011;
   27383: result <= 12'b001111110010;
   27384: result <= 12'b001111110010;
   27385: result <= 12'b001111110010;
   27386: result <= 12'b001111110010;
   27387: result <= 12'b001111110010;
   27388: result <= 12'b001111110010;
   27389: result <= 12'b001111110001;
   27390: result <= 12'b001111110001;
   27391: result <= 12'b001111110001;
   27392: result <= 12'b001111110001;
   27393: result <= 12'b001111110001;
   27394: result <= 12'b001111110001;
   27395: result <= 12'b001111110000;
   27396: result <= 12'b001111110000;
   27397: result <= 12'b001111110000;
   27398: result <= 12'b001111110000;
   27399: result <= 12'b001111110000;
   27400: result <= 12'b001111110000;
   27401: result <= 12'b001111101111;
   27402: result <= 12'b001111101111;
   27403: result <= 12'b001111101111;
   27404: result <= 12'b001111101111;
   27405: result <= 12'b001111101111;
   27406: result <= 12'b001111101111;
   27407: result <= 12'b001111101110;
   27408: result <= 12'b001111101110;
   27409: result <= 12'b001111101110;
   27410: result <= 12'b001111101110;
   27411: result <= 12'b001111101110;
   27412: result <= 12'b001111101110;
   27413: result <= 12'b001111101101;
   27414: result <= 12'b001111101101;
   27415: result <= 12'b001111101101;
   27416: result <= 12'b001111101101;
   27417: result <= 12'b001111101101;
   27418: result <= 12'b001111101101;
   27419: result <= 12'b001111101100;
   27420: result <= 12'b001111101100;
   27421: result <= 12'b001111101100;
   27422: result <= 12'b001111101100;
   27423: result <= 12'b001111101100;
   27424: result <= 12'b001111101011;
   27425: result <= 12'b001111101011;
   27426: result <= 12'b001111101011;
   27427: result <= 12'b001111101011;
   27428: result <= 12'b001111101011;
   27429: result <= 12'b001111101011;
   27430: result <= 12'b001111101010;
   27431: result <= 12'b001111101010;
   27432: result <= 12'b001111101010;
   27433: result <= 12'b001111101010;
   27434: result <= 12'b001111101010;
   27435: result <= 12'b001111101010;
   27436: result <= 12'b001111101001;
   27437: result <= 12'b001111101001;
   27438: result <= 12'b001111101001;
   27439: result <= 12'b001111101001;
   27440: result <= 12'b001111101001;
   27441: result <= 12'b001111101001;
   27442: result <= 12'b001111101000;
   27443: result <= 12'b001111101000;
   27444: result <= 12'b001111101000;
   27445: result <= 12'b001111101000;
   27446: result <= 12'b001111101000;
   27447: result <= 12'b001111101000;
   27448: result <= 12'b001111100111;
   27449: result <= 12'b001111100111;
   27450: result <= 12'b001111100111;
   27451: result <= 12'b001111100111;
   27452: result <= 12'b001111100111;
   27453: result <= 12'b001111100111;
   27454: result <= 12'b001111100110;
   27455: result <= 12'b001111100110;
   27456: result <= 12'b001111100110;
   27457: result <= 12'b001111100110;
   27458: result <= 12'b001111100110;
   27459: result <= 12'b001111100101;
   27460: result <= 12'b001111100101;
   27461: result <= 12'b001111100101;
   27462: result <= 12'b001111100101;
   27463: result <= 12'b001111100101;
   27464: result <= 12'b001111100101;
   27465: result <= 12'b001111100100;
   27466: result <= 12'b001111100100;
   27467: result <= 12'b001111100100;
   27468: result <= 12'b001111100100;
   27469: result <= 12'b001111100100;
   27470: result <= 12'b001111100100;
   27471: result <= 12'b001111100011;
   27472: result <= 12'b001111100011;
   27473: result <= 12'b001111100011;
   27474: result <= 12'b001111100011;
   27475: result <= 12'b001111100011;
   27476: result <= 12'b001111100011;
   27477: result <= 12'b001111100010;
   27478: result <= 12'b001111100010;
   27479: result <= 12'b001111100010;
   27480: result <= 12'b001111100010;
   27481: result <= 12'b001111100010;
   27482: result <= 12'b001111100010;
   27483: result <= 12'b001111100001;
   27484: result <= 12'b001111100001;
   27485: result <= 12'b001111100001;
   27486: result <= 12'b001111100001;
   27487: result <= 12'b001111100001;
   27488: result <= 12'b001111100001;
   27489: result <= 12'b001111100000;
   27490: result <= 12'b001111100000;
   27491: result <= 12'b001111100000;
   27492: result <= 12'b001111100000;
   27493: result <= 12'b001111100000;
   27494: result <= 12'b001111011111;
   27495: result <= 12'b001111011111;
   27496: result <= 12'b001111011111;
   27497: result <= 12'b001111011111;
   27498: result <= 12'b001111011111;
   27499: result <= 12'b001111011111;
   27500: result <= 12'b001111011110;
   27501: result <= 12'b001111011110;
   27502: result <= 12'b001111011110;
   27503: result <= 12'b001111011110;
   27504: result <= 12'b001111011110;
   27505: result <= 12'b001111011110;
   27506: result <= 12'b001111011101;
   27507: result <= 12'b001111011101;
   27508: result <= 12'b001111011101;
   27509: result <= 12'b001111011101;
   27510: result <= 12'b001111011101;
   27511: result <= 12'b001111011101;
   27512: result <= 12'b001111011100;
   27513: result <= 12'b001111011100;
   27514: result <= 12'b001111011100;
   27515: result <= 12'b001111011100;
   27516: result <= 12'b001111011100;
   27517: result <= 12'b001111011100;
   27518: result <= 12'b001111011011;
   27519: result <= 12'b001111011011;
   27520: result <= 12'b001111011011;
   27521: result <= 12'b001111011011;
   27522: result <= 12'b001111011011;
   27523: result <= 12'b001111011010;
   27524: result <= 12'b001111011010;
   27525: result <= 12'b001111011010;
   27526: result <= 12'b001111011010;
   27527: result <= 12'b001111011010;
   27528: result <= 12'b001111011010;
   27529: result <= 12'b001111011001;
   27530: result <= 12'b001111011001;
   27531: result <= 12'b001111011001;
   27532: result <= 12'b001111011001;
   27533: result <= 12'b001111011001;
   27534: result <= 12'b001111011001;
   27535: result <= 12'b001111011000;
   27536: result <= 12'b001111011000;
   27537: result <= 12'b001111011000;
   27538: result <= 12'b001111011000;
   27539: result <= 12'b001111011000;
   27540: result <= 12'b001111011000;
   27541: result <= 12'b001111010111;
   27542: result <= 12'b001111010111;
   27543: result <= 12'b001111010111;
   27544: result <= 12'b001111010111;
   27545: result <= 12'b001111010111;
   27546: result <= 12'b001111010111;
   27547: result <= 12'b001111010110;
   27548: result <= 12'b001111010110;
   27549: result <= 12'b001111010110;
   27550: result <= 12'b001111010110;
   27551: result <= 12'b001111010110;
   27552: result <= 12'b001111010110;
   27553: result <= 12'b001111010101;
   27554: result <= 12'b001111010101;
   27555: result <= 12'b001111010101;
   27556: result <= 12'b001111010101;
   27557: result <= 12'b001111010101;
   27558: result <= 12'b001111010100;
   27559: result <= 12'b001111010100;
   27560: result <= 12'b001111010100;
   27561: result <= 12'b001111010100;
   27562: result <= 12'b001111010100;
   27563: result <= 12'b001111010100;
   27564: result <= 12'b001111010011;
   27565: result <= 12'b001111010011;
   27566: result <= 12'b001111010011;
   27567: result <= 12'b001111010011;
   27568: result <= 12'b001111010011;
   27569: result <= 12'b001111010011;
   27570: result <= 12'b001111010010;
   27571: result <= 12'b001111010010;
   27572: result <= 12'b001111010010;
   27573: result <= 12'b001111010010;
   27574: result <= 12'b001111010010;
   27575: result <= 12'b001111010010;
   27576: result <= 12'b001111010001;
   27577: result <= 12'b001111010001;
   27578: result <= 12'b001111010001;
   27579: result <= 12'b001111010001;
   27580: result <= 12'b001111010001;
   27581: result <= 12'b001111010001;
   27582: result <= 12'b001111010000;
   27583: result <= 12'b001111010000;
   27584: result <= 12'b001111010000;
   27585: result <= 12'b001111010000;
   27586: result <= 12'b001111010000;
   27587: result <= 12'b001111001111;
   27588: result <= 12'b001111001111;
   27589: result <= 12'b001111001111;
   27590: result <= 12'b001111001111;
   27591: result <= 12'b001111001111;
   27592: result <= 12'b001111001111;
   27593: result <= 12'b001111001110;
   27594: result <= 12'b001111001110;
   27595: result <= 12'b001111001110;
   27596: result <= 12'b001111001110;
   27597: result <= 12'b001111001110;
   27598: result <= 12'b001111001110;
   27599: result <= 12'b001111001101;
   27600: result <= 12'b001111001101;
   27601: result <= 12'b001111001101;
   27602: result <= 12'b001111001101;
   27603: result <= 12'b001111001101;
   27604: result <= 12'b001111001101;
   27605: result <= 12'b001111001100;
   27606: result <= 12'b001111001100;
   27607: result <= 12'b001111001100;
   27608: result <= 12'b001111001100;
   27609: result <= 12'b001111001100;
   27610: result <= 12'b001111001011;
   27611: result <= 12'b001111001011;
   27612: result <= 12'b001111001011;
   27613: result <= 12'b001111001011;
   27614: result <= 12'b001111001011;
   27615: result <= 12'b001111001011;
   27616: result <= 12'b001111001010;
   27617: result <= 12'b001111001010;
   27618: result <= 12'b001111001010;
   27619: result <= 12'b001111001010;
   27620: result <= 12'b001111001010;
   27621: result <= 12'b001111001010;
   27622: result <= 12'b001111001001;
   27623: result <= 12'b001111001001;
   27624: result <= 12'b001111001001;
   27625: result <= 12'b001111001001;
   27626: result <= 12'b001111001001;
   27627: result <= 12'b001111001001;
   27628: result <= 12'b001111001000;
   27629: result <= 12'b001111001000;
   27630: result <= 12'b001111001000;
   27631: result <= 12'b001111001000;
   27632: result <= 12'b001111001000;
   27633: result <= 12'b001111001000;
   27634: result <= 12'b001111000111;
   27635: result <= 12'b001111000111;
   27636: result <= 12'b001111000111;
   27637: result <= 12'b001111000111;
   27638: result <= 12'b001111000111;
   27639: result <= 12'b001111000110;
   27640: result <= 12'b001111000110;
   27641: result <= 12'b001111000110;
   27642: result <= 12'b001111000110;
   27643: result <= 12'b001111000110;
   27644: result <= 12'b001111000110;
   27645: result <= 12'b001111000101;
   27646: result <= 12'b001111000101;
   27647: result <= 12'b001111000101;
   27648: result <= 12'b001111000101;
   27649: result <= 12'b001111000101;
   27650: result <= 12'b001111000101;
   27651: result <= 12'b001111000100;
   27652: result <= 12'b001111000100;
   27653: result <= 12'b001111000100;
   27654: result <= 12'b001111000100;
   27655: result <= 12'b001111000100;
   27656: result <= 12'b001111000100;
   27657: result <= 12'b001111000011;
   27658: result <= 12'b001111000011;
   27659: result <= 12'b001111000011;
   27660: result <= 12'b001111000011;
   27661: result <= 12'b001111000011;
   27662: result <= 12'b001111000010;
   27663: result <= 12'b001111000010;
   27664: result <= 12'b001111000010;
   27665: result <= 12'b001111000010;
   27666: result <= 12'b001111000010;
   27667: result <= 12'b001111000010;
   27668: result <= 12'b001111000001;
   27669: result <= 12'b001111000001;
   27670: result <= 12'b001111000001;
   27671: result <= 12'b001111000001;
   27672: result <= 12'b001111000001;
   27673: result <= 12'b001111000001;
   27674: result <= 12'b001111000000;
   27675: result <= 12'b001111000000;
   27676: result <= 12'b001111000000;
   27677: result <= 12'b001111000000;
   27678: result <= 12'b001111000000;
   27679: result <= 12'b001111000000;
   27680: result <= 12'b001110111111;
   27681: result <= 12'b001110111111;
   27682: result <= 12'b001110111111;
   27683: result <= 12'b001110111111;
   27684: result <= 12'b001110111111;
   27685: result <= 12'b001110111111;
   27686: result <= 12'b001110111110;
   27687: result <= 12'b001110111110;
   27688: result <= 12'b001110111110;
   27689: result <= 12'b001110111110;
   27690: result <= 12'b001110111110;
   27691: result <= 12'b001110111101;
   27692: result <= 12'b001110111101;
   27693: result <= 12'b001110111101;
   27694: result <= 12'b001110111101;
   27695: result <= 12'b001110111101;
   27696: result <= 12'b001110111101;
   27697: result <= 12'b001110111100;
   27698: result <= 12'b001110111100;
   27699: result <= 12'b001110111100;
   27700: result <= 12'b001110111100;
   27701: result <= 12'b001110111100;
   27702: result <= 12'b001110111100;
   27703: result <= 12'b001110111011;
   27704: result <= 12'b001110111011;
   27705: result <= 12'b001110111011;
   27706: result <= 12'b001110111011;
   27707: result <= 12'b001110111011;
   27708: result <= 12'b001110111011;
   27709: result <= 12'b001110111010;
   27710: result <= 12'b001110111010;
   27711: result <= 12'b001110111010;
   27712: result <= 12'b001110111010;
   27713: result <= 12'b001110111010;
   27714: result <= 12'b001110111001;
   27715: result <= 12'b001110111001;
   27716: result <= 12'b001110111001;
   27717: result <= 12'b001110111001;
   27718: result <= 12'b001110111001;
   27719: result <= 12'b001110111001;
   27720: result <= 12'b001110111000;
   27721: result <= 12'b001110111000;
   27722: result <= 12'b001110111000;
   27723: result <= 12'b001110111000;
   27724: result <= 12'b001110111000;
   27725: result <= 12'b001110111000;
   27726: result <= 12'b001110110111;
   27727: result <= 12'b001110110111;
   27728: result <= 12'b001110110111;
   27729: result <= 12'b001110110111;
   27730: result <= 12'b001110110111;
   27731: result <= 12'b001110110111;
   27732: result <= 12'b001110110110;
   27733: result <= 12'b001110110110;
   27734: result <= 12'b001110110110;
   27735: result <= 12'b001110110110;
   27736: result <= 12'b001110110110;
   27737: result <= 12'b001110110101;
   27738: result <= 12'b001110110101;
   27739: result <= 12'b001110110101;
   27740: result <= 12'b001110110101;
   27741: result <= 12'b001110110101;
   27742: result <= 12'b001110110101;
   27743: result <= 12'b001110110100;
   27744: result <= 12'b001110110100;
   27745: result <= 12'b001110110100;
   27746: result <= 12'b001110110100;
   27747: result <= 12'b001110110100;
   27748: result <= 12'b001110110100;
   27749: result <= 12'b001110110011;
   27750: result <= 12'b001110110011;
   27751: result <= 12'b001110110011;
   27752: result <= 12'b001110110011;
   27753: result <= 12'b001110110011;
   27754: result <= 12'b001110110011;
   27755: result <= 12'b001110110010;
   27756: result <= 12'b001110110010;
   27757: result <= 12'b001110110010;
   27758: result <= 12'b001110110010;
   27759: result <= 12'b001110110010;
   27760: result <= 12'b001110110001;
   27761: result <= 12'b001110110001;
   27762: result <= 12'b001110110001;
   27763: result <= 12'b001110110001;
   27764: result <= 12'b001110110001;
   27765: result <= 12'b001110110001;
   27766: result <= 12'b001110110000;
   27767: result <= 12'b001110110000;
   27768: result <= 12'b001110110000;
   27769: result <= 12'b001110110000;
   27770: result <= 12'b001110110000;
   27771: result <= 12'b001110110000;
   27772: result <= 12'b001110101111;
   27773: result <= 12'b001110101111;
   27774: result <= 12'b001110101111;
   27775: result <= 12'b001110101111;
   27776: result <= 12'b001110101111;
   27777: result <= 12'b001110101111;
   27778: result <= 12'b001110101110;
   27779: result <= 12'b001110101110;
   27780: result <= 12'b001110101110;
   27781: result <= 12'b001110101110;
   27782: result <= 12'b001110101110;
   27783: result <= 12'b001110101101;
   27784: result <= 12'b001110101101;
   27785: result <= 12'b001110101101;
   27786: result <= 12'b001110101101;
   27787: result <= 12'b001110101101;
   27788: result <= 12'b001110101101;
   27789: result <= 12'b001110101100;
   27790: result <= 12'b001110101100;
   27791: result <= 12'b001110101100;
   27792: result <= 12'b001110101100;
   27793: result <= 12'b001110101100;
   27794: result <= 12'b001110101100;
   27795: result <= 12'b001110101011;
   27796: result <= 12'b001110101011;
   27797: result <= 12'b001110101011;
   27798: result <= 12'b001110101011;
   27799: result <= 12'b001110101011;
   27800: result <= 12'b001110101010;
   27801: result <= 12'b001110101010;
   27802: result <= 12'b001110101010;
   27803: result <= 12'b001110101010;
   27804: result <= 12'b001110101010;
   27805: result <= 12'b001110101010;
   27806: result <= 12'b001110101001;
   27807: result <= 12'b001110101001;
   27808: result <= 12'b001110101001;
   27809: result <= 12'b001110101001;
   27810: result <= 12'b001110101001;
   27811: result <= 12'b001110101001;
   27812: result <= 12'b001110101000;
   27813: result <= 12'b001110101000;
   27814: result <= 12'b001110101000;
   27815: result <= 12'b001110101000;
   27816: result <= 12'b001110101000;
   27817: result <= 12'b001110101000;
   27818: result <= 12'b001110100111;
   27819: result <= 12'b001110100111;
   27820: result <= 12'b001110100111;
   27821: result <= 12'b001110100111;
   27822: result <= 12'b001110100111;
   27823: result <= 12'b001110100110;
   27824: result <= 12'b001110100110;
   27825: result <= 12'b001110100110;
   27826: result <= 12'b001110100110;
   27827: result <= 12'b001110100110;
   27828: result <= 12'b001110100110;
   27829: result <= 12'b001110100101;
   27830: result <= 12'b001110100101;
   27831: result <= 12'b001110100101;
   27832: result <= 12'b001110100101;
   27833: result <= 12'b001110100101;
   27834: result <= 12'b001110100101;
   27835: result <= 12'b001110100100;
   27836: result <= 12'b001110100100;
   27837: result <= 12'b001110100100;
   27838: result <= 12'b001110100100;
   27839: result <= 12'b001110100100;
   27840: result <= 12'b001110100100;
   27841: result <= 12'b001110100011;
   27842: result <= 12'b001110100011;
   27843: result <= 12'b001110100011;
   27844: result <= 12'b001110100011;
   27845: result <= 12'b001110100011;
   27846: result <= 12'b001110100010;
   27847: result <= 12'b001110100010;
   27848: result <= 12'b001110100010;
   27849: result <= 12'b001110100010;
   27850: result <= 12'b001110100010;
   27851: result <= 12'b001110100010;
   27852: result <= 12'b001110100001;
   27853: result <= 12'b001110100001;
   27854: result <= 12'b001110100001;
   27855: result <= 12'b001110100001;
   27856: result <= 12'b001110100001;
   27857: result <= 12'b001110100001;
   27858: result <= 12'b001110100000;
   27859: result <= 12'b001110100000;
   27860: result <= 12'b001110100000;
   27861: result <= 12'b001110100000;
   27862: result <= 12'b001110100000;
   27863: result <= 12'b001110011111;
   27864: result <= 12'b001110011111;
   27865: result <= 12'b001110011111;
   27866: result <= 12'b001110011111;
   27867: result <= 12'b001110011111;
   27868: result <= 12'b001110011111;
   27869: result <= 12'b001110011110;
   27870: result <= 12'b001110011110;
   27871: result <= 12'b001110011110;
   27872: result <= 12'b001110011110;
   27873: result <= 12'b001110011110;
   27874: result <= 12'b001110011110;
   27875: result <= 12'b001110011101;
   27876: result <= 12'b001110011101;
   27877: result <= 12'b001110011101;
   27878: result <= 12'b001110011101;
   27879: result <= 12'b001110011101;
   27880: result <= 12'b001110011101;
   27881: result <= 12'b001110011100;
   27882: result <= 12'b001110011100;
   27883: result <= 12'b001110011100;
   27884: result <= 12'b001110011100;
   27885: result <= 12'b001110011100;
   27886: result <= 12'b001110011011;
   27887: result <= 12'b001110011011;
   27888: result <= 12'b001110011011;
   27889: result <= 12'b001110011011;
   27890: result <= 12'b001110011011;
   27891: result <= 12'b001110011011;
   27892: result <= 12'b001110011010;
   27893: result <= 12'b001110011010;
   27894: result <= 12'b001110011010;
   27895: result <= 12'b001110011010;
   27896: result <= 12'b001110011010;
   27897: result <= 12'b001110011010;
   27898: result <= 12'b001110011001;
   27899: result <= 12'b001110011001;
   27900: result <= 12'b001110011001;
   27901: result <= 12'b001110011001;
   27902: result <= 12'b001110011001;
   27903: result <= 12'b001110011000;
   27904: result <= 12'b001110011000;
   27905: result <= 12'b001110011000;
   27906: result <= 12'b001110011000;
   27907: result <= 12'b001110011000;
   27908: result <= 12'b001110011000;
   27909: result <= 12'b001110010111;
   27910: result <= 12'b001110010111;
   27911: result <= 12'b001110010111;
   27912: result <= 12'b001110010111;
   27913: result <= 12'b001110010111;
   27914: result <= 12'b001110010111;
   27915: result <= 12'b001110010110;
   27916: result <= 12'b001110010110;
   27917: result <= 12'b001110010110;
   27918: result <= 12'b001110010110;
   27919: result <= 12'b001110010110;
   27920: result <= 12'b001110010101;
   27921: result <= 12'b001110010101;
   27922: result <= 12'b001110010101;
   27923: result <= 12'b001110010101;
   27924: result <= 12'b001110010101;
   27925: result <= 12'b001110010101;
   27926: result <= 12'b001110010100;
   27927: result <= 12'b001110010100;
   27928: result <= 12'b001110010100;
   27929: result <= 12'b001110010100;
   27930: result <= 12'b001110010100;
   27931: result <= 12'b001110010100;
   27932: result <= 12'b001110010011;
   27933: result <= 12'b001110010011;
   27934: result <= 12'b001110010011;
   27935: result <= 12'b001110010011;
   27936: result <= 12'b001110010011;
   27937: result <= 12'b001110010011;
   27938: result <= 12'b001110010010;
   27939: result <= 12'b001110010010;
   27940: result <= 12'b001110010010;
   27941: result <= 12'b001110010010;
   27942: result <= 12'b001110010010;
   27943: result <= 12'b001110010001;
   27944: result <= 12'b001110010001;
   27945: result <= 12'b001110010001;
   27946: result <= 12'b001110010001;
   27947: result <= 12'b001110010001;
   27948: result <= 12'b001110010001;
   27949: result <= 12'b001110010000;
   27950: result <= 12'b001110010000;
   27951: result <= 12'b001110010000;
   27952: result <= 12'b001110010000;
   27953: result <= 12'b001110010000;
   27954: result <= 12'b001110010000;
   27955: result <= 12'b001110001111;
   27956: result <= 12'b001110001111;
   27957: result <= 12'b001110001111;
   27958: result <= 12'b001110001111;
   27959: result <= 12'b001110001111;
   27960: result <= 12'b001110001110;
   27961: result <= 12'b001110001110;
   27962: result <= 12'b001110001110;
   27963: result <= 12'b001110001110;
   27964: result <= 12'b001110001110;
   27965: result <= 12'b001110001110;
   27966: result <= 12'b001110001101;
   27967: result <= 12'b001110001101;
   27968: result <= 12'b001110001101;
   27969: result <= 12'b001110001101;
   27970: result <= 12'b001110001101;
   27971: result <= 12'b001110001101;
   27972: result <= 12'b001110001100;
   27973: result <= 12'b001110001100;
   27974: result <= 12'b001110001100;
   27975: result <= 12'b001110001100;
   27976: result <= 12'b001110001100;
   27977: result <= 12'b001110001011;
   27978: result <= 12'b001110001011;
   27979: result <= 12'b001110001011;
   27980: result <= 12'b001110001011;
   27981: result <= 12'b001110001011;
   27982: result <= 12'b001110001011;
   27983: result <= 12'b001110001010;
   27984: result <= 12'b001110001010;
   27985: result <= 12'b001110001010;
   27986: result <= 12'b001110001010;
   27987: result <= 12'b001110001010;
   27988: result <= 12'b001110001010;
   27989: result <= 12'b001110001001;
   27990: result <= 12'b001110001001;
   27991: result <= 12'b001110001001;
   27992: result <= 12'b001110001001;
   27993: result <= 12'b001110001001;
   27994: result <= 12'b001110001000;
   27995: result <= 12'b001110001000;
   27996: result <= 12'b001110001000;
   27997: result <= 12'b001110001000;
   27998: result <= 12'b001110001000;
   27999: result <= 12'b001110001000;
   28000: result <= 12'b001110000111;
   28001: result <= 12'b001110000111;
   28002: result <= 12'b001110000111;
   28003: result <= 12'b001110000111;
   28004: result <= 12'b001110000111;
   28005: result <= 12'b001110000111;
   28006: result <= 12'b001110000110;
   28007: result <= 12'b001110000110;
   28008: result <= 12'b001110000110;
   28009: result <= 12'b001110000110;
   28010: result <= 12'b001110000110;
   28011: result <= 12'b001110000101;
   28012: result <= 12'b001110000101;
   28013: result <= 12'b001110000101;
   28014: result <= 12'b001110000101;
   28015: result <= 12'b001110000101;
   28016: result <= 12'b001110000101;
   28017: result <= 12'b001110000100;
   28018: result <= 12'b001110000100;
   28019: result <= 12'b001110000100;
   28020: result <= 12'b001110000100;
   28021: result <= 12'b001110000100;
   28022: result <= 12'b001110000100;
   28023: result <= 12'b001110000011;
   28024: result <= 12'b001110000011;
   28025: result <= 12'b001110000011;
   28026: result <= 12'b001110000011;
   28027: result <= 12'b001110000011;
   28028: result <= 12'b001110000010;
   28029: result <= 12'b001110000010;
   28030: result <= 12'b001110000010;
   28031: result <= 12'b001110000010;
   28032: result <= 12'b001110000010;
   28033: result <= 12'b001110000010;
   28034: result <= 12'b001110000001;
   28035: result <= 12'b001110000001;
   28036: result <= 12'b001110000001;
   28037: result <= 12'b001110000001;
   28038: result <= 12'b001110000001;
   28039: result <= 12'b001110000001;
   28040: result <= 12'b001110000000;
   28041: result <= 12'b001110000000;
   28042: result <= 12'b001110000000;
   28043: result <= 12'b001110000000;
   28044: result <= 12'b001110000000;
   28045: result <= 12'b001101111111;
   28046: result <= 12'b001101111111;
   28047: result <= 12'b001101111111;
   28048: result <= 12'b001101111111;
   28049: result <= 12'b001101111111;
   28050: result <= 12'b001101111111;
   28051: result <= 12'b001101111110;
   28052: result <= 12'b001101111110;
   28053: result <= 12'b001101111110;
   28054: result <= 12'b001101111110;
   28055: result <= 12'b001101111110;
   28056: result <= 12'b001101111110;
   28057: result <= 12'b001101111101;
   28058: result <= 12'b001101111101;
   28059: result <= 12'b001101111101;
   28060: result <= 12'b001101111101;
   28061: result <= 12'b001101111101;
   28062: result <= 12'b001101111100;
   28063: result <= 12'b001101111100;
   28064: result <= 12'b001101111100;
   28065: result <= 12'b001101111100;
   28066: result <= 12'b001101111100;
   28067: result <= 12'b001101111100;
   28068: result <= 12'b001101111011;
   28069: result <= 12'b001101111011;
   28070: result <= 12'b001101111011;
   28071: result <= 12'b001101111011;
   28072: result <= 12'b001101111011;
   28073: result <= 12'b001101111011;
   28074: result <= 12'b001101111010;
   28075: result <= 12'b001101111010;
   28076: result <= 12'b001101111010;
   28077: result <= 12'b001101111010;
   28078: result <= 12'b001101111010;
   28079: result <= 12'b001101111001;
   28080: result <= 12'b001101111001;
   28081: result <= 12'b001101111001;
   28082: result <= 12'b001101111001;
   28083: result <= 12'b001101111001;
   28084: result <= 12'b001101111001;
   28085: result <= 12'b001101111000;
   28086: result <= 12'b001101111000;
   28087: result <= 12'b001101111000;
   28088: result <= 12'b001101111000;
   28089: result <= 12'b001101111000;
   28090: result <= 12'b001101111000;
   28091: result <= 12'b001101110111;
   28092: result <= 12'b001101110111;
   28093: result <= 12'b001101110111;
   28094: result <= 12'b001101110111;
   28095: result <= 12'b001101110111;
   28096: result <= 12'b001101110110;
   28097: result <= 12'b001101110110;
   28098: result <= 12'b001101110110;
   28099: result <= 12'b001101110110;
   28100: result <= 12'b001101110110;
   28101: result <= 12'b001101110110;
   28102: result <= 12'b001101110101;
   28103: result <= 12'b001101110101;
   28104: result <= 12'b001101110101;
   28105: result <= 12'b001101110101;
   28106: result <= 12'b001101110101;
   28107: result <= 12'b001101110101;
   28108: result <= 12'b001101110100;
   28109: result <= 12'b001101110100;
   28110: result <= 12'b001101110100;
   28111: result <= 12'b001101110100;
   28112: result <= 12'b001101110100;
   28113: result <= 12'b001101110011;
   28114: result <= 12'b001101110011;
   28115: result <= 12'b001101110011;
   28116: result <= 12'b001101110011;
   28117: result <= 12'b001101110011;
   28118: result <= 12'b001101110011;
   28119: result <= 12'b001101110010;
   28120: result <= 12'b001101110010;
   28121: result <= 12'b001101110010;
   28122: result <= 12'b001101110010;
   28123: result <= 12'b001101110010;
   28124: result <= 12'b001101110010;
   28125: result <= 12'b001101110001;
   28126: result <= 12'b001101110001;
   28127: result <= 12'b001101110001;
   28128: result <= 12'b001101110001;
   28129: result <= 12'b001101110001;
   28130: result <= 12'b001101110000;
   28131: result <= 12'b001101110000;
   28132: result <= 12'b001101110000;
   28133: result <= 12'b001101110000;
   28134: result <= 12'b001101110000;
   28135: result <= 12'b001101110000;
   28136: result <= 12'b001101101111;
   28137: result <= 12'b001101101111;
   28138: result <= 12'b001101101111;
   28139: result <= 12'b001101101111;
   28140: result <= 12'b001101101111;
   28141: result <= 12'b001101101111;
   28142: result <= 12'b001101101110;
   28143: result <= 12'b001101101110;
   28144: result <= 12'b001101101110;
   28145: result <= 12'b001101101110;
   28146: result <= 12'b001101101110;
   28147: result <= 12'b001101101101;
   28148: result <= 12'b001101101101;
   28149: result <= 12'b001101101101;
   28150: result <= 12'b001101101101;
   28151: result <= 12'b001101101101;
   28152: result <= 12'b001101101101;
   28153: result <= 12'b001101101100;
   28154: result <= 12'b001101101100;
   28155: result <= 12'b001101101100;
   28156: result <= 12'b001101101100;
   28157: result <= 12'b001101101100;
   28158: result <= 12'b001101101011;
   28159: result <= 12'b001101101011;
   28160: result <= 12'b001101101011;
   28161: result <= 12'b001101101011;
   28162: result <= 12'b001101101011;
   28163: result <= 12'b001101101011;
   28164: result <= 12'b001101101010;
   28165: result <= 12'b001101101010;
   28166: result <= 12'b001101101010;
   28167: result <= 12'b001101101010;
   28168: result <= 12'b001101101010;
   28169: result <= 12'b001101101010;
   28170: result <= 12'b001101101001;
   28171: result <= 12'b001101101001;
   28172: result <= 12'b001101101001;
   28173: result <= 12'b001101101001;
   28174: result <= 12'b001101101001;
   28175: result <= 12'b001101101000;
   28176: result <= 12'b001101101000;
   28177: result <= 12'b001101101000;
   28178: result <= 12'b001101101000;
   28179: result <= 12'b001101101000;
   28180: result <= 12'b001101101000;
   28181: result <= 12'b001101100111;
   28182: result <= 12'b001101100111;
   28183: result <= 12'b001101100111;
   28184: result <= 12'b001101100111;
   28185: result <= 12'b001101100111;
   28186: result <= 12'b001101100111;
   28187: result <= 12'b001101100110;
   28188: result <= 12'b001101100110;
   28189: result <= 12'b001101100110;
   28190: result <= 12'b001101100110;
   28191: result <= 12'b001101100110;
   28192: result <= 12'b001101100101;
   28193: result <= 12'b001101100101;
   28194: result <= 12'b001101100101;
   28195: result <= 12'b001101100101;
   28196: result <= 12'b001101100101;
   28197: result <= 12'b001101100101;
   28198: result <= 12'b001101100100;
   28199: result <= 12'b001101100100;
   28200: result <= 12'b001101100100;
   28201: result <= 12'b001101100100;
   28202: result <= 12'b001101100100;
   28203: result <= 12'b001101100011;
   28204: result <= 12'b001101100011;
   28205: result <= 12'b001101100011;
   28206: result <= 12'b001101100011;
   28207: result <= 12'b001101100011;
   28208: result <= 12'b001101100011;
   28209: result <= 12'b001101100010;
   28210: result <= 12'b001101100010;
   28211: result <= 12'b001101100010;
   28212: result <= 12'b001101100010;
   28213: result <= 12'b001101100010;
   28214: result <= 12'b001101100010;
   28215: result <= 12'b001101100001;
   28216: result <= 12'b001101100001;
   28217: result <= 12'b001101100001;
   28218: result <= 12'b001101100001;
   28219: result <= 12'b001101100001;
   28220: result <= 12'b001101100000;
   28221: result <= 12'b001101100000;
   28222: result <= 12'b001101100000;
   28223: result <= 12'b001101100000;
   28224: result <= 12'b001101100000;
   28225: result <= 12'b001101100000;
   28226: result <= 12'b001101011111;
   28227: result <= 12'b001101011111;
   28228: result <= 12'b001101011111;
   28229: result <= 12'b001101011111;
   28230: result <= 12'b001101011111;
   28231: result <= 12'b001101011111;
   28232: result <= 12'b001101011110;
   28233: result <= 12'b001101011110;
   28234: result <= 12'b001101011110;
   28235: result <= 12'b001101011110;
   28236: result <= 12'b001101011110;
   28237: result <= 12'b001101011101;
   28238: result <= 12'b001101011101;
   28239: result <= 12'b001101011101;
   28240: result <= 12'b001101011101;
   28241: result <= 12'b001101011101;
   28242: result <= 12'b001101011101;
   28243: result <= 12'b001101011100;
   28244: result <= 12'b001101011100;
   28245: result <= 12'b001101011100;
   28246: result <= 12'b001101011100;
   28247: result <= 12'b001101011100;
   28248: result <= 12'b001101011011;
   28249: result <= 12'b001101011011;
   28250: result <= 12'b001101011011;
   28251: result <= 12'b001101011011;
   28252: result <= 12'b001101011011;
   28253: result <= 12'b001101011011;
   28254: result <= 12'b001101011010;
   28255: result <= 12'b001101011010;
   28256: result <= 12'b001101011010;
   28257: result <= 12'b001101011010;
   28258: result <= 12'b001101011010;
   28259: result <= 12'b001101011010;
   28260: result <= 12'b001101011001;
   28261: result <= 12'b001101011001;
   28262: result <= 12'b001101011001;
   28263: result <= 12'b001101011001;
   28264: result <= 12'b001101011001;
   28265: result <= 12'b001101011000;
   28266: result <= 12'b001101011000;
   28267: result <= 12'b001101011000;
   28268: result <= 12'b001101011000;
   28269: result <= 12'b001101011000;
   28270: result <= 12'b001101011000;
   28271: result <= 12'b001101010111;
   28272: result <= 12'b001101010111;
   28273: result <= 12'b001101010111;
   28274: result <= 12'b001101010111;
   28275: result <= 12'b001101010111;
   28276: result <= 12'b001101010110;
   28277: result <= 12'b001101010110;
   28278: result <= 12'b001101010110;
   28279: result <= 12'b001101010110;
   28280: result <= 12'b001101010110;
   28281: result <= 12'b001101010110;
   28282: result <= 12'b001101010101;
   28283: result <= 12'b001101010101;
   28284: result <= 12'b001101010101;
   28285: result <= 12'b001101010101;
   28286: result <= 12'b001101010101;
   28287: result <= 12'b001101010101;
   28288: result <= 12'b001101010100;
   28289: result <= 12'b001101010100;
   28290: result <= 12'b001101010100;
   28291: result <= 12'b001101010100;
   28292: result <= 12'b001101010100;
   28293: result <= 12'b001101010011;
   28294: result <= 12'b001101010011;
   28295: result <= 12'b001101010011;
   28296: result <= 12'b001101010011;
   28297: result <= 12'b001101010011;
   28298: result <= 12'b001101010011;
   28299: result <= 12'b001101010010;
   28300: result <= 12'b001101010010;
   28301: result <= 12'b001101010010;
   28302: result <= 12'b001101010010;
   28303: result <= 12'b001101010010;
   28304: result <= 12'b001101010001;
   28305: result <= 12'b001101010001;
   28306: result <= 12'b001101010001;
   28307: result <= 12'b001101010001;
   28308: result <= 12'b001101010001;
   28309: result <= 12'b001101010001;
   28310: result <= 12'b001101010000;
   28311: result <= 12'b001101010000;
   28312: result <= 12'b001101010000;
   28313: result <= 12'b001101010000;
   28314: result <= 12'b001101010000;
   28315: result <= 12'b001101010000;
   28316: result <= 12'b001101001111;
   28317: result <= 12'b001101001111;
   28318: result <= 12'b001101001111;
   28319: result <= 12'b001101001111;
   28320: result <= 12'b001101001111;
   28321: result <= 12'b001101001110;
   28322: result <= 12'b001101001110;
   28323: result <= 12'b001101001110;
   28324: result <= 12'b001101001110;
   28325: result <= 12'b001101001110;
   28326: result <= 12'b001101001110;
   28327: result <= 12'b001101001101;
   28328: result <= 12'b001101001101;
   28329: result <= 12'b001101001101;
   28330: result <= 12'b001101001101;
   28331: result <= 12'b001101001101;
   28332: result <= 12'b001101001100;
   28333: result <= 12'b001101001100;
   28334: result <= 12'b001101001100;
   28335: result <= 12'b001101001100;
   28336: result <= 12'b001101001100;
   28337: result <= 12'b001101001100;
   28338: result <= 12'b001101001011;
   28339: result <= 12'b001101001011;
   28340: result <= 12'b001101001011;
   28341: result <= 12'b001101001011;
   28342: result <= 12'b001101001011;
   28343: result <= 12'b001101001011;
   28344: result <= 12'b001101001010;
   28345: result <= 12'b001101001010;
   28346: result <= 12'b001101001010;
   28347: result <= 12'b001101001010;
   28348: result <= 12'b001101001010;
   28349: result <= 12'b001101001001;
   28350: result <= 12'b001101001001;
   28351: result <= 12'b001101001001;
   28352: result <= 12'b001101001001;
   28353: result <= 12'b001101001001;
   28354: result <= 12'b001101001001;
   28355: result <= 12'b001101001000;
   28356: result <= 12'b001101001000;
   28357: result <= 12'b001101001000;
   28358: result <= 12'b001101001000;
   28359: result <= 12'b001101001000;
   28360: result <= 12'b001101000111;
   28361: result <= 12'b001101000111;
   28362: result <= 12'b001101000111;
   28363: result <= 12'b001101000111;
   28364: result <= 12'b001101000111;
   28365: result <= 12'b001101000111;
   28366: result <= 12'b001101000110;
   28367: result <= 12'b001101000110;
   28368: result <= 12'b001101000110;
   28369: result <= 12'b001101000110;
   28370: result <= 12'b001101000110;
   28371: result <= 12'b001101000110;
   28372: result <= 12'b001101000101;
   28373: result <= 12'b001101000101;
   28374: result <= 12'b001101000101;
   28375: result <= 12'b001101000101;
   28376: result <= 12'b001101000101;
   28377: result <= 12'b001101000100;
   28378: result <= 12'b001101000100;
   28379: result <= 12'b001101000100;
   28380: result <= 12'b001101000100;
   28381: result <= 12'b001101000100;
   28382: result <= 12'b001101000100;
   28383: result <= 12'b001101000011;
   28384: result <= 12'b001101000011;
   28385: result <= 12'b001101000011;
   28386: result <= 12'b001101000011;
   28387: result <= 12'b001101000011;
   28388: result <= 12'b001101000010;
   28389: result <= 12'b001101000010;
   28390: result <= 12'b001101000010;
   28391: result <= 12'b001101000010;
   28392: result <= 12'b001101000010;
   28393: result <= 12'b001101000010;
   28394: result <= 12'b001101000001;
   28395: result <= 12'b001101000001;
   28396: result <= 12'b001101000001;
   28397: result <= 12'b001101000001;
   28398: result <= 12'b001101000001;
   28399: result <= 12'b001101000000;
   28400: result <= 12'b001101000000;
   28401: result <= 12'b001101000000;
   28402: result <= 12'b001101000000;
   28403: result <= 12'b001101000000;
   28404: result <= 12'b001101000000;
   28405: result <= 12'b001100111111;
   28406: result <= 12'b001100111111;
   28407: result <= 12'b001100111111;
   28408: result <= 12'b001100111111;
   28409: result <= 12'b001100111111;
   28410: result <= 12'b001100111111;
   28411: result <= 12'b001100111110;
   28412: result <= 12'b001100111110;
   28413: result <= 12'b001100111110;
   28414: result <= 12'b001100111110;
   28415: result <= 12'b001100111110;
   28416: result <= 12'b001100111101;
   28417: result <= 12'b001100111101;
   28418: result <= 12'b001100111101;
   28419: result <= 12'b001100111101;
   28420: result <= 12'b001100111101;
   28421: result <= 12'b001100111101;
   28422: result <= 12'b001100111100;
   28423: result <= 12'b001100111100;
   28424: result <= 12'b001100111100;
   28425: result <= 12'b001100111100;
   28426: result <= 12'b001100111100;
   28427: result <= 12'b001100111011;
   28428: result <= 12'b001100111011;
   28429: result <= 12'b001100111011;
   28430: result <= 12'b001100111011;
   28431: result <= 12'b001100111011;
   28432: result <= 12'b001100111011;
   28433: result <= 12'b001100111010;
   28434: result <= 12'b001100111010;
   28435: result <= 12'b001100111010;
   28436: result <= 12'b001100111010;
   28437: result <= 12'b001100111010;
   28438: result <= 12'b001100111001;
   28439: result <= 12'b001100111001;
   28440: result <= 12'b001100111001;
   28441: result <= 12'b001100111001;
   28442: result <= 12'b001100111001;
   28443: result <= 12'b001100111001;
   28444: result <= 12'b001100111000;
   28445: result <= 12'b001100111000;
   28446: result <= 12'b001100111000;
   28447: result <= 12'b001100111000;
   28448: result <= 12'b001100111000;
   28449: result <= 12'b001100111000;
   28450: result <= 12'b001100110111;
   28451: result <= 12'b001100110111;
   28452: result <= 12'b001100110111;
   28453: result <= 12'b001100110111;
   28454: result <= 12'b001100110111;
   28455: result <= 12'b001100110110;
   28456: result <= 12'b001100110110;
   28457: result <= 12'b001100110110;
   28458: result <= 12'b001100110110;
   28459: result <= 12'b001100110110;
   28460: result <= 12'b001100110110;
   28461: result <= 12'b001100110101;
   28462: result <= 12'b001100110101;
   28463: result <= 12'b001100110101;
   28464: result <= 12'b001100110101;
   28465: result <= 12'b001100110101;
   28466: result <= 12'b001100110100;
   28467: result <= 12'b001100110100;
   28468: result <= 12'b001100110100;
   28469: result <= 12'b001100110100;
   28470: result <= 12'b001100110100;
   28471: result <= 12'b001100110100;
   28472: result <= 12'b001100110011;
   28473: result <= 12'b001100110011;
   28474: result <= 12'b001100110011;
   28475: result <= 12'b001100110011;
   28476: result <= 12'b001100110011;
   28477: result <= 12'b001100110010;
   28478: result <= 12'b001100110010;
   28479: result <= 12'b001100110010;
   28480: result <= 12'b001100110010;
   28481: result <= 12'b001100110010;
   28482: result <= 12'b001100110010;
   28483: result <= 12'b001100110001;
   28484: result <= 12'b001100110001;
   28485: result <= 12'b001100110001;
   28486: result <= 12'b001100110001;
   28487: result <= 12'b001100110001;
   28488: result <= 12'b001100110000;
   28489: result <= 12'b001100110000;
   28490: result <= 12'b001100110000;
   28491: result <= 12'b001100110000;
   28492: result <= 12'b001100110000;
   28493: result <= 12'b001100110000;
   28494: result <= 12'b001100101111;
   28495: result <= 12'b001100101111;
   28496: result <= 12'b001100101111;
   28497: result <= 12'b001100101111;
   28498: result <= 12'b001100101111;
   28499: result <= 12'b001100101111;
   28500: result <= 12'b001100101110;
   28501: result <= 12'b001100101110;
   28502: result <= 12'b001100101110;
   28503: result <= 12'b001100101110;
   28504: result <= 12'b001100101110;
   28505: result <= 12'b001100101101;
   28506: result <= 12'b001100101101;
   28507: result <= 12'b001100101101;
   28508: result <= 12'b001100101101;
   28509: result <= 12'b001100101101;
   28510: result <= 12'b001100101101;
   28511: result <= 12'b001100101100;
   28512: result <= 12'b001100101100;
   28513: result <= 12'b001100101100;
   28514: result <= 12'b001100101100;
   28515: result <= 12'b001100101100;
   28516: result <= 12'b001100101011;
   28517: result <= 12'b001100101011;
   28518: result <= 12'b001100101011;
   28519: result <= 12'b001100101011;
   28520: result <= 12'b001100101011;
   28521: result <= 12'b001100101011;
   28522: result <= 12'b001100101010;
   28523: result <= 12'b001100101010;
   28524: result <= 12'b001100101010;
   28525: result <= 12'b001100101010;
   28526: result <= 12'b001100101010;
   28527: result <= 12'b001100101001;
   28528: result <= 12'b001100101001;
   28529: result <= 12'b001100101001;
   28530: result <= 12'b001100101001;
   28531: result <= 12'b001100101001;
   28532: result <= 12'b001100101001;
   28533: result <= 12'b001100101000;
   28534: result <= 12'b001100101000;
   28535: result <= 12'b001100101000;
   28536: result <= 12'b001100101000;
   28537: result <= 12'b001100101000;
   28538: result <= 12'b001100100111;
   28539: result <= 12'b001100100111;
   28540: result <= 12'b001100100111;
   28541: result <= 12'b001100100111;
   28542: result <= 12'b001100100111;
   28543: result <= 12'b001100100111;
   28544: result <= 12'b001100100110;
   28545: result <= 12'b001100100110;
   28546: result <= 12'b001100100110;
   28547: result <= 12'b001100100110;
   28548: result <= 12'b001100100110;
   28549: result <= 12'b001100100101;
   28550: result <= 12'b001100100101;
   28551: result <= 12'b001100100101;
   28552: result <= 12'b001100100101;
   28553: result <= 12'b001100100101;
   28554: result <= 12'b001100100101;
   28555: result <= 12'b001100100100;
   28556: result <= 12'b001100100100;
   28557: result <= 12'b001100100100;
   28558: result <= 12'b001100100100;
   28559: result <= 12'b001100100100;
   28560: result <= 12'b001100100100;
   28561: result <= 12'b001100100011;
   28562: result <= 12'b001100100011;
   28563: result <= 12'b001100100011;
   28564: result <= 12'b001100100011;
   28565: result <= 12'b001100100011;
   28566: result <= 12'b001100100010;
   28567: result <= 12'b001100100010;
   28568: result <= 12'b001100100010;
   28569: result <= 12'b001100100010;
   28570: result <= 12'b001100100010;
   28571: result <= 12'b001100100010;
   28572: result <= 12'b001100100001;
   28573: result <= 12'b001100100001;
   28574: result <= 12'b001100100001;
   28575: result <= 12'b001100100001;
   28576: result <= 12'b001100100001;
   28577: result <= 12'b001100100000;
   28578: result <= 12'b001100100000;
   28579: result <= 12'b001100100000;
   28580: result <= 12'b001100100000;
   28581: result <= 12'b001100100000;
   28582: result <= 12'b001100100000;
   28583: result <= 12'b001100011111;
   28584: result <= 12'b001100011111;
   28585: result <= 12'b001100011111;
   28586: result <= 12'b001100011111;
   28587: result <= 12'b001100011111;
   28588: result <= 12'b001100011110;
   28589: result <= 12'b001100011110;
   28590: result <= 12'b001100011110;
   28591: result <= 12'b001100011110;
   28592: result <= 12'b001100011110;
   28593: result <= 12'b001100011110;
   28594: result <= 12'b001100011101;
   28595: result <= 12'b001100011101;
   28596: result <= 12'b001100011101;
   28597: result <= 12'b001100011101;
   28598: result <= 12'b001100011101;
   28599: result <= 12'b001100011100;
   28600: result <= 12'b001100011100;
   28601: result <= 12'b001100011100;
   28602: result <= 12'b001100011100;
   28603: result <= 12'b001100011100;
   28604: result <= 12'b001100011100;
   28605: result <= 12'b001100011011;
   28606: result <= 12'b001100011011;
   28607: result <= 12'b001100011011;
   28608: result <= 12'b001100011011;
   28609: result <= 12'b001100011011;
   28610: result <= 12'b001100011010;
   28611: result <= 12'b001100011010;
   28612: result <= 12'b001100011010;
   28613: result <= 12'b001100011010;
   28614: result <= 12'b001100011010;
   28615: result <= 12'b001100011010;
   28616: result <= 12'b001100011001;
   28617: result <= 12'b001100011001;
   28618: result <= 12'b001100011001;
   28619: result <= 12'b001100011001;
   28620: result <= 12'b001100011001;
   28621: result <= 12'b001100011000;
   28622: result <= 12'b001100011000;
   28623: result <= 12'b001100011000;
   28624: result <= 12'b001100011000;
   28625: result <= 12'b001100011000;
   28626: result <= 12'b001100011000;
   28627: result <= 12'b001100010111;
   28628: result <= 12'b001100010111;
   28629: result <= 12'b001100010111;
   28630: result <= 12'b001100010111;
   28631: result <= 12'b001100010111;
   28632: result <= 12'b001100010110;
   28633: result <= 12'b001100010110;
   28634: result <= 12'b001100010110;
   28635: result <= 12'b001100010110;
   28636: result <= 12'b001100010110;
   28637: result <= 12'b001100010110;
   28638: result <= 12'b001100010101;
   28639: result <= 12'b001100010101;
   28640: result <= 12'b001100010101;
   28641: result <= 12'b001100010101;
   28642: result <= 12'b001100010101;
   28643: result <= 12'b001100010100;
   28644: result <= 12'b001100010100;
   28645: result <= 12'b001100010100;
   28646: result <= 12'b001100010100;
   28647: result <= 12'b001100010100;
   28648: result <= 12'b001100010100;
   28649: result <= 12'b001100010011;
   28650: result <= 12'b001100010011;
   28651: result <= 12'b001100010011;
   28652: result <= 12'b001100010011;
   28653: result <= 12'b001100010011;
   28654: result <= 12'b001100010010;
   28655: result <= 12'b001100010010;
   28656: result <= 12'b001100010010;
   28657: result <= 12'b001100010010;
   28658: result <= 12'b001100010010;
   28659: result <= 12'b001100010010;
   28660: result <= 12'b001100010001;
   28661: result <= 12'b001100010001;
   28662: result <= 12'b001100010001;
   28663: result <= 12'b001100010001;
   28664: result <= 12'b001100010001;
   28665: result <= 12'b001100010001;
   28666: result <= 12'b001100010000;
   28667: result <= 12'b001100010000;
   28668: result <= 12'b001100010000;
   28669: result <= 12'b001100010000;
   28670: result <= 12'b001100010000;
   28671: result <= 12'b001100001111;
   28672: result <= 12'b001100001111;
   28673: result <= 12'b001100001111;
   28674: result <= 12'b001100001111;
   28675: result <= 12'b001100001111;
   28676: result <= 12'b001100001111;
   28677: result <= 12'b001100001110;
   28678: result <= 12'b001100001110;
   28679: result <= 12'b001100001110;
   28680: result <= 12'b001100001110;
   28681: result <= 12'b001100001110;
   28682: result <= 12'b001100001101;
   28683: result <= 12'b001100001101;
   28684: result <= 12'b001100001101;
   28685: result <= 12'b001100001101;
   28686: result <= 12'b001100001101;
   28687: result <= 12'b001100001101;
   28688: result <= 12'b001100001100;
   28689: result <= 12'b001100001100;
   28690: result <= 12'b001100001100;
   28691: result <= 12'b001100001100;
   28692: result <= 12'b001100001100;
   28693: result <= 12'b001100001011;
   28694: result <= 12'b001100001011;
   28695: result <= 12'b001100001011;
   28696: result <= 12'b001100001011;
   28697: result <= 12'b001100001011;
   28698: result <= 12'b001100001011;
   28699: result <= 12'b001100001010;
   28700: result <= 12'b001100001010;
   28701: result <= 12'b001100001010;
   28702: result <= 12'b001100001010;
   28703: result <= 12'b001100001010;
   28704: result <= 12'b001100001001;
   28705: result <= 12'b001100001001;
   28706: result <= 12'b001100001001;
   28707: result <= 12'b001100001001;
   28708: result <= 12'b001100001001;
   28709: result <= 12'b001100001001;
   28710: result <= 12'b001100001000;
   28711: result <= 12'b001100001000;
   28712: result <= 12'b001100001000;
   28713: result <= 12'b001100001000;
   28714: result <= 12'b001100001000;
   28715: result <= 12'b001100000111;
   28716: result <= 12'b001100000111;
   28717: result <= 12'b001100000111;
   28718: result <= 12'b001100000111;
   28719: result <= 12'b001100000111;
   28720: result <= 12'b001100000111;
   28721: result <= 12'b001100000110;
   28722: result <= 12'b001100000110;
   28723: result <= 12'b001100000110;
   28724: result <= 12'b001100000110;
   28725: result <= 12'b001100000110;
   28726: result <= 12'b001100000101;
   28727: result <= 12'b001100000101;
   28728: result <= 12'b001100000101;
   28729: result <= 12'b001100000101;
   28730: result <= 12'b001100000101;
   28731: result <= 12'b001100000101;
   28732: result <= 12'b001100000100;
   28733: result <= 12'b001100000100;
   28734: result <= 12'b001100000100;
   28735: result <= 12'b001100000100;
   28736: result <= 12'b001100000100;
   28737: result <= 12'b001100000011;
   28738: result <= 12'b001100000011;
   28739: result <= 12'b001100000011;
   28740: result <= 12'b001100000011;
   28741: result <= 12'b001100000011;
   28742: result <= 12'b001100000011;
   28743: result <= 12'b001100000010;
   28744: result <= 12'b001100000010;
   28745: result <= 12'b001100000010;
   28746: result <= 12'b001100000010;
   28747: result <= 12'b001100000010;
   28748: result <= 12'b001100000001;
   28749: result <= 12'b001100000001;
   28750: result <= 12'b001100000001;
   28751: result <= 12'b001100000001;
   28752: result <= 12'b001100000001;
   28753: result <= 12'b001100000001;
   28754: result <= 12'b001100000000;
   28755: result <= 12'b001100000000;
   28756: result <= 12'b001100000000;
   28757: result <= 12'b001100000000;
   28758: result <= 12'b001100000000;
   28759: result <= 12'b001011111111;
   28760: result <= 12'b001011111111;
   28761: result <= 12'b001011111111;
   28762: result <= 12'b001011111111;
   28763: result <= 12'b001011111111;
   28764: result <= 12'b001011111111;
   28765: result <= 12'b001011111110;
   28766: result <= 12'b001011111110;
   28767: result <= 12'b001011111110;
   28768: result <= 12'b001011111110;
   28769: result <= 12'b001011111110;
   28770: result <= 12'b001011111101;
   28771: result <= 12'b001011111101;
   28772: result <= 12'b001011111101;
   28773: result <= 12'b001011111101;
   28774: result <= 12'b001011111101;
   28775: result <= 12'b001011111101;
   28776: result <= 12'b001011111100;
   28777: result <= 12'b001011111100;
   28778: result <= 12'b001011111100;
   28779: result <= 12'b001011111100;
   28780: result <= 12'b001011111100;
   28781: result <= 12'b001011111011;
   28782: result <= 12'b001011111011;
   28783: result <= 12'b001011111011;
   28784: result <= 12'b001011111011;
   28785: result <= 12'b001011111011;
   28786: result <= 12'b001011111011;
   28787: result <= 12'b001011111010;
   28788: result <= 12'b001011111010;
   28789: result <= 12'b001011111010;
   28790: result <= 12'b001011111010;
   28791: result <= 12'b001011111010;
   28792: result <= 12'b001011111001;
   28793: result <= 12'b001011111001;
   28794: result <= 12'b001011111001;
   28795: result <= 12'b001011111001;
   28796: result <= 12'b001011111001;
   28797: result <= 12'b001011111001;
   28798: result <= 12'b001011111000;
   28799: result <= 12'b001011111000;
   28800: result <= 12'b001011111000;
   28801: result <= 12'b001011111000;
   28802: result <= 12'b001011111000;
   28803: result <= 12'b001011110111;
   28804: result <= 12'b001011110111;
   28805: result <= 12'b001011110111;
   28806: result <= 12'b001011110111;
   28807: result <= 12'b001011110111;
   28808: result <= 12'b001011110110;
   28809: result <= 12'b001011110110;
   28810: result <= 12'b001011110110;
   28811: result <= 12'b001011110110;
   28812: result <= 12'b001011110110;
   28813: result <= 12'b001011110110;
   28814: result <= 12'b001011110101;
   28815: result <= 12'b001011110101;
   28816: result <= 12'b001011110101;
   28817: result <= 12'b001011110101;
   28818: result <= 12'b001011110101;
   28819: result <= 12'b001011110100;
   28820: result <= 12'b001011110100;
   28821: result <= 12'b001011110100;
   28822: result <= 12'b001011110100;
   28823: result <= 12'b001011110100;
   28824: result <= 12'b001011110100;
   28825: result <= 12'b001011110011;
   28826: result <= 12'b001011110011;
   28827: result <= 12'b001011110011;
   28828: result <= 12'b001011110011;
   28829: result <= 12'b001011110011;
   28830: result <= 12'b001011110010;
   28831: result <= 12'b001011110010;
   28832: result <= 12'b001011110010;
   28833: result <= 12'b001011110010;
   28834: result <= 12'b001011110010;
   28835: result <= 12'b001011110010;
   28836: result <= 12'b001011110001;
   28837: result <= 12'b001011110001;
   28838: result <= 12'b001011110001;
   28839: result <= 12'b001011110001;
   28840: result <= 12'b001011110001;
   28841: result <= 12'b001011110000;
   28842: result <= 12'b001011110000;
   28843: result <= 12'b001011110000;
   28844: result <= 12'b001011110000;
   28845: result <= 12'b001011110000;
   28846: result <= 12'b001011110000;
   28847: result <= 12'b001011101111;
   28848: result <= 12'b001011101111;
   28849: result <= 12'b001011101111;
   28850: result <= 12'b001011101111;
   28851: result <= 12'b001011101111;
   28852: result <= 12'b001011101110;
   28853: result <= 12'b001011101110;
   28854: result <= 12'b001011101110;
   28855: result <= 12'b001011101110;
   28856: result <= 12'b001011101110;
   28857: result <= 12'b001011101110;
   28858: result <= 12'b001011101101;
   28859: result <= 12'b001011101101;
   28860: result <= 12'b001011101101;
   28861: result <= 12'b001011101101;
   28862: result <= 12'b001011101101;
   28863: result <= 12'b001011101100;
   28864: result <= 12'b001011101100;
   28865: result <= 12'b001011101100;
   28866: result <= 12'b001011101100;
   28867: result <= 12'b001011101100;
   28868: result <= 12'b001011101100;
   28869: result <= 12'b001011101011;
   28870: result <= 12'b001011101011;
   28871: result <= 12'b001011101011;
   28872: result <= 12'b001011101011;
   28873: result <= 12'b001011101011;
   28874: result <= 12'b001011101010;
   28875: result <= 12'b001011101010;
   28876: result <= 12'b001011101010;
   28877: result <= 12'b001011101010;
   28878: result <= 12'b001011101010;
   28879: result <= 12'b001011101010;
   28880: result <= 12'b001011101001;
   28881: result <= 12'b001011101001;
   28882: result <= 12'b001011101001;
   28883: result <= 12'b001011101001;
   28884: result <= 12'b001011101001;
   28885: result <= 12'b001011101000;
   28886: result <= 12'b001011101000;
   28887: result <= 12'b001011101000;
   28888: result <= 12'b001011101000;
   28889: result <= 12'b001011101000;
   28890: result <= 12'b001011101000;
   28891: result <= 12'b001011100111;
   28892: result <= 12'b001011100111;
   28893: result <= 12'b001011100111;
   28894: result <= 12'b001011100111;
   28895: result <= 12'b001011100111;
   28896: result <= 12'b001011100110;
   28897: result <= 12'b001011100110;
   28898: result <= 12'b001011100110;
   28899: result <= 12'b001011100110;
   28900: result <= 12'b001011100110;
   28901: result <= 12'b001011100110;
   28902: result <= 12'b001011100101;
   28903: result <= 12'b001011100101;
   28904: result <= 12'b001011100101;
   28905: result <= 12'b001011100101;
   28906: result <= 12'b001011100101;
   28907: result <= 12'b001011100100;
   28908: result <= 12'b001011100100;
   28909: result <= 12'b001011100100;
   28910: result <= 12'b001011100100;
   28911: result <= 12'b001011100100;
   28912: result <= 12'b001011100011;
   28913: result <= 12'b001011100011;
   28914: result <= 12'b001011100011;
   28915: result <= 12'b001011100011;
   28916: result <= 12'b001011100011;
   28917: result <= 12'b001011100011;
   28918: result <= 12'b001011100010;
   28919: result <= 12'b001011100010;
   28920: result <= 12'b001011100010;
   28921: result <= 12'b001011100010;
   28922: result <= 12'b001011100010;
   28923: result <= 12'b001011100001;
   28924: result <= 12'b001011100001;
   28925: result <= 12'b001011100001;
   28926: result <= 12'b001011100001;
   28927: result <= 12'b001011100001;
   28928: result <= 12'b001011100001;
   28929: result <= 12'b001011100000;
   28930: result <= 12'b001011100000;
   28931: result <= 12'b001011100000;
   28932: result <= 12'b001011100000;
   28933: result <= 12'b001011100000;
   28934: result <= 12'b001011011111;
   28935: result <= 12'b001011011111;
   28936: result <= 12'b001011011111;
   28937: result <= 12'b001011011111;
   28938: result <= 12'b001011011111;
   28939: result <= 12'b001011011111;
   28940: result <= 12'b001011011110;
   28941: result <= 12'b001011011110;
   28942: result <= 12'b001011011110;
   28943: result <= 12'b001011011110;
   28944: result <= 12'b001011011110;
   28945: result <= 12'b001011011101;
   28946: result <= 12'b001011011101;
   28947: result <= 12'b001011011101;
   28948: result <= 12'b001011011101;
   28949: result <= 12'b001011011101;
   28950: result <= 12'b001011011101;
   28951: result <= 12'b001011011100;
   28952: result <= 12'b001011011100;
   28953: result <= 12'b001011011100;
   28954: result <= 12'b001011011100;
   28955: result <= 12'b001011011100;
   28956: result <= 12'b001011011011;
   28957: result <= 12'b001011011011;
   28958: result <= 12'b001011011011;
   28959: result <= 12'b001011011011;
   28960: result <= 12'b001011011011;
   28961: result <= 12'b001011011011;
   28962: result <= 12'b001011011010;
   28963: result <= 12'b001011011010;
   28964: result <= 12'b001011011010;
   28965: result <= 12'b001011011010;
   28966: result <= 12'b001011011010;
   28967: result <= 12'b001011011001;
   28968: result <= 12'b001011011001;
   28969: result <= 12'b001011011001;
   28970: result <= 12'b001011011001;
   28971: result <= 12'b001011011001;
   28972: result <= 12'b001011011000;
   28973: result <= 12'b001011011000;
   28974: result <= 12'b001011011000;
   28975: result <= 12'b001011011000;
   28976: result <= 12'b001011011000;
   28977: result <= 12'b001011011000;
   28978: result <= 12'b001011010111;
   28979: result <= 12'b001011010111;
   28980: result <= 12'b001011010111;
   28981: result <= 12'b001011010111;
   28982: result <= 12'b001011010111;
   28983: result <= 12'b001011010110;
   28984: result <= 12'b001011010110;
   28985: result <= 12'b001011010110;
   28986: result <= 12'b001011010110;
   28987: result <= 12'b001011010110;
   28988: result <= 12'b001011010110;
   28989: result <= 12'b001011010101;
   28990: result <= 12'b001011010101;
   28991: result <= 12'b001011010101;
   28992: result <= 12'b001011010101;
   28993: result <= 12'b001011010101;
   28994: result <= 12'b001011010100;
   28995: result <= 12'b001011010100;
   28996: result <= 12'b001011010100;
   28997: result <= 12'b001011010100;
   28998: result <= 12'b001011010100;
   28999: result <= 12'b001011010100;
   29000: result <= 12'b001011010011;
   29001: result <= 12'b001011010011;
   29002: result <= 12'b001011010011;
   29003: result <= 12'b001011010011;
   29004: result <= 12'b001011010011;
   29005: result <= 12'b001011010010;
   29006: result <= 12'b001011010010;
   29007: result <= 12'b001011010010;
   29008: result <= 12'b001011010010;
   29009: result <= 12'b001011010010;
   29010: result <= 12'b001011010010;
   29011: result <= 12'b001011010001;
   29012: result <= 12'b001011010001;
   29013: result <= 12'b001011010001;
   29014: result <= 12'b001011010001;
   29015: result <= 12'b001011010001;
   29016: result <= 12'b001011010000;
   29017: result <= 12'b001011010000;
   29018: result <= 12'b001011010000;
   29019: result <= 12'b001011010000;
   29020: result <= 12'b001011010000;
   29021: result <= 12'b001011001111;
   29022: result <= 12'b001011001111;
   29023: result <= 12'b001011001111;
   29024: result <= 12'b001011001111;
   29025: result <= 12'b001011001111;
   29026: result <= 12'b001011001111;
   29027: result <= 12'b001011001110;
   29028: result <= 12'b001011001110;
   29029: result <= 12'b001011001110;
   29030: result <= 12'b001011001110;
   29031: result <= 12'b001011001110;
   29032: result <= 12'b001011001101;
   29033: result <= 12'b001011001101;
   29034: result <= 12'b001011001101;
   29035: result <= 12'b001011001101;
   29036: result <= 12'b001011001101;
   29037: result <= 12'b001011001101;
   29038: result <= 12'b001011001100;
   29039: result <= 12'b001011001100;
   29040: result <= 12'b001011001100;
   29041: result <= 12'b001011001100;
   29042: result <= 12'b001011001100;
   29043: result <= 12'b001011001011;
   29044: result <= 12'b001011001011;
   29045: result <= 12'b001011001011;
   29046: result <= 12'b001011001011;
   29047: result <= 12'b001011001011;
   29048: result <= 12'b001011001011;
   29049: result <= 12'b001011001010;
   29050: result <= 12'b001011001010;
   29051: result <= 12'b001011001010;
   29052: result <= 12'b001011001010;
   29053: result <= 12'b001011001010;
   29054: result <= 12'b001011001001;
   29055: result <= 12'b001011001001;
   29056: result <= 12'b001011001001;
   29057: result <= 12'b001011001001;
   29058: result <= 12'b001011001001;
   29059: result <= 12'b001011001001;
   29060: result <= 12'b001011001000;
   29061: result <= 12'b001011001000;
   29062: result <= 12'b001011001000;
   29063: result <= 12'b001011001000;
   29064: result <= 12'b001011001000;
   29065: result <= 12'b001011000111;
   29066: result <= 12'b001011000111;
   29067: result <= 12'b001011000111;
   29068: result <= 12'b001011000111;
   29069: result <= 12'b001011000111;
   29070: result <= 12'b001011000110;
   29071: result <= 12'b001011000110;
   29072: result <= 12'b001011000110;
   29073: result <= 12'b001011000110;
   29074: result <= 12'b001011000110;
   29075: result <= 12'b001011000110;
   29076: result <= 12'b001011000101;
   29077: result <= 12'b001011000101;
   29078: result <= 12'b001011000101;
   29079: result <= 12'b001011000101;
   29080: result <= 12'b001011000101;
   29081: result <= 12'b001011000100;
   29082: result <= 12'b001011000100;
   29083: result <= 12'b001011000100;
   29084: result <= 12'b001011000100;
   29085: result <= 12'b001011000100;
   29086: result <= 12'b001011000100;
   29087: result <= 12'b001011000011;
   29088: result <= 12'b001011000011;
   29089: result <= 12'b001011000011;
   29090: result <= 12'b001011000011;
   29091: result <= 12'b001011000011;
   29092: result <= 12'b001011000010;
   29093: result <= 12'b001011000010;
   29094: result <= 12'b001011000010;
   29095: result <= 12'b001011000010;
   29096: result <= 12'b001011000010;
   29097: result <= 12'b001011000010;
   29098: result <= 12'b001011000001;
   29099: result <= 12'b001011000001;
   29100: result <= 12'b001011000001;
   29101: result <= 12'b001011000001;
   29102: result <= 12'b001011000001;
   29103: result <= 12'b001011000000;
   29104: result <= 12'b001011000000;
   29105: result <= 12'b001011000000;
   29106: result <= 12'b001011000000;
   29107: result <= 12'b001011000000;
   29108: result <= 12'b001010111111;
   29109: result <= 12'b001010111111;
   29110: result <= 12'b001010111111;
   29111: result <= 12'b001010111111;
   29112: result <= 12'b001010111111;
   29113: result <= 12'b001010111111;
   29114: result <= 12'b001010111110;
   29115: result <= 12'b001010111110;
   29116: result <= 12'b001010111110;
   29117: result <= 12'b001010111110;
   29118: result <= 12'b001010111110;
   29119: result <= 12'b001010111101;
   29120: result <= 12'b001010111101;
   29121: result <= 12'b001010111101;
   29122: result <= 12'b001010111101;
   29123: result <= 12'b001010111101;
   29124: result <= 12'b001010111101;
   29125: result <= 12'b001010111100;
   29126: result <= 12'b001010111100;
   29127: result <= 12'b001010111100;
   29128: result <= 12'b001010111100;
   29129: result <= 12'b001010111100;
   29130: result <= 12'b001010111011;
   29131: result <= 12'b001010111011;
   29132: result <= 12'b001010111011;
   29133: result <= 12'b001010111011;
   29134: result <= 12'b001010111011;
   29135: result <= 12'b001010111011;
   29136: result <= 12'b001010111010;
   29137: result <= 12'b001010111010;
   29138: result <= 12'b001010111010;
   29139: result <= 12'b001010111010;
   29140: result <= 12'b001010111010;
   29141: result <= 12'b001010111001;
   29142: result <= 12'b001010111001;
   29143: result <= 12'b001010111001;
   29144: result <= 12'b001010111001;
   29145: result <= 12'b001010111001;
   29146: result <= 12'b001010111000;
   29147: result <= 12'b001010111000;
   29148: result <= 12'b001010111000;
   29149: result <= 12'b001010111000;
   29150: result <= 12'b001010111000;
   29151: result <= 12'b001010111000;
   29152: result <= 12'b001010110111;
   29153: result <= 12'b001010110111;
   29154: result <= 12'b001010110111;
   29155: result <= 12'b001010110111;
   29156: result <= 12'b001010110111;
   29157: result <= 12'b001010110110;
   29158: result <= 12'b001010110110;
   29159: result <= 12'b001010110110;
   29160: result <= 12'b001010110110;
   29161: result <= 12'b001010110110;
   29162: result <= 12'b001010110110;
   29163: result <= 12'b001010110101;
   29164: result <= 12'b001010110101;
   29165: result <= 12'b001010110101;
   29166: result <= 12'b001010110101;
   29167: result <= 12'b001010110101;
   29168: result <= 12'b001010110100;
   29169: result <= 12'b001010110100;
   29170: result <= 12'b001010110100;
   29171: result <= 12'b001010110100;
   29172: result <= 12'b001010110100;
   29173: result <= 12'b001010110011;
   29174: result <= 12'b001010110011;
   29175: result <= 12'b001010110011;
   29176: result <= 12'b001010110011;
   29177: result <= 12'b001010110011;
   29178: result <= 12'b001010110011;
   29179: result <= 12'b001010110010;
   29180: result <= 12'b001010110010;
   29181: result <= 12'b001010110010;
   29182: result <= 12'b001010110010;
   29183: result <= 12'b001010110010;
   29184: result <= 12'b001010110001;
   29185: result <= 12'b001010110001;
   29186: result <= 12'b001010110001;
   29187: result <= 12'b001010110001;
   29188: result <= 12'b001010110001;
   29189: result <= 12'b001010110001;
   29190: result <= 12'b001010110000;
   29191: result <= 12'b001010110000;
   29192: result <= 12'b001010110000;
   29193: result <= 12'b001010110000;
   29194: result <= 12'b001010110000;
   29195: result <= 12'b001010101111;
   29196: result <= 12'b001010101111;
   29197: result <= 12'b001010101111;
   29198: result <= 12'b001010101111;
   29199: result <= 12'b001010101111;
   29200: result <= 12'b001010101110;
   29201: result <= 12'b001010101110;
   29202: result <= 12'b001010101110;
   29203: result <= 12'b001010101110;
   29204: result <= 12'b001010101110;
   29205: result <= 12'b001010101110;
   29206: result <= 12'b001010101101;
   29207: result <= 12'b001010101101;
   29208: result <= 12'b001010101101;
   29209: result <= 12'b001010101101;
   29210: result <= 12'b001010101101;
   29211: result <= 12'b001010101100;
   29212: result <= 12'b001010101100;
   29213: result <= 12'b001010101100;
   29214: result <= 12'b001010101100;
   29215: result <= 12'b001010101100;
   29216: result <= 12'b001010101100;
   29217: result <= 12'b001010101011;
   29218: result <= 12'b001010101011;
   29219: result <= 12'b001010101011;
   29220: result <= 12'b001010101011;
   29221: result <= 12'b001010101011;
   29222: result <= 12'b001010101010;
   29223: result <= 12'b001010101010;
   29224: result <= 12'b001010101010;
   29225: result <= 12'b001010101010;
   29226: result <= 12'b001010101010;
   29227: result <= 12'b001010101001;
   29228: result <= 12'b001010101001;
   29229: result <= 12'b001010101001;
   29230: result <= 12'b001010101001;
   29231: result <= 12'b001010101001;
   29232: result <= 12'b001010101001;
   29233: result <= 12'b001010101000;
   29234: result <= 12'b001010101000;
   29235: result <= 12'b001010101000;
   29236: result <= 12'b001010101000;
   29237: result <= 12'b001010101000;
   29238: result <= 12'b001010100111;
   29239: result <= 12'b001010100111;
   29240: result <= 12'b001010100111;
   29241: result <= 12'b001010100111;
   29242: result <= 12'b001010100111;
   29243: result <= 12'b001010100111;
   29244: result <= 12'b001010100110;
   29245: result <= 12'b001010100110;
   29246: result <= 12'b001010100110;
   29247: result <= 12'b001010100110;
   29248: result <= 12'b001010100110;
   29249: result <= 12'b001010100101;
   29250: result <= 12'b001010100101;
   29251: result <= 12'b001010100101;
   29252: result <= 12'b001010100101;
   29253: result <= 12'b001010100101;
   29254: result <= 12'b001010100100;
   29255: result <= 12'b001010100100;
   29256: result <= 12'b001010100100;
   29257: result <= 12'b001010100100;
   29258: result <= 12'b001010100100;
   29259: result <= 12'b001010100100;
   29260: result <= 12'b001010100011;
   29261: result <= 12'b001010100011;
   29262: result <= 12'b001010100011;
   29263: result <= 12'b001010100011;
   29264: result <= 12'b001010100011;
   29265: result <= 12'b001010100010;
   29266: result <= 12'b001010100010;
   29267: result <= 12'b001010100010;
   29268: result <= 12'b001010100010;
   29269: result <= 12'b001010100010;
   29270: result <= 12'b001010100010;
   29271: result <= 12'b001010100001;
   29272: result <= 12'b001010100001;
   29273: result <= 12'b001010100001;
   29274: result <= 12'b001010100001;
   29275: result <= 12'b001010100001;
   29276: result <= 12'b001010100000;
   29277: result <= 12'b001010100000;
   29278: result <= 12'b001010100000;
   29279: result <= 12'b001010100000;
   29280: result <= 12'b001010100000;
   29281: result <= 12'b001010011111;
   29282: result <= 12'b001010011111;
   29283: result <= 12'b001010011111;
   29284: result <= 12'b001010011111;
   29285: result <= 12'b001010011111;
   29286: result <= 12'b001010011111;
   29287: result <= 12'b001010011110;
   29288: result <= 12'b001010011110;
   29289: result <= 12'b001010011110;
   29290: result <= 12'b001010011110;
   29291: result <= 12'b001010011110;
   29292: result <= 12'b001010011101;
   29293: result <= 12'b001010011101;
   29294: result <= 12'b001010011101;
   29295: result <= 12'b001010011101;
   29296: result <= 12'b001010011101;
   29297: result <= 12'b001010011101;
   29298: result <= 12'b001010011100;
   29299: result <= 12'b001010011100;
   29300: result <= 12'b001010011100;
   29301: result <= 12'b001010011100;
   29302: result <= 12'b001010011100;
   29303: result <= 12'b001010011011;
   29304: result <= 12'b001010011011;
   29305: result <= 12'b001010011011;
   29306: result <= 12'b001010011011;
   29307: result <= 12'b001010011011;
   29308: result <= 12'b001010011010;
   29309: result <= 12'b001010011010;
   29310: result <= 12'b001010011010;
   29311: result <= 12'b001010011010;
   29312: result <= 12'b001010011010;
   29313: result <= 12'b001010011010;
   29314: result <= 12'b001010011001;
   29315: result <= 12'b001010011001;
   29316: result <= 12'b001010011001;
   29317: result <= 12'b001010011001;
   29318: result <= 12'b001010011001;
   29319: result <= 12'b001010011000;
   29320: result <= 12'b001010011000;
   29321: result <= 12'b001010011000;
   29322: result <= 12'b001010011000;
   29323: result <= 12'b001010011000;
   29324: result <= 12'b001010011000;
   29325: result <= 12'b001010010111;
   29326: result <= 12'b001010010111;
   29327: result <= 12'b001010010111;
   29328: result <= 12'b001010010111;
   29329: result <= 12'b001010010111;
   29330: result <= 12'b001010010110;
   29331: result <= 12'b001010010110;
   29332: result <= 12'b001010010110;
   29333: result <= 12'b001010010110;
   29334: result <= 12'b001010010110;
   29335: result <= 12'b001010010101;
   29336: result <= 12'b001010010101;
   29337: result <= 12'b001010010101;
   29338: result <= 12'b001010010101;
   29339: result <= 12'b001010010101;
   29340: result <= 12'b001010010101;
   29341: result <= 12'b001010010100;
   29342: result <= 12'b001010010100;
   29343: result <= 12'b001010010100;
   29344: result <= 12'b001010010100;
   29345: result <= 12'b001010010100;
   29346: result <= 12'b001010010011;
   29347: result <= 12'b001010010011;
   29348: result <= 12'b001010010011;
   29349: result <= 12'b001010010011;
   29350: result <= 12'b001010010011;
   29351: result <= 12'b001010010010;
   29352: result <= 12'b001010010010;
   29353: result <= 12'b001010010010;
   29354: result <= 12'b001010010010;
   29355: result <= 12'b001010010010;
   29356: result <= 12'b001010010010;
   29357: result <= 12'b001010010001;
   29358: result <= 12'b001010010001;
   29359: result <= 12'b001010010001;
   29360: result <= 12'b001010010001;
   29361: result <= 12'b001010010001;
   29362: result <= 12'b001010010000;
   29363: result <= 12'b001010010000;
   29364: result <= 12'b001010010000;
   29365: result <= 12'b001010010000;
   29366: result <= 12'b001010010000;
   29367: result <= 12'b001010010000;
   29368: result <= 12'b001010001111;
   29369: result <= 12'b001010001111;
   29370: result <= 12'b001010001111;
   29371: result <= 12'b001010001111;
   29372: result <= 12'b001010001111;
   29373: result <= 12'b001010001110;
   29374: result <= 12'b001010001110;
   29375: result <= 12'b001010001110;
   29376: result <= 12'b001010001110;
   29377: result <= 12'b001010001110;
   29378: result <= 12'b001010001101;
   29379: result <= 12'b001010001101;
   29380: result <= 12'b001010001101;
   29381: result <= 12'b001010001101;
   29382: result <= 12'b001010001101;
   29383: result <= 12'b001010001101;
   29384: result <= 12'b001010001100;
   29385: result <= 12'b001010001100;
   29386: result <= 12'b001010001100;
   29387: result <= 12'b001010001100;
   29388: result <= 12'b001010001100;
   29389: result <= 12'b001010001011;
   29390: result <= 12'b001010001011;
   29391: result <= 12'b001010001011;
   29392: result <= 12'b001010001011;
   29393: result <= 12'b001010001011;
   29394: result <= 12'b001010001010;
   29395: result <= 12'b001010001010;
   29396: result <= 12'b001010001010;
   29397: result <= 12'b001010001010;
   29398: result <= 12'b001010001010;
   29399: result <= 12'b001010001010;
   29400: result <= 12'b001010001001;
   29401: result <= 12'b001010001001;
   29402: result <= 12'b001010001001;
   29403: result <= 12'b001010001001;
   29404: result <= 12'b001010001001;
   29405: result <= 12'b001010001000;
   29406: result <= 12'b001010001000;
   29407: result <= 12'b001010001000;
   29408: result <= 12'b001010001000;
   29409: result <= 12'b001010001000;
   29410: result <= 12'b001010001000;
   29411: result <= 12'b001010000111;
   29412: result <= 12'b001010000111;
   29413: result <= 12'b001010000111;
   29414: result <= 12'b001010000111;
   29415: result <= 12'b001010000111;
   29416: result <= 12'b001010000110;
   29417: result <= 12'b001010000110;
   29418: result <= 12'b001010000110;
   29419: result <= 12'b001010000110;
   29420: result <= 12'b001010000110;
   29421: result <= 12'b001010000101;
   29422: result <= 12'b001010000101;
   29423: result <= 12'b001010000101;
   29424: result <= 12'b001010000101;
   29425: result <= 12'b001010000101;
   29426: result <= 12'b001010000101;
   29427: result <= 12'b001010000100;
   29428: result <= 12'b001010000100;
   29429: result <= 12'b001010000100;
   29430: result <= 12'b001010000100;
   29431: result <= 12'b001010000100;
   29432: result <= 12'b001010000011;
   29433: result <= 12'b001010000011;
   29434: result <= 12'b001010000011;
   29435: result <= 12'b001010000011;
   29436: result <= 12'b001010000011;
   29437: result <= 12'b001010000010;
   29438: result <= 12'b001010000010;
   29439: result <= 12'b001010000010;
   29440: result <= 12'b001010000010;
   29441: result <= 12'b001010000010;
   29442: result <= 12'b001010000010;
   29443: result <= 12'b001010000001;
   29444: result <= 12'b001010000001;
   29445: result <= 12'b001010000001;
   29446: result <= 12'b001010000001;
   29447: result <= 12'b001010000001;
   29448: result <= 12'b001010000000;
   29449: result <= 12'b001010000000;
   29450: result <= 12'b001010000000;
   29451: result <= 12'b001010000000;
   29452: result <= 12'b001010000000;
   29453: result <= 12'b001001111111;
   29454: result <= 12'b001001111111;
   29455: result <= 12'b001001111111;
   29456: result <= 12'b001001111111;
   29457: result <= 12'b001001111111;
   29458: result <= 12'b001001111111;
   29459: result <= 12'b001001111110;
   29460: result <= 12'b001001111110;
   29461: result <= 12'b001001111110;
   29462: result <= 12'b001001111110;
   29463: result <= 12'b001001111110;
   29464: result <= 12'b001001111101;
   29465: result <= 12'b001001111101;
   29466: result <= 12'b001001111101;
   29467: result <= 12'b001001111101;
   29468: result <= 12'b001001111101;
   29469: result <= 12'b001001111101;
   29470: result <= 12'b001001111100;
   29471: result <= 12'b001001111100;
   29472: result <= 12'b001001111100;
   29473: result <= 12'b001001111100;
   29474: result <= 12'b001001111100;
   29475: result <= 12'b001001111011;
   29476: result <= 12'b001001111011;
   29477: result <= 12'b001001111011;
   29478: result <= 12'b001001111011;
   29479: result <= 12'b001001111011;
   29480: result <= 12'b001001111010;
   29481: result <= 12'b001001111010;
   29482: result <= 12'b001001111010;
   29483: result <= 12'b001001111010;
   29484: result <= 12'b001001111010;
   29485: result <= 12'b001001111010;
   29486: result <= 12'b001001111001;
   29487: result <= 12'b001001111001;
   29488: result <= 12'b001001111001;
   29489: result <= 12'b001001111001;
   29490: result <= 12'b001001111001;
   29491: result <= 12'b001001111000;
   29492: result <= 12'b001001111000;
   29493: result <= 12'b001001111000;
   29494: result <= 12'b001001111000;
   29495: result <= 12'b001001111000;
   29496: result <= 12'b001001110111;
   29497: result <= 12'b001001110111;
   29498: result <= 12'b001001110111;
   29499: result <= 12'b001001110111;
   29500: result <= 12'b001001110111;
   29501: result <= 12'b001001110111;
   29502: result <= 12'b001001110110;
   29503: result <= 12'b001001110110;
   29504: result <= 12'b001001110110;
   29505: result <= 12'b001001110110;
   29506: result <= 12'b001001110110;
   29507: result <= 12'b001001110101;
   29508: result <= 12'b001001110101;
   29509: result <= 12'b001001110101;
   29510: result <= 12'b001001110101;
   29511: result <= 12'b001001110101;
   29512: result <= 12'b001001110100;
   29513: result <= 12'b001001110100;
   29514: result <= 12'b001001110100;
   29515: result <= 12'b001001110100;
   29516: result <= 12'b001001110100;
   29517: result <= 12'b001001110100;
   29518: result <= 12'b001001110011;
   29519: result <= 12'b001001110011;
   29520: result <= 12'b001001110011;
   29521: result <= 12'b001001110011;
   29522: result <= 12'b001001110011;
   29523: result <= 12'b001001110010;
   29524: result <= 12'b001001110010;
   29525: result <= 12'b001001110010;
   29526: result <= 12'b001001110010;
   29527: result <= 12'b001001110010;
   29528: result <= 12'b001001110001;
   29529: result <= 12'b001001110001;
   29530: result <= 12'b001001110001;
   29531: result <= 12'b001001110001;
   29532: result <= 12'b001001110001;
   29533: result <= 12'b001001110001;
   29534: result <= 12'b001001110000;
   29535: result <= 12'b001001110000;
   29536: result <= 12'b001001110000;
   29537: result <= 12'b001001110000;
   29538: result <= 12'b001001110000;
   29539: result <= 12'b001001101111;
   29540: result <= 12'b001001101111;
   29541: result <= 12'b001001101111;
   29542: result <= 12'b001001101111;
   29543: result <= 12'b001001101111;
   29544: result <= 12'b001001101110;
   29545: result <= 12'b001001101110;
   29546: result <= 12'b001001101110;
   29547: result <= 12'b001001101110;
   29548: result <= 12'b001001101110;
   29549: result <= 12'b001001101110;
   29550: result <= 12'b001001101101;
   29551: result <= 12'b001001101101;
   29552: result <= 12'b001001101101;
   29553: result <= 12'b001001101101;
   29554: result <= 12'b001001101101;
   29555: result <= 12'b001001101100;
   29556: result <= 12'b001001101100;
   29557: result <= 12'b001001101100;
   29558: result <= 12'b001001101100;
   29559: result <= 12'b001001101100;
   29560: result <= 12'b001001101100;
   29561: result <= 12'b001001101011;
   29562: result <= 12'b001001101011;
   29563: result <= 12'b001001101011;
   29564: result <= 12'b001001101011;
   29565: result <= 12'b001001101011;
   29566: result <= 12'b001001101010;
   29567: result <= 12'b001001101010;
   29568: result <= 12'b001001101010;
   29569: result <= 12'b001001101010;
   29570: result <= 12'b001001101010;
   29571: result <= 12'b001001101001;
   29572: result <= 12'b001001101001;
   29573: result <= 12'b001001101001;
   29574: result <= 12'b001001101001;
   29575: result <= 12'b001001101001;
   29576: result <= 12'b001001101001;
   29577: result <= 12'b001001101000;
   29578: result <= 12'b001001101000;
   29579: result <= 12'b001001101000;
   29580: result <= 12'b001001101000;
   29581: result <= 12'b001001101000;
   29582: result <= 12'b001001100111;
   29583: result <= 12'b001001100111;
   29584: result <= 12'b001001100111;
   29585: result <= 12'b001001100111;
   29586: result <= 12'b001001100111;
   29587: result <= 12'b001001100110;
   29588: result <= 12'b001001100110;
   29589: result <= 12'b001001100110;
   29590: result <= 12'b001001100110;
   29591: result <= 12'b001001100110;
   29592: result <= 12'b001001100110;
   29593: result <= 12'b001001100101;
   29594: result <= 12'b001001100101;
   29595: result <= 12'b001001100101;
   29596: result <= 12'b001001100101;
   29597: result <= 12'b001001100101;
   29598: result <= 12'b001001100100;
   29599: result <= 12'b001001100100;
   29600: result <= 12'b001001100100;
   29601: result <= 12'b001001100100;
   29602: result <= 12'b001001100100;
   29603: result <= 12'b001001100011;
   29604: result <= 12'b001001100011;
   29605: result <= 12'b001001100011;
   29606: result <= 12'b001001100011;
   29607: result <= 12'b001001100011;
   29608: result <= 12'b001001100011;
   29609: result <= 12'b001001100010;
   29610: result <= 12'b001001100010;
   29611: result <= 12'b001001100010;
   29612: result <= 12'b001001100010;
   29613: result <= 12'b001001100010;
   29614: result <= 12'b001001100001;
   29615: result <= 12'b001001100001;
   29616: result <= 12'b001001100001;
   29617: result <= 12'b001001100001;
   29618: result <= 12'b001001100001;
   29619: result <= 12'b001001100000;
   29620: result <= 12'b001001100000;
   29621: result <= 12'b001001100000;
   29622: result <= 12'b001001100000;
   29623: result <= 12'b001001100000;
   29624: result <= 12'b001001100000;
   29625: result <= 12'b001001011111;
   29626: result <= 12'b001001011111;
   29627: result <= 12'b001001011111;
   29628: result <= 12'b001001011111;
   29629: result <= 12'b001001011111;
   29630: result <= 12'b001001011110;
   29631: result <= 12'b001001011110;
   29632: result <= 12'b001001011110;
   29633: result <= 12'b001001011110;
   29634: result <= 12'b001001011110;
   29635: result <= 12'b001001011101;
   29636: result <= 12'b001001011101;
   29637: result <= 12'b001001011101;
   29638: result <= 12'b001001011101;
   29639: result <= 12'b001001011101;
   29640: result <= 12'b001001011101;
   29641: result <= 12'b001001011100;
   29642: result <= 12'b001001011100;
   29643: result <= 12'b001001011100;
   29644: result <= 12'b001001011100;
   29645: result <= 12'b001001011100;
   29646: result <= 12'b001001011011;
   29647: result <= 12'b001001011011;
   29648: result <= 12'b001001011011;
   29649: result <= 12'b001001011011;
   29650: result <= 12'b001001011011;
   29651: result <= 12'b001001011010;
   29652: result <= 12'b001001011010;
   29653: result <= 12'b001001011010;
   29654: result <= 12'b001001011010;
   29655: result <= 12'b001001011010;
   29656: result <= 12'b001001011010;
   29657: result <= 12'b001001011001;
   29658: result <= 12'b001001011001;
   29659: result <= 12'b001001011001;
   29660: result <= 12'b001001011001;
   29661: result <= 12'b001001011001;
   29662: result <= 12'b001001011000;
   29663: result <= 12'b001001011000;
   29664: result <= 12'b001001011000;
   29665: result <= 12'b001001011000;
   29666: result <= 12'b001001011000;
   29667: result <= 12'b001001010111;
   29668: result <= 12'b001001010111;
   29669: result <= 12'b001001010111;
   29670: result <= 12'b001001010111;
   29671: result <= 12'b001001010111;
   29672: result <= 12'b001001010111;
   29673: result <= 12'b001001010110;
   29674: result <= 12'b001001010110;
   29675: result <= 12'b001001010110;
   29676: result <= 12'b001001010110;
   29677: result <= 12'b001001010110;
   29678: result <= 12'b001001010101;
   29679: result <= 12'b001001010101;
   29680: result <= 12'b001001010101;
   29681: result <= 12'b001001010101;
   29682: result <= 12'b001001010101;
   29683: result <= 12'b001001010100;
   29684: result <= 12'b001001010100;
   29685: result <= 12'b001001010100;
   29686: result <= 12'b001001010100;
   29687: result <= 12'b001001010100;
   29688: result <= 12'b001001010100;
   29689: result <= 12'b001001010011;
   29690: result <= 12'b001001010011;
   29691: result <= 12'b001001010011;
   29692: result <= 12'b001001010011;
   29693: result <= 12'b001001010011;
   29694: result <= 12'b001001010010;
   29695: result <= 12'b001001010010;
   29696: result <= 12'b001001010010;
   29697: result <= 12'b001001010010;
   29698: result <= 12'b001001010010;
   29699: result <= 12'b001001010001;
   29700: result <= 12'b001001010001;
   29701: result <= 12'b001001010001;
   29702: result <= 12'b001001010001;
   29703: result <= 12'b001001010001;
   29704: result <= 12'b001001010000;
   29705: result <= 12'b001001010000;
   29706: result <= 12'b001001010000;
   29707: result <= 12'b001001010000;
   29708: result <= 12'b001001010000;
   29709: result <= 12'b001001010000;
   29710: result <= 12'b001001001111;
   29711: result <= 12'b001001001111;
   29712: result <= 12'b001001001111;
   29713: result <= 12'b001001001111;
   29714: result <= 12'b001001001111;
   29715: result <= 12'b001001001110;
   29716: result <= 12'b001001001110;
   29717: result <= 12'b001001001110;
   29718: result <= 12'b001001001110;
   29719: result <= 12'b001001001110;
   29720: result <= 12'b001001001101;
   29721: result <= 12'b001001001101;
   29722: result <= 12'b001001001101;
   29723: result <= 12'b001001001101;
   29724: result <= 12'b001001001101;
   29725: result <= 12'b001001001101;
   29726: result <= 12'b001001001100;
   29727: result <= 12'b001001001100;
   29728: result <= 12'b001001001100;
   29729: result <= 12'b001001001100;
   29730: result <= 12'b001001001100;
   29731: result <= 12'b001001001011;
   29732: result <= 12'b001001001011;
   29733: result <= 12'b001001001011;
   29734: result <= 12'b001001001011;
   29735: result <= 12'b001001001011;
   29736: result <= 12'b001001001010;
   29737: result <= 12'b001001001010;
   29738: result <= 12'b001001001010;
   29739: result <= 12'b001001001010;
   29740: result <= 12'b001001001010;
   29741: result <= 12'b001001001010;
   29742: result <= 12'b001001001001;
   29743: result <= 12'b001001001001;
   29744: result <= 12'b001001001001;
   29745: result <= 12'b001001001001;
   29746: result <= 12'b001001001001;
   29747: result <= 12'b001001001000;
   29748: result <= 12'b001001001000;
   29749: result <= 12'b001001001000;
   29750: result <= 12'b001001001000;
   29751: result <= 12'b001001001000;
   29752: result <= 12'b001001000111;
   29753: result <= 12'b001001000111;
   29754: result <= 12'b001001000111;
   29755: result <= 12'b001001000111;
   29756: result <= 12'b001001000111;
   29757: result <= 12'b001001000111;
   29758: result <= 12'b001001000110;
   29759: result <= 12'b001001000110;
   29760: result <= 12'b001001000110;
   29761: result <= 12'b001001000110;
   29762: result <= 12'b001001000110;
   29763: result <= 12'b001001000101;
   29764: result <= 12'b001001000101;
   29765: result <= 12'b001001000101;
   29766: result <= 12'b001001000101;
   29767: result <= 12'b001001000101;
   29768: result <= 12'b001001000100;
   29769: result <= 12'b001001000100;
   29770: result <= 12'b001001000100;
   29771: result <= 12'b001001000100;
   29772: result <= 12'b001001000100;
   29773: result <= 12'b001001000100;
   29774: result <= 12'b001001000011;
   29775: result <= 12'b001001000011;
   29776: result <= 12'b001001000011;
   29777: result <= 12'b001001000011;
   29778: result <= 12'b001001000011;
   29779: result <= 12'b001001000010;
   29780: result <= 12'b001001000010;
   29781: result <= 12'b001001000010;
   29782: result <= 12'b001001000010;
   29783: result <= 12'b001001000010;
   29784: result <= 12'b001001000001;
   29785: result <= 12'b001001000001;
   29786: result <= 12'b001001000001;
   29787: result <= 12'b001001000001;
   29788: result <= 12'b001001000001;
   29789: result <= 12'b001001000001;
   29790: result <= 12'b001001000000;
   29791: result <= 12'b001001000000;
   29792: result <= 12'b001001000000;
   29793: result <= 12'b001001000000;
   29794: result <= 12'b001001000000;
   29795: result <= 12'b001000111111;
   29796: result <= 12'b001000111111;
   29797: result <= 12'b001000111111;
   29798: result <= 12'b001000111111;
   29799: result <= 12'b001000111111;
   29800: result <= 12'b001000111110;
   29801: result <= 12'b001000111110;
   29802: result <= 12'b001000111110;
   29803: result <= 12'b001000111110;
   29804: result <= 12'b001000111110;
   29805: result <= 12'b001000111101;
   29806: result <= 12'b001000111101;
   29807: result <= 12'b001000111101;
   29808: result <= 12'b001000111101;
   29809: result <= 12'b001000111101;
   29810: result <= 12'b001000111101;
   29811: result <= 12'b001000111100;
   29812: result <= 12'b001000111100;
   29813: result <= 12'b001000111100;
   29814: result <= 12'b001000111100;
   29815: result <= 12'b001000111100;
   29816: result <= 12'b001000111011;
   29817: result <= 12'b001000111011;
   29818: result <= 12'b001000111011;
   29819: result <= 12'b001000111011;
   29820: result <= 12'b001000111011;
   29821: result <= 12'b001000111010;
   29822: result <= 12'b001000111010;
   29823: result <= 12'b001000111010;
   29824: result <= 12'b001000111010;
   29825: result <= 12'b001000111010;
   29826: result <= 12'b001000111010;
   29827: result <= 12'b001000111001;
   29828: result <= 12'b001000111001;
   29829: result <= 12'b001000111001;
   29830: result <= 12'b001000111001;
   29831: result <= 12'b001000111001;
   29832: result <= 12'b001000111000;
   29833: result <= 12'b001000111000;
   29834: result <= 12'b001000111000;
   29835: result <= 12'b001000111000;
   29836: result <= 12'b001000111000;
   29837: result <= 12'b001000110111;
   29838: result <= 12'b001000110111;
   29839: result <= 12'b001000110111;
   29840: result <= 12'b001000110111;
   29841: result <= 12'b001000110111;
   29842: result <= 12'b001000110111;
   29843: result <= 12'b001000110110;
   29844: result <= 12'b001000110110;
   29845: result <= 12'b001000110110;
   29846: result <= 12'b001000110110;
   29847: result <= 12'b001000110110;
   29848: result <= 12'b001000110101;
   29849: result <= 12'b001000110101;
   29850: result <= 12'b001000110101;
   29851: result <= 12'b001000110101;
   29852: result <= 12'b001000110101;
   29853: result <= 12'b001000110100;
   29854: result <= 12'b001000110100;
   29855: result <= 12'b001000110100;
   29856: result <= 12'b001000110100;
   29857: result <= 12'b001000110100;
   29858: result <= 12'b001000110011;
   29859: result <= 12'b001000110011;
   29860: result <= 12'b001000110011;
   29861: result <= 12'b001000110011;
   29862: result <= 12'b001000110011;
   29863: result <= 12'b001000110011;
   29864: result <= 12'b001000110010;
   29865: result <= 12'b001000110010;
   29866: result <= 12'b001000110010;
   29867: result <= 12'b001000110010;
   29868: result <= 12'b001000110010;
   29869: result <= 12'b001000110001;
   29870: result <= 12'b001000110001;
   29871: result <= 12'b001000110001;
   29872: result <= 12'b001000110001;
   29873: result <= 12'b001000110001;
   29874: result <= 12'b001000110000;
   29875: result <= 12'b001000110000;
   29876: result <= 12'b001000110000;
   29877: result <= 12'b001000110000;
   29878: result <= 12'b001000110000;
   29879: result <= 12'b001000110000;
   29880: result <= 12'b001000101111;
   29881: result <= 12'b001000101111;
   29882: result <= 12'b001000101111;
   29883: result <= 12'b001000101111;
   29884: result <= 12'b001000101111;
   29885: result <= 12'b001000101110;
   29886: result <= 12'b001000101110;
   29887: result <= 12'b001000101110;
   29888: result <= 12'b001000101110;
   29889: result <= 12'b001000101110;
   29890: result <= 12'b001000101101;
   29891: result <= 12'b001000101101;
   29892: result <= 12'b001000101101;
   29893: result <= 12'b001000101101;
   29894: result <= 12'b001000101101;
   29895: result <= 12'b001000101101;
   29896: result <= 12'b001000101100;
   29897: result <= 12'b001000101100;
   29898: result <= 12'b001000101100;
   29899: result <= 12'b001000101100;
   29900: result <= 12'b001000101100;
   29901: result <= 12'b001000101011;
   29902: result <= 12'b001000101011;
   29903: result <= 12'b001000101011;
   29904: result <= 12'b001000101011;
   29905: result <= 12'b001000101011;
   29906: result <= 12'b001000101010;
   29907: result <= 12'b001000101010;
   29908: result <= 12'b001000101010;
   29909: result <= 12'b001000101010;
   29910: result <= 12'b001000101010;
   29911: result <= 12'b001000101001;
   29912: result <= 12'b001000101001;
   29913: result <= 12'b001000101001;
   29914: result <= 12'b001000101001;
   29915: result <= 12'b001000101001;
   29916: result <= 12'b001000101001;
   29917: result <= 12'b001000101000;
   29918: result <= 12'b001000101000;
   29919: result <= 12'b001000101000;
   29920: result <= 12'b001000101000;
   29921: result <= 12'b001000101000;
   29922: result <= 12'b001000100111;
   29923: result <= 12'b001000100111;
   29924: result <= 12'b001000100111;
   29925: result <= 12'b001000100111;
   29926: result <= 12'b001000100111;
   29927: result <= 12'b001000100110;
   29928: result <= 12'b001000100110;
   29929: result <= 12'b001000100110;
   29930: result <= 12'b001000100110;
   29931: result <= 12'b001000100110;
   29932: result <= 12'b001000100110;
   29933: result <= 12'b001000100101;
   29934: result <= 12'b001000100101;
   29935: result <= 12'b001000100101;
   29936: result <= 12'b001000100101;
   29937: result <= 12'b001000100101;
   29938: result <= 12'b001000100100;
   29939: result <= 12'b001000100100;
   29940: result <= 12'b001000100100;
   29941: result <= 12'b001000100100;
   29942: result <= 12'b001000100100;
   29943: result <= 12'b001000100011;
   29944: result <= 12'b001000100011;
   29945: result <= 12'b001000100011;
   29946: result <= 12'b001000100011;
   29947: result <= 12'b001000100011;
   29948: result <= 12'b001000100010;
   29949: result <= 12'b001000100010;
   29950: result <= 12'b001000100010;
   29951: result <= 12'b001000100010;
   29952: result <= 12'b001000100010;
   29953: result <= 12'b001000100010;
   29954: result <= 12'b001000100001;
   29955: result <= 12'b001000100001;
   29956: result <= 12'b001000100001;
   29957: result <= 12'b001000100001;
   29958: result <= 12'b001000100001;
   29959: result <= 12'b001000100000;
   29960: result <= 12'b001000100000;
   29961: result <= 12'b001000100000;
   29962: result <= 12'b001000100000;
   29963: result <= 12'b001000100000;
   29964: result <= 12'b001000011111;
   29965: result <= 12'b001000011111;
   29966: result <= 12'b001000011111;
   29967: result <= 12'b001000011111;
   29968: result <= 12'b001000011111;
   29969: result <= 12'b001000011111;
   29970: result <= 12'b001000011110;
   29971: result <= 12'b001000011110;
   29972: result <= 12'b001000011110;
   29973: result <= 12'b001000011110;
   29974: result <= 12'b001000011110;
   29975: result <= 12'b001000011101;
   29976: result <= 12'b001000011101;
   29977: result <= 12'b001000011101;
   29978: result <= 12'b001000011101;
   29979: result <= 12'b001000011101;
   29980: result <= 12'b001000011100;
   29981: result <= 12'b001000011100;
   29982: result <= 12'b001000011100;
   29983: result <= 12'b001000011100;
   29984: result <= 12'b001000011100;
   29985: result <= 12'b001000011011;
   29986: result <= 12'b001000011011;
   29987: result <= 12'b001000011011;
   29988: result <= 12'b001000011011;
   29989: result <= 12'b001000011011;
   29990: result <= 12'b001000011011;
   29991: result <= 12'b001000011010;
   29992: result <= 12'b001000011010;
   29993: result <= 12'b001000011010;
   29994: result <= 12'b001000011010;
   29995: result <= 12'b001000011010;
   29996: result <= 12'b001000011001;
   29997: result <= 12'b001000011001;
   29998: result <= 12'b001000011001;
   29999: result <= 12'b001000011001;
   30000: result <= 12'b001000011001;
   30001: result <= 12'b001000011000;
   30002: result <= 12'b001000011000;
   30003: result <= 12'b001000011000;
   30004: result <= 12'b001000011000;
   30005: result <= 12'b001000011000;
   30006: result <= 12'b001000011000;
   30007: result <= 12'b001000010111;
   30008: result <= 12'b001000010111;
   30009: result <= 12'b001000010111;
   30010: result <= 12'b001000010111;
   30011: result <= 12'b001000010111;
   30012: result <= 12'b001000010110;
   30013: result <= 12'b001000010110;
   30014: result <= 12'b001000010110;
   30015: result <= 12'b001000010110;
   30016: result <= 12'b001000010110;
   30017: result <= 12'b001000010101;
   30018: result <= 12'b001000010101;
   30019: result <= 12'b001000010101;
   30020: result <= 12'b001000010101;
   30021: result <= 12'b001000010101;
   30022: result <= 12'b001000010100;
   30023: result <= 12'b001000010100;
   30024: result <= 12'b001000010100;
   30025: result <= 12'b001000010100;
   30026: result <= 12'b001000010100;
   30027: result <= 12'b001000010100;
   30028: result <= 12'b001000010011;
   30029: result <= 12'b001000010011;
   30030: result <= 12'b001000010011;
   30031: result <= 12'b001000010011;
   30032: result <= 12'b001000010011;
   30033: result <= 12'b001000010010;
   30034: result <= 12'b001000010010;
   30035: result <= 12'b001000010010;
   30036: result <= 12'b001000010010;
   30037: result <= 12'b001000010010;
   30038: result <= 12'b001000010001;
   30039: result <= 12'b001000010001;
   30040: result <= 12'b001000010001;
   30041: result <= 12'b001000010001;
   30042: result <= 12'b001000010001;
   30043: result <= 12'b001000010000;
   30044: result <= 12'b001000010000;
   30045: result <= 12'b001000010000;
   30046: result <= 12'b001000010000;
   30047: result <= 12'b001000010000;
   30048: result <= 12'b001000010000;
   30049: result <= 12'b001000001111;
   30050: result <= 12'b001000001111;
   30051: result <= 12'b001000001111;
   30052: result <= 12'b001000001111;
   30053: result <= 12'b001000001111;
   30054: result <= 12'b001000001110;
   30055: result <= 12'b001000001110;
   30056: result <= 12'b001000001110;
   30057: result <= 12'b001000001110;
   30058: result <= 12'b001000001110;
   30059: result <= 12'b001000001101;
   30060: result <= 12'b001000001101;
   30061: result <= 12'b001000001101;
   30062: result <= 12'b001000001101;
   30063: result <= 12'b001000001101;
   30064: result <= 12'b001000001101;
   30065: result <= 12'b001000001100;
   30066: result <= 12'b001000001100;
   30067: result <= 12'b001000001100;
   30068: result <= 12'b001000001100;
   30069: result <= 12'b001000001100;
   30070: result <= 12'b001000001011;
   30071: result <= 12'b001000001011;
   30072: result <= 12'b001000001011;
   30073: result <= 12'b001000001011;
   30074: result <= 12'b001000001011;
   30075: result <= 12'b001000001010;
   30076: result <= 12'b001000001010;
   30077: result <= 12'b001000001010;
   30078: result <= 12'b001000001010;
   30079: result <= 12'b001000001010;
   30080: result <= 12'b001000001001;
   30081: result <= 12'b001000001001;
   30082: result <= 12'b001000001001;
   30083: result <= 12'b001000001001;
   30084: result <= 12'b001000001001;
   30085: result <= 12'b001000001001;
   30086: result <= 12'b001000001000;
   30087: result <= 12'b001000001000;
   30088: result <= 12'b001000001000;
   30089: result <= 12'b001000001000;
   30090: result <= 12'b001000001000;
   30091: result <= 12'b001000000111;
   30092: result <= 12'b001000000111;
   30093: result <= 12'b001000000111;
   30094: result <= 12'b001000000111;
   30095: result <= 12'b001000000111;
   30096: result <= 12'b001000000110;
   30097: result <= 12'b001000000110;
   30098: result <= 12'b001000000110;
   30099: result <= 12'b001000000110;
   30100: result <= 12'b001000000110;
   30101: result <= 12'b001000000101;
   30102: result <= 12'b001000000101;
   30103: result <= 12'b001000000101;
   30104: result <= 12'b001000000101;
   30105: result <= 12'b001000000101;
   30106: result <= 12'b001000000101;
   30107: result <= 12'b001000000100;
   30108: result <= 12'b001000000100;
   30109: result <= 12'b001000000100;
   30110: result <= 12'b001000000100;
   30111: result <= 12'b001000000100;
   30112: result <= 12'b001000000011;
   30113: result <= 12'b001000000011;
   30114: result <= 12'b001000000011;
   30115: result <= 12'b001000000011;
   30116: result <= 12'b001000000011;
   30117: result <= 12'b001000000010;
   30118: result <= 12'b001000000010;
   30119: result <= 12'b001000000010;
   30120: result <= 12'b001000000010;
   30121: result <= 12'b001000000010;
   30122: result <= 12'b001000000001;
   30123: result <= 12'b001000000001;
   30124: result <= 12'b001000000001;
   30125: result <= 12'b001000000001;
   30126: result <= 12'b001000000001;
   30127: result <= 12'b001000000001;
   30128: result <= 12'b001000000000;
   30129: result <= 12'b001000000000;
   30130: result <= 12'b001000000000;
   30131: result <= 12'b001000000000;
   30132: result <= 12'b001000000000;
   30133: result <= 12'b000111111111;
   30134: result <= 12'b000111111111;
   30135: result <= 12'b000111111111;
   30136: result <= 12'b000111111111;
   30137: result <= 12'b000111111111;
   30138: result <= 12'b000111111110;
   30139: result <= 12'b000111111110;
   30140: result <= 12'b000111111110;
   30141: result <= 12'b000111111110;
   30142: result <= 12'b000111111110;
   30143: result <= 12'b000111111101;
   30144: result <= 12'b000111111101;
   30145: result <= 12'b000111111101;
   30146: result <= 12'b000111111101;
   30147: result <= 12'b000111111101;
   30148: result <= 12'b000111111101;
   30149: result <= 12'b000111111100;
   30150: result <= 12'b000111111100;
   30151: result <= 12'b000111111100;
   30152: result <= 12'b000111111100;
   30153: result <= 12'b000111111100;
   30154: result <= 12'b000111111011;
   30155: result <= 12'b000111111011;
   30156: result <= 12'b000111111011;
   30157: result <= 12'b000111111011;
   30158: result <= 12'b000111111011;
   30159: result <= 12'b000111111010;
   30160: result <= 12'b000111111010;
   30161: result <= 12'b000111111010;
   30162: result <= 12'b000111111010;
   30163: result <= 12'b000111111010;
   30164: result <= 12'b000111111001;
   30165: result <= 12'b000111111001;
   30166: result <= 12'b000111111001;
   30167: result <= 12'b000111111001;
   30168: result <= 12'b000111111001;
   30169: result <= 12'b000111111001;
   30170: result <= 12'b000111111000;
   30171: result <= 12'b000111111000;
   30172: result <= 12'b000111111000;
   30173: result <= 12'b000111111000;
   30174: result <= 12'b000111111000;
   30175: result <= 12'b000111110111;
   30176: result <= 12'b000111110111;
   30177: result <= 12'b000111110111;
   30178: result <= 12'b000111110111;
   30179: result <= 12'b000111110111;
   30180: result <= 12'b000111110110;
   30181: result <= 12'b000111110110;
   30182: result <= 12'b000111110110;
   30183: result <= 12'b000111110110;
   30184: result <= 12'b000111110110;
   30185: result <= 12'b000111110110;
   30186: result <= 12'b000111110101;
   30187: result <= 12'b000111110101;
   30188: result <= 12'b000111110101;
   30189: result <= 12'b000111110101;
   30190: result <= 12'b000111110101;
   30191: result <= 12'b000111110100;
   30192: result <= 12'b000111110100;
   30193: result <= 12'b000111110100;
   30194: result <= 12'b000111110100;
   30195: result <= 12'b000111110100;
   30196: result <= 12'b000111110011;
   30197: result <= 12'b000111110011;
   30198: result <= 12'b000111110011;
   30199: result <= 12'b000111110011;
   30200: result <= 12'b000111110011;
   30201: result <= 12'b000111110010;
   30202: result <= 12'b000111110010;
   30203: result <= 12'b000111110010;
   30204: result <= 12'b000111110010;
   30205: result <= 12'b000111110010;
   30206: result <= 12'b000111110010;
   30207: result <= 12'b000111110001;
   30208: result <= 12'b000111110001;
   30209: result <= 12'b000111110001;
   30210: result <= 12'b000111110001;
   30211: result <= 12'b000111110001;
   30212: result <= 12'b000111110000;
   30213: result <= 12'b000111110000;
   30214: result <= 12'b000111110000;
   30215: result <= 12'b000111110000;
   30216: result <= 12'b000111110000;
   30217: result <= 12'b000111101111;
   30218: result <= 12'b000111101111;
   30219: result <= 12'b000111101111;
   30220: result <= 12'b000111101111;
   30221: result <= 12'b000111101111;
   30222: result <= 12'b000111101110;
   30223: result <= 12'b000111101110;
   30224: result <= 12'b000111101110;
   30225: result <= 12'b000111101110;
   30226: result <= 12'b000111101110;
   30227: result <= 12'b000111101110;
   30228: result <= 12'b000111101101;
   30229: result <= 12'b000111101101;
   30230: result <= 12'b000111101101;
   30231: result <= 12'b000111101101;
   30232: result <= 12'b000111101101;
   30233: result <= 12'b000111101100;
   30234: result <= 12'b000111101100;
   30235: result <= 12'b000111101100;
   30236: result <= 12'b000111101100;
   30237: result <= 12'b000111101100;
   30238: result <= 12'b000111101011;
   30239: result <= 12'b000111101011;
   30240: result <= 12'b000111101011;
   30241: result <= 12'b000111101011;
   30242: result <= 12'b000111101011;
   30243: result <= 12'b000111101010;
   30244: result <= 12'b000111101010;
   30245: result <= 12'b000111101010;
   30246: result <= 12'b000111101010;
   30247: result <= 12'b000111101010;
   30248: result <= 12'b000111101010;
   30249: result <= 12'b000111101001;
   30250: result <= 12'b000111101001;
   30251: result <= 12'b000111101001;
   30252: result <= 12'b000111101001;
   30253: result <= 12'b000111101001;
   30254: result <= 12'b000111101000;
   30255: result <= 12'b000111101000;
   30256: result <= 12'b000111101000;
   30257: result <= 12'b000111101000;
   30258: result <= 12'b000111101000;
   30259: result <= 12'b000111100111;
   30260: result <= 12'b000111100111;
   30261: result <= 12'b000111100111;
   30262: result <= 12'b000111100111;
   30263: result <= 12'b000111100111;
   30264: result <= 12'b000111100110;
   30265: result <= 12'b000111100110;
   30266: result <= 12'b000111100110;
   30267: result <= 12'b000111100110;
   30268: result <= 12'b000111100110;
   30269: result <= 12'b000111100101;
   30270: result <= 12'b000111100101;
   30271: result <= 12'b000111100101;
   30272: result <= 12'b000111100101;
   30273: result <= 12'b000111100101;
   30274: result <= 12'b000111100101;
   30275: result <= 12'b000111100100;
   30276: result <= 12'b000111100100;
   30277: result <= 12'b000111100100;
   30278: result <= 12'b000111100100;
   30279: result <= 12'b000111100100;
   30280: result <= 12'b000111100011;
   30281: result <= 12'b000111100011;
   30282: result <= 12'b000111100011;
   30283: result <= 12'b000111100011;
   30284: result <= 12'b000111100011;
   30285: result <= 12'b000111100010;
   30286: result <= 12'b000111100010;
   30287: result <= 12'b000111100010;
   30288: result <= 12'b000111100010;
   30289: result <= 12'b000111100010;
   30290: result <= 12'b000111100001;
   30291: result <= 12'b000111100001;
   30292: result <= 12'b000111100001;
   30293: result <= 12'b000111100001;
   30294: result <= 12'b000111100001;
   30295: result <= 12'b000111100001;
   30296: result <= 12'b000111100000;
   30297: result <= 12'b000111100000;
   30298: result <= 12'b000111100000;
   30299: result <= 12'b000111100000;
   30300: result <= 12'b000111100000;
   30301: result <= 12'b000111011111;
   30302: result <= 12'b000111011111;
   30303: result <= 12'b000111011111;
   30304: result <= 12'b000111011111;
   30305: result <= 12'b000111011111;
   30306: result <= 12'b000111011110;
   30307: result <= 12'b000111011110;
   30308: result <= 12'b000111011110;
   30309: result <= 12'b000111011110;
   30310: result <= 12'b000111011110;
   30311: result <= 12'b000111011101;
   30312: result <= 12'b000111011101;
   30313: result <= 12'b000111011101;
   30314: result <= 12'b000111011101;
   30315: result <= 12'b000111011101;
   30316: result <= 12'b000111011101;
   30317: result <= 12'b000111011100;
   30318: result <= 12'b000111011100;
   30319: result <= 12'b000111011100;
   30320: result <= 12'b000111011100;
   30321: result <= 12'b000111011100;
   30322: result <= 12'b000111011011;
   30323: result <= 12'b000111011011;
   30324: result <= 12'b000111011011;
   30325: result <= 12'b000111011011;
   30326: result <= 12'b000111011011;
   30327: result <= 12'b000111011010;
   30328: result <= 12'b000111011010;
   30329: result <= 12'b000111011010;
   30330: result <= 12'b000111011010;
   30331: result <= 12'b000111011010;
   30332: result <= 12'b000111011001;
   30333: result <= 12'b000111011001;
   30334: result <= 12'b000111011001;
   30335: result <= 12'b000111011001;
   30336: result <= 12'b000111011001;
   30337: result <= 12'b000111011001;
   30338: result <= 12'b000111011000;
   30339: result <= 12'b000111011000;
   30340: result <= 12'b000111011000;
   30341: result <= 12'b000111011000;
   30342: result <= 12'b000111011000;
   30343: result <= 12'b000111010111;
   30344: result <= 12'b000111010111;
   30345: result <= 12'b000111010111;
   30346: result <= 12'b000111010111;
   30347: result <= 12'b000111010111;
   30348: result <= 12'b000111010110;
   30349: result <= 12'b000111010110;
   30350: result <= 12'b000111010110;
   30351: result <= 12'b000111010110;
   30352: result <= 12'b000111010110;
   30353: result <= 12'b000111010101;
   30354: result <= 12'b000111010101;
   30355: result <= 12'b000111010101;
   30356: result <= 12'b000111010101;
   30357: result <= 12'b000111010101;
   30358: result <= 12'b000111010101;
   30359: result <= 12'b000111010100;
   30360: result <= 12'b000111010100;
   30361: result <= 12'b000111010100;
   30362: result <= 12'b000111010100;
   30363: result <= 12'b000111010100;
   30364: result <= 12'b000111010011;
   30365: result <= 12'b000111010011;
   30366: result <= 12'b000111010011;
   30367: result <= 12'b000111010011;
   30368: result <= 12'b000111010011;
   30369: result <= 12'b000111010010;
   30370: result <= 12'b000111010010;
   30371: result <= 12'b000111010010;
   30372: result <= 12'b000111010010;
   30373: result <= 12'b000111010010;
   30374: result <= 12'b000111010001;
   30375: result <= 12'b000111010001;
   30376: result <= 12'b000111010001;
   30377: result <= 12'b000111010001;
   30378: result <= 12'b000111010001;
   30379: result <= 12'b000111010000;
   30380: result <= 12'b000111010000;
   30381: result <= 12'b000111010000;
   30382: result <= 12'b000111010000;
   30383: result <= 12'b000111010000;
   30384: result <= 12'b000111010000;
   30385: result <= 12'b000111001111;
   30386: result <= 12'b000111001111;
   30387: result <= 12'b000111001111;
   30388: result <= 12'b000111001111;
   30389: result <= 12'b000111001111;
   30390: result <= 12'b000111001110;
   30391: result <= 12'b000111001110;
   30392: result <= 12'b000111001110;
   30393: result <= 12'b000111001110;
   30394: result <= 12'b000111001110;
   30395: result <= 12'b000111001101;
   30396: result <= 12'b000111001101;
   30397: result <= 12'b000111001101;
   30398: result <= 12'b000111001101;
   30399: result <= 12'b000111001101;
   30400: result <= 12'b000111001100;
   30401: result <= 12'b000111001100;
   30402: result <= 12'b000111001100;
   30403: result <= 12'b000111001100;
   30404: result <= 12'b000111001100;
   30405: result <= 12'b000111001100;
   30406: result <= 12'b000111001011;
   30407: result <= 12'b000111001011;
   30408: result <= 12'b000111001011;
   30409: result <= 12'b000111001011;
   30410: result <= 12'b000111001011;
   30411: result <= 12'b000111001010;
   30412: result <= 12'b000111001010;
   30413: result <= 12'b000111001010;
   30414: result <= 12'b000111001010;
   30415: result <= 12'b000111001010;
   30416: result <= 12'b000111001001;
   30417: result <= 12'b000111001001;
   30418: result <= 12'b000111001001;
   30419: result <= 12'b000111001001;
   30420: result <= 12'b000111001001;
   30421: result <= 12'b000111001000;
   30422: result <= 12'b000111001000;
   30423: result <= 12'b000111001000;
   30424: result <= 12'b000111001000;
   30425: result <= 12'b000111001000;
   30426: result <= 12'b000111000111;
   30427: result <= 12'b000111000111;
   30428: result <= 12'b000111000111;
   30429: result <= 12'b000111000111;
   30430: result <= 12'b000111000111;
   30431: result <= 12'b000111000111;
   30432: result <= 12'b000111000110;
   30433: result <= 12'b000111000110;
   30434: result <= 12'b000111000110;
   30435: result <= 12'b000111000110;
   30436: result <= 12'b000111000110;
   30437: result <= 12'b000111000101;
   30438: result <= 12'b000111000101;
   30439: result <= 12'b000111000101;
   30440: result <= 12'b000111000101;
   30441: result <= 12'b000111000101;
   30442: result <= 12'b000111000100;
   30443: result <= 12'b000111000100;
   30444: result <= 12'b000111000100;
   30445: result <= 12'b000111000100;
   30446: result <= 12'b000111000100;
   30447: result <= 12'b000111000011;
   30448: result <= 12'b000111000011;
   30449: result <= 12'b000111000011;
   30450: result <= 12'b000111000011;
   30451: result <= 12'b000111000011;
   30452: result <= 12'b000111000011;
   30453: result <= 12'b000111000010;
   30454: result <= 12'b000111000010;
   30455: result <= 12'b000111000010;
   30456: result <= 12'b000111000010;
   30457: result <= 12'b000111000010;
   30458: result <= 12'b000111000001;
   30459: result <= 12'b000111000001;
   30460: result <= 12'b000111000001;
   30461: result <= 12'b000111000001;
   30462: result <= 12'b000111000001;
   30463: result <= 12'b000111000000;
   30464: result <= 12'b000111000000;
   30465: result <= 12'b000111000000;
   30466: result <= 12'b000111000000;
   30467: result <= 12'b000111000000;
   30468: result <= 12'b000110111111;
   30469: result <= 12'b000110111111;
   30470: result <= 12'b000110111111;
   30471: result <= 12'b000110111111;
   30472: result <= 12'b000110111111;
   30473: result <= 12'b000110111110;
   30474: result <= 12'b000110111110;
   30475: result <= 12'b000110111110;
   30476: result <= 12'b000110111110;
   30477: result <= 12'b000110111110;
   30478: result <= 12'b000110111110;
   30479: result <= 12'b000110111101;
   30480: result <= 12'b000110111101;
   30481: result <= 12'b000110111101;
   30482: result <= 12'b000110111101;
   30483: result <= 12'b000110111101;
   30484: result <= 12'b000110111100;
   30485: result <= 12'b000110111100;
   30486: result <= 12'b000110111100;
   30487: result <= 12'b000110111100;
   30488: result <= 12'b000110111100;
   30489: result <= 12'b000110111011;
   30490: result <= 12'b000110111011;
   30491: result <= 12'b000110111011;
   30492: result <= 12'b000110111011;
   30493: result <= 12'b000110111011;
   30494: result <= 12'b000110111010;
   30495: result <= 12'b000110111010;
   30496: result <= 12'b000110111010;
   30497: result <= 12'b000110111010;
   30498: result <= 12'b000110111010;
   30499: result <= 12'b000110111010;
   30500: result <= 12'b000110111001;
   30501: result <= 12'b000110111001;
   30502: result <= 12'b000110111001;
   30503: result <= 12'b000110111001;
   30504: result <= 12'b000110111001;
   30505: result <= 12'b000110111000;
   30506: result <= 12'b000110111000;
   30507: result <= 12'b000110111000;
   30508: result <= 12'b000110111000;
   30509: result <= 12'b000110111000;
   30510: result <= 12'b000110110111;
   30511: result <= 12'b000110110111;
   30512: result <= 12'b000110110111;
   30513: result <= 12'b000110110111;
   30514: result <= 12'b000110110111;
   30515: result <= 12'b000110110110;
   30516: result <= 12'b000110110110;
   30517: result <= 12'b000110110110;
   30518: result <= 12'b000110110110;
   30519: result <= 12'b000110110110;
   30520: result <= 12'b000110110101;
   30521: result <= 12'b000110110101;
   30522: result <= 12'b000110110101;
   30523: result <= 12'b000110110101;
   30524: result <= 12'b000110110101;
   30525: result <= 12'b000110110101;
   30526: result <= 12'b000110110100;
   30527: result <= 12'b000110110100;
   30528: result <= 12'b000110110100;
   30529: result <= 12'b000110110100;
   30530: result <= 12'b000110110100;
   30531: result <= 12'b000110110011;
   30532: result <= 12'b000110110011;
   30533: result <= 12'b000110110011;
   30534: result <= 12'b000110110011;
   30535: result <= 12'b000110110011;
   30536: result <= 12'b000110110010;
   30537: result <= 12'b000110110010;
   30538: result <= 12'b000110110010;
   30539: result <= 12'b000110110010;
   30540: result <= 12'b000110110010;
   30541: result <= 12'b000110110001;
   30542: result <= 12'b000110110001;
   30543: result <= 12'b000110110001;
   30544: result <= 12'b000110110001;
   30545: result <= 12'b000110110001;
   30546: result <= 12'b000110110000;
   30547: result <= 12'b000110110000;
   30548: result <= 12'b000110110000;
   30549: result <= 12'b000110110000;
   30550: result <= 12'b000110110000;
   30551: result <= 12'b000110110000;
   30552: result <= 12'b000110101111;
   30553: result <= 12'b000110101111;
   30554: result <= 12'b000110101111;
   30555: result <= 12'b000110101111;
   30556: result <= 12'b000110101111;
   30557: result <= 12'b000110101110;
   30558: result <= 12'b000110101110;
   30559: result <= 12'b000110101110;
   30560: result <= 12'b000110101110;
   30561: result <= 12'b000110101110;
   30562: result <= 12'b000110101101;
   30563: result <= 12'b000110101101;
   30564: result <= 12'b000110101101;
   30565: result <= 12'b000110101101;
   30566: result <= 12'b000110101101;
   30567: result <= 12'b000110101100;
   30568: result <= 12'b000110101100;
   30569: result <= 12'b000110101100;
   30570: result <= 12'b000110101100;
   30571: result <= 12'b000110101100;
   30572: result <= 12'b000110101100;
   30573: result <= 12'b000110101011;
   30574: result <= 12'b000110101011;
   30575: result <= 12'b000110101011;
   30576: result <= 12'b000110101011;
   30577: result <= 12'b000110101011;
   30578: result <= 12'b000110101010;
   30579: result <= 12'b000110101010;
   30580: result <= 12'b000110101010;
   30581: result <= 12'b000110101010;
   30582: result <= 12'b000110101010;
   30583: result <= 12'b000110101001;
   30584: result <= 12'b000110101001;
   30585: result <= 12'b000110101001;
   30586: result <= 12'b000110101001;
   30587: result <= 12'b000110101001;
   30588: result <= 12'b000110101000;
   30589: result <= 12'b000110101000;
   30590: result <= 12'b000110101000;
   30591: result <= 12'b000110101000;
   30592: result <= 12'b000110101000;
   30593: result <= 12'b000110100111;
   30594: result <= 12'b000110100111;
   30595: result <= 12'b000110100111;
   30596: result <= 12'b000110100111;
   30597: result <= 12'b000110100111;
   30598: result <= 12'b000110100111;
   30599: result <= 12'b000110100110;
   30600: result <= 12'b000110100110;
   30601: result <= 12'b000110100110;
   30602: result <= 12'b000110100110;
   30603: result <= 12'b000110100110;
   30604: result <= 12'b000110100101;
   30605: result <= 12'b000110100101;
   30606: result <= 12'b000110100101;
   30607: result <= 12'b000110100101;
   30608: result <= 12'b000110100101;
   30609: result <= 12'b000110100100;
   30610: result <= 12'b000110100100;
   30611: result <= 12'b000110100100;
   30612: result <= 12'b000110100100;
   30613: result <= 12'b000110100100;
   30614: result <= 12'b000110100011;
   30615: result <= 12'b000110100011;
   30616: result <= 12'b000110100011;
   30617: result <= 12'b000110100011;
   30618: result <= 12'b000110100011;
   30619: result <= 12'b000110100010;
   30620: result <= 12'b000110100010;
   30621: result <= 12'b000110100010;
   30622: result <= 12'b000110100010;
   30623: result <= 12'b000110100010;
   30624: result <= 12'b000110100010;
   30625: result <= 12'b000110100001;
   30626: result <= 12'b000110100001;
   30627: result <= 12'b000110100001;
   30628: result <= 12'b000110100001;
   30629: result <= 12'b000110100001;
   30630: result <= 12'b000110100000;
   30631: result <= 12'b000110100000;
   30632: result <= 12'b000110100000;
   30633: result <= 12'b000110100000;
   30634: result <= 12'b000110100000;
   30635: result <= 12'b000110011111;
   30636: result <= 12'b000110011111;
   30637: result <= 12'b000110011111;
   30638: result <= 12'b000110011111;
   30639: result <= 12'b000110011111;
   30640: result <= 12'b000110011110;
   30641: result <= 12'b000110011110;
   30642: result <= 12'b000110011110;
   30643: result <= 12'b000110011110;
   30644: result <= 12'b000110011110;
   30645: result <= 12'b000110011101;
   30646: result <= 12'b000110011101;
   30647: result <= 12'b000110011101;
   30648: result <= 12'b000110011101;
   30649: result <= 12'b000110011101;
   30650: result <= 12'b000110011101;
   30651: result <= 12'b000110011100;
   30652: result <= 12'b000110011100;
   30653: result <= 12'b000110011100;
   30654: result <= 12'b000110011100;
   30655: result <= 12'b000110011100;
   30656: result <= 12'b000110011011;
   30657: result <= 12'b000110011011;
   30658: result <= 12'b000110011011;
   30659: result <= 12'b000110011011;
   30660: result <= 12'b000110011011;
   30661: result <= 12'b000110011010;
   30662: result <= 12'b000110011010;
   30663: result <= 12'b000110011010;
   30664: result <= 12'b000110011010;
   30665: result <= 12'b000110011010;
   30666: result <= 12'b000110011001;
   30667: result <= 12'b000110011001;
   30668: result <= 12'b000110011001;
   30669: result <= 12'b000110011001;
   30670: result <= 12'b000110011001;
   30671: result <= 12'b000110011000;
   30672: result <= 12'b000110011000;
   30673: result <= 12'b000110011000;
   30674: result <= 12'b000110011000;
   30675: result <= 12'b000110011000;
   30676: result <= 12'b000110011000;
   30677: result <= 12'b000110010111;
   30678: result <= 12'b000110010111;
   30679: result <= 12'b000110010111;
   30680: result <= 12'b000110010111;
   30681: result <= 12'b000110010111;
   30682: result <= 12'b000110010110;
   30683: result <= 12'b000110010110;
   30684: result <= 12'b000110010110;
   30685: result <= 12'b000110010110;
   30686: result <= 12'b000110010110;
   30687: result <= 12'b000110010101;
   30688: result <= 12'b000110010101;
   30689: result <= 12'b000110010101;
   30690: result <= 12'b000110010101;
   30691: result <= 12'b000110010101;
   30692: result <= 12'b000110010100;
   30693: result <= 12'b000110010100;
   30694: result <= 12'b000110010100;
   30695: result <= 12'b000110010100;
   30696: result <= 12'b000110010100;
   30697: result <= 12'b000110010011;
   30698: result <= 12'b000110010011;
   30699: result <= 12'b000110010011;
   30700: result <= 12'b000110010011;
   30701: result <= 12'b000110010011;
   30702: result <= 12'b000110010011;
   30703: result <= 12'b000110010010;
   30704: result <= 12'b000110010010;
   30705: result <= 12'b000110010010;
   30706: result <= 12'b000110010010;
   30707: result <= 12'b000110010010;
   30708: result <= 12'b000110010001;
   30709: result <= 12'b000110010001;
   30710: result <= 12'b000110010001;
   30711: result <= 12'b000110010001;
   30712: result <= 12'b000110010001;
   30713: result <= 12'b000110010000;
   30714: result <= 12'b000110010000;
   30715: result <= 12'b000110010000;
   30716: result <= 12'b000110010000;
   30717: result <= 12'b000110010000;
   30718: result <= 12'b000110001111;
   30719: result <= 12'b000110001111;
   30720: result <= 12'b000110001111;
   30721: result <= 12'b000110001111;
   30722: result <= 12'b000110001111;
   30723: result <= 12'b000110001110;
   30724: result <= 12'b000110001110;
   30725: result <= 12'b000110001110;
   30726: result <= 12'b000110001110;
   30727: result <= 12'b000110001110;
   30728: result <= 12'b000110001110;
   30729: result <= 12'b000110001101;
   30730: result <= 12'b000110001101;
   30731: result <= 12'b000110001101;
   30732: result <= 12'b000110001101;
   30733: result <= 12'b000110001101;
   30734: result <= 12'b000110001100;
   30735: result <= 12'b000110001100;
   30736: result <= 12'b000110001100;
   30737: result <= 12'b000110001100;
   30738: result <= 12'b000110001100;
   30739: result <= 12'b000110001011;
   30740: result <= 12'b000110001011;
   30741: result <= 12'b000110001011;
   30742: result <= 12'b000110001011;
   30743: result <= 12'b000110001011;
   30744: result <= 12'b000110001010;
   30745: result <= 12'b000110001010;
   30746: result <= 12'b000110001010;
   30747: result <= 12'b000110001010;
   30748: result <= 12'b000110001010;
   30749: result <= 12'b000110001001;
   30750: result <= 12'b000110001001;
   30751: result <= 12'b000110001001;
   30752: result <= 12'b000110001001;
   30753: result <= 12'b000110001001;
   30754: result <= 12'b000110001000;
   30755: result <= 12'b000110001000;
   30756: result <= 12'b000110001000;
   30757: result <= 12'b000110001000;
   30758: result <= 12'b000110001000;
   30759: result <= 12'b000110001000;
   30760: result <= 12'b000110000111;
   30761: result <= 12'b000110000111;
   30762: result <= 12'b000110000111;
   30763: result <= 12'b000110000111;
   30764: result <= 12'b000110000111;
   30765: result <= 12'b000110000110;
   30766: result <= 12'b000110000110;
   30767: result <= 12'b000110000110;
   30768: result <= 12'b000110000110;
   30769: result <= 12'b000110000110;
   30770: result <= 12'b000110000101;
   30771: result <= 12'b000110000101;
   30772: result <= 12'b000110000101;
   30773: result <= 12'b000110000101;
   30774: result <= 12'b000110000101;
   30775: result <= 12'b000110000100;
   30776: result <= 12'b000110000100;
   30777: result <= 12'b000110000100;
   30778: result <= 12'b000110000100;
   30779: result <= 12'b000110000100;
   30780: result <= 12'b000110000011;
   30781: result <= 12'b000110000011;
   30782: result <= 12'b000110000011;
   30783: result <= 12'b000110000011;
   30784: result <= 12'b000110000011;
   30785: result <= 12'b000110000011;
   30786: result <= 12'b000110000010;
   30787: result <= 12'b000110000010;
   30788: result <= 12'b000110000010;
   30789: result <= 12'b000110000010;
   30790: result <= 12'b000110000010;
   30791: result <= 12'b000110000001;
   30792: result <= 12'b000110000001;
   30793: result <= 12'b000110000001;
   30794: result <= 12'b000110000001;
   30795: result <= 12'b000110000001;
   30796: result <= 12'b000110000000;
   30797: result <= 12'b000110000000;
   30798: result <= 12'b000110000000;
   30799: result <= 12'b000110000000;
   30800: result <= 12'b000110000000;
   30801: result <= 12'b000101111111;
   30802: result <= 12'b000101111111;
   30803: result <= 12'b000101111111;
   30804: result <= 12'b000101111111;
   30805: result <= 12'b000101111111;
   30806: result <= 12'b000101111110;
   30807: result <= 12'b000101111110;
   30808: result <= 12'b000101111110;
   30809: result <= 12'b000101111110;
   30810: result <= 12'b000101111110;
   30811: result <= 12'b000101111110;
   30812: result <= 12'b000101111101;
   30813: result <= 12'b000101111101;
   30814: result <= 12'b000101111101;
   30815: result <= 12'b000101111101;
   30816: result <= 12'b000101111101;
   30817: result <= 12'b000101111100;
   30818: result <= 12'b000101111100;
   30819: result <= 12'b000101111100;
   30820: result <= 12'b000101111100;
   30821: result <= 12'b000101111100;
   30822: result <= 12'b000101111011;
   30823: result <= 12'b000101111011;
   30824: result <= 12'b000101111011;
   30825: result <= 12'b000101111011;
   30826: result <= 12'b000101111011;
   30827: result <= 12'b000101111010;
   30828: result <= 12'b000101111010;
   30829: result <= 12'b000101111010;
   30830: result <= 12'b000101111010;
   30831: result <= 12'b000101111010;
   30832: result <= 12'b000101111001;
   30833: result <= 12'b000101111001;
   30834: result <= 12'b000101111001;
   30835: result <= 12'b000101111001;
   30836: result <= 12'b000101111001;
   30837: result <= 12'b000101111000;
   30838: result <= 12'b000101111000;
   30839: result <= 12'b000101111000;
   30840: result <= 12'b000101111000;
   30841: result <= 12'b000101111000;
   30842: result <= 12'b000101111000;
   30843: result <= 12'b000101110111;
   30844: result <= 12'b000101110111;
   30845: result <= 12'b000101110111;
   30846: result <= 12'b000101110111;
   30847: result <= 12'b000101110111;
   30848: result <= 12'b000101110110;
   30849: result <= 12'b000101110110;
   30850: result <= 12'b000101110110;
   30851: result <= 12'b000101110110;
   30852: result <= 12'b000101110110;
   30853: result <= 12'b000101110101;
   30854: result <= 12'b000101110101;
   30855: result <= 12'b000101110101;
   30856: result <= 12'b000101110101;
   30857: result <= 12'b000101110101;
   30858: result <= 12'b000101110100;
   30859: result <= 12'b000101110100;
   30860: result <= 12'b000101110100;
   30861: result <= 12'b000101110100;
   30862: result <= 12'b000101110100;
   30863: result <= 12'b000101110011;
   30864: result <= 12'b000101110011;
   30865: result <= 12'b000101110011;
   30866: result <= 12'b000101110011;
   30867: result <= 12'b000101110011;
   30868: result <= 12'b000101110011;
   30869: result <= 12'b000101110010;
   30870: result <= 12'b000101110010;
   30871: result <= 12'b000101110010;
   30872: result <= 12'b000101110010;
   30873: result <= 12'b000101110010;
   30874: result <= 12'b000101110001;
   30875: result <= 12'b000101110001;
   30876: result <= 12'b000101110001;
   30877: result <= 12'b000101110001;
   30878: result <= 12'b000101110001;
   30879: result <= 12'b000101110000;
   30880: result <= 12'b000101110000;
   30881: result <= 12'b000101110000;
   30882: result <= 12'b000101110000;
   30883: result <= 12'b000101110000;
   30884: result <= 12'b000101101111;
   30885: result <= 12'b000101101111;
   30886: result <= 12'b000101101111;
   30887: result <= 12'b000101101111;
   30888: result <= 12'b000101101111;
   30889: result <= 12'b000101101110;
   30890: result <= 12'b000101101110;
   30891: result <= 12'b000101101110;
   30892: result <= 12'b000101101110;
   30893: result <= 12'b000101101110;
   30894: result <= 12'b000101101101;
   30895: result <= 12'b000101101101;
   30896: result <= 12'b000101101101;
   30897: result <= 12'b000101101101;
   30898: result <= 12'b000101101101;
   30899: result <= 12'b000101101101;
   30900: result <= 12'b000101101100;
   30901: result <= 12'b000101101100;
   30902: result <= 12'b000101101100;
   30903: result <= 12'b000101101100;
   30904: result <= 12'b000101101100;
   30905: result <= 12'b000101101011;
   30906: result <= 12'b000101101011;
   30907: result <= 12'b000101101011;
   30908: result <= 12'b000101101011;
   30909: result <= 12'b000101101011;
   30910: result <= 12'b000101101010;
   30911: result <= 12'b000101101010;
   30912: result <= 12'b000101101010;
   30913: result <= 12'b000101101010;
   30914: result <= 12'b000101101010;
   30915: result <= 12'b000101101001;
   30916: result <= 12'b000101101001;
   30917: result <= 12'b000101101001;
   30918: result <= 12'b000101101001;
   30919: result <= 12'b000101101001;
   30920: result <= 12'b000101101000;
   30921: result <= 12'b000101101000;
   30922: result <= 12'b000101101000;
   30923: result <= 12'b000101101000;
   30924: result <= 12'b000101101000;
   30925: result <= 12'b000101100111;
   30926: result <= 12'b000101100111;
   30927: result <= 12'b000101100111;
   30928: result <= 12'b000101100111;
   30929: result <= 12'b000101100111;
   30930: result <= 12'b000101100111;
   30931: result <= 12'b000101100110;
   30932: result <= 12'b000101100110;
   30933: result <= 12'b000101100110;
   30934: result <= 12'b000101100110;
   30935: result <= 12'b000101100110;
   30936: result <= 12'b000101100101;
   30937: result <= 12'b000101100101;
   30938: result <= 12'b000101100101;
   30939: result <= 12'b000101100101;
   30940: result <= 12'b000101100101;
   30941: result <= 12'b000101100100;
   30942: result <= 12'b000101100100;
   30943: result <= 12'b000101100100;
   30944: result <= 12'b000101100100;
   30945: result <= 12'b000101100100;
   30946: result <= 12'b000101100011;
   30947: result <= 12'b000101100011;
   30948: result <= 12'b000101100011;
   30949: result <= 12'b000101100011;
   30950: result <= 12'b000101100011;
   30951: result <= 12'b000101100010;
   30952: result <= 12'b000101100010;
   30953: result <= 12'b000101100010;
   30954: result <= 12'b000101100010;
   30955: result <= 12'b000101100010;
   30956: result <= 12'b000101100001;
   30957: result <= 12'b000101100001;
   30958: result <= 12'b000101100001;
   30959: result <= 12'b000101100001;
   30960: result <= 12'b000101100001;
   30961: result <= 12'b000101100001;
   30962: result <= 12'b000101100000;
   30963: result <= 12'b000101100000;
   30964: result <= 12'b000101100000;
   30965: result <= 12'b000101100000;
   30966: result <= 12'b000101100000;
   30967: result <= 12'b000101011111;
   30968: result <= 12'b000101011111;
   30969: result <= 12'b000101011111;
   30970: result <= 12'b000101011111;
   30971: result <= 12'b000101011111;
   30972: result <= 12'b000101011110;
   30973: result <= 12'b000101011110;
   30974: result <= 12'b000101011110;
   30975: result <= 12'b000101011110;
   30976: result <= 12'b000101011110;
   30977: result <= 12'b000101011101;
   30978: result <= 12'b000101011101;
   30979: result <= 12'b000101011101;
   30980: result <= 12'b000101011101;
   30981: result <= 12'b000101011101;
   30982: result <= 12'b000101011100;
   30983: result <= 12'b000101011100;
   30984: result <= 12'b000101011100;
   30985: result <= 12'b000101011100;
   30986: result <= 12'b000101011100;
   30987: result <= 12'b000101011100;
   30988: result <= 12'b000101011011;
   30989: result <= 12'b000101011011;
   30990: result <= 12'b000101011011;
   30991: result <= 12'b000101011011;
   30992: result <= 12'b000101011011;
   30993: result <= 12'b000101011010;
   30994: result <= 12'b000101011010;
   30995: result <= 12'b000101011010;
   30996: result <= 12'b000101011010;
   30997: result <= 12'b000101011010;
   30998: result <= 12'b000101011001;
   30999: result <= 12'b000101011001;
   31000: result <= 12'b000101011001;
   31001: result <= 12'b000101011001;
   31002: result <= 12'b000101011001;
   31003: result <= 12'b000101011000;
   31004: result <= 12'b000101011000;
   31005: result <= 12'b000101011000;
   31006: result <= 12'b000101011000;
   31007: result <= 12'b000101011000;
   31008: result <= 12'b000101010111;
   31009: result <= 12'b000101010111;
   31010: result <= 12'b000101010111;
   31011: result <= 12'b000101010111;
   31012: result <= 12'b000101010111;
   31013: result <= 12'b000101010110;
   31014: result <= 12'b000101010110;
   31015: result <= 12'b000101010110;
   31016: result <= 12'b000101010110;
   31017: result <= 12'b000101010110;
   31018: result <= 12'b000101010110;
   31019: result <= 12'b000101010101;
   31020: result <= 12'b000101010101;
   31021: result <= 12'b000101010101;
   31022: result <= 12'b000101010101;
   31023: result <= 12'b000101010101;
   31024: result <= 12'b000101010100;
   31025: result <= 12'b000101010100;
   31026: result <= 12'b000101010100;
   31027: result <= 12'b000101010100;
   31028: result <= 12'b000101010100;
   31029: result <= 12'b000101010011;
   31030: result <= 12'b000101010011;
   31031: result <= 12'b000101010011;
   31032: result <= 12'b000101010011;
   31033: result <= 12'b000101010011;
   31034: result <= 12'b000101010010;
   31035: result <= 12'b000101010010;
   31036: result <= 12'b000101010010;
   31037: result <= 12'b000101010010;
   31038: result <= 12'b000101010010;
   31039: result <= 12'b000101010001;
   31040: result <= 12'b000101010001;
   31041: result <= 12'b000101010001;
   31042: result <= 12'b000101010001;
   31043: result <= 12'b000101010001;
   31044: result <= 12'b000101010000;
   31045: result <= 12'b000101010000;
   31046: result <= 12'b000101010000;
   31047: result <= 12'b000101010000;
   31048: result <= 12'b000101010000;
   31049: result <= 12'b000101001111;
   31050: result <= 12'b000101001111;
   31051: result <= 12'b000101001111;
   31052: result <= 12'b000101001111;
   31053: result <= 12'b000101001111;
   31054: result <= 12'b000101001111;
   31055: result <= 12'b000101001110;
   31056: result <= 12'b000101001110;
   31057: result <= 12'b000101001110;
   31058: result <= 12'b000101001110;
   31059: result <= 12'b000101001110;
   31060: result <= 12'b000101001101;
   31061: result <= 12'b000101001101;
   31062: result <= 12'b000101001101;
   31063: result <= 12'b000101001101;
   31064: result <= 12'b000101001101;
   31065: result <= 12'b000101001100;
   31066: result <= 12'b000101001100;
   31067: result <= 12'b000101001100;
   31068: result <= 12'b000101001100;
   31069: result <= 12'b000101001100;
   31070: result <= 12'b000101001011;
   31071: result <= 12'b000101001011;
   31072: result <= 12'b000101001011;
   31073: result <= 12'b000101001011;
   31074: result <= 12'b000101001011;
   31075: result <= 12'b000101001010;
   31076: result <= 12'b000101001010;
   31077: result <= 12'b000101001010;
   31078: result <= 12'b000101001010;
   31079: result <= 12'b000101001010;
   31080: result <= 12'b000101001001;
   31081: result <= 12'b000101001001;
   31082: result <= 12'b000101001001;
   31083: result <= 12'b000101001001;
   31084: result <= 12'b000101001001;
   31085: result <= 12'b000101001001;
   31086: result <= 12'b000101001000;
   31087: result <= 12'b000101001000;
   31088: result <= 12'b000101001000;
   31089: result <= 12'b000101001000;
   31090: result <= 12'b000101001000;
   31091: result <= 12'b000101000111;
   31092: result <= 12'b000101000111;
   31093: result <= 12'b000101000111;
   31094: result <= 12'b000101000111;
   31095: result <= 12'b000101000111;
   31096: result <= 12'b000101000110;
   31097: result <= 12'b000101000110;
   31098: result <= 12'b000101000110;
   31099: result <= 12'b000101000110;
   31100: result <= 12'b000101000110;
   31101: result <= 12'b000101000101;
   31102: result <= 12'b000101000101;
   31103: result <= 12'b000101000101;
   31104: result <= 12'b000101000101;
   31105: result <= 12'b000101000101;
   31106: result <= 12'b000101000100;
   31107: result <= 12'b000101000100;
   31108: result <= 12'b000101000100;
   31109: result <= 12'b000101000100;
   31110: result <= 12'b000101000100;
   31111: result <= 12'b000101000011;
   31112: result <= 12'b000101000011;
   31113: result <= 12'b000101000011;
   31114: result <= 12'b000101000011;
   31115: result <= 12'b000101000011;
   31116: result <= 12'b000101000011;
   31117: result <= 12'b000101000010;
   31118: result <= 12'b000101000010;
   31119: result <= 12'b000101000010;
   31120: result <= 12'b000101000010;
   31121: result <= 12'b000101000010;
   31122: result <= 12'b000101000001;
   31123: result <= 12'b000101000001;
   31124: result <= 12'b000101000001;
   31125: result <= 12'b000101000001;
   31126: result <= 12'b000101000001;
   31127: result <= 12'b000101000000;
   31128: result <= 12'b000101000000;
   31129: result <= 12'b000101000000;
   31130: result <= 12'b000101000000;
   31131: result <= 12'b000101000000;
   31132: result <= 12'b000100111111;
   31133: result <= 12'b000100111111;
   31134: result <= 12'b000100111111;
   31135: result <= 12'b000100111111;
   31136: result <= 12'b000100111111;
   31137: result <= 12'b000100111110;
   31138: result <= 12'b000100111110;
   31139: result <= 12'b000100111110;
   31140: result <= 12'b000100111110;
   31141: result <= 12'b000100111110;
   31142: result <= 12'b000100111101;
   31143: result <= 12'b000100111101;
   31144: result <= 12'b000100111101;
   31145: result <= 12'b000100111101;
   31146: result <= 12'b000100111101;
   31147: result <= 12'b000100111101;
   31148: result <= 12'b000100111100;
   31149: result <= 12'b000100111100;
   31150: result <= 12'b000100111100;
   31151: result <= 12'b000100111100;
   31152: result <= 12'b000100111100;
   31153: result <= 12'b000100111011;
   31154: result <= 12'b000100111011;
   31155: result <= 12'b000100111011;
   31156: result <= 12'b000100111011;
   31157: result <= 12'b000100111011;
   31158: result <= 12'b000100111010;
   31159: result <= 12'b000100111010;
   31160: result <= 12'b000100111010;
   31161: result <= 12'b000100111010;
   31162: result <= 12'b000100111010;
   31163: result <= 12'b000100111001;
   31164: result <= 12'b000100111001;
   31165: result <= 12'b000100111001;
   31166: result <= 12'b000100111001;
   31167: result <= 12'b000100111001;
   31168: result <= 12'b000100111000;
   31169: result <= 12'b000100111000;
   31170: result <= 12'b000100111000;
   31171: result <= 12'b000100111000;
   31172: result <= 12'b000100111000;
   31173: result <= 12'b000100110111;
   31174: result <= 12'b000100110111;
   31175: result <= 12'b000100110111;
   31176: result <= 12'b000100110111;
   31177: result <= 12'b000100110111;
   31178: result <= 12'b000100110110;
   31179: result <= 12'b000100110110;
   31180: result <= 12'b000100110110;
   31181: result <= 12'b000100110110;
   31182: result <= 12'b000100110110;
   31183: result <= 12'b000100110110;
   31184: result <= 12'b000100110101;
   31185: result <= 12'b000100110101;
   31186: result <= 12'b000100110101;
   31187: result <= 12'b000100110101;
   31188: result <= 12'b000100110101;
   31189: result <= 12'b000100110100;
   31190: result <= 12'b000100110100;
   31191: result <= 12'b000100110100;
   31192: result <= 12'b000100110100;
   31193: result <= 12'b000100110100;
   31194: result <= 12'b000100110011;
   31195: result <= 12'b000100110011;
   31196: result <= 12'b000100110011;
   31197: result <= 12'b000100110011;
   31198: result <= 12'b000100110011;
   31199: result <= 12'b000100110010;
   31200: result <= 12'b000100110010;
   31201: result <= 12'b000100110010;
   31202: result <= 12'b000100110010;
   31203: result <= 12'b000100110010;
   31204: result <= 12'b000100110001;
   31205: result <= 12'b000100110001;
   31206: result <= 12'b000100110001;
   31207: result <= 12'b000100110001;
   31208: result <= 12'b000100110001;
   31209: result <= 12'b000100110000;
   31210: result <= 12'b000100110000;
   31211: result <= 12'b000100110000;
   31212: result <= 12'b000100110000;
   31213: result <= 12'b000100110000;
   31214: result <= 12'b000100101111;
   31215: result <= 12'b000100101111;
   31216: result <= 12'b000100101111;
   31217: result <= 12'b000100101111;
   31218: result <= 12'b000100101111;
   31219: result <= 12'b000100101111;
   31220: result <= 12'b000100101110;
   31221: result <= 12'b000100101110;
   31222: result <= 12'b000100101110;
   31223: result <= 12'b000100101110;
   31224: result <= 12'b000100101110;
   31225: result <= 12'b000100101101;
   31226: result <= 12'b000100101101;
   31227: result <= 12'b000100101101;
   31228: result <= 12'b000100101101;
   31229: result <= 12'b000100101101;
   31230: result <= 12'b000100101100;
   31231: result <= 12'b000100101100;
   31232: result <= 12'b000100101100;
   31233: result <= 12'b000100101100;
   31234: result <= 12'b000100101100;
   31235: result <= 12'b000100101011;
   31236: result <= 12'b000100101011;
   31237: result <= 12'b000100101011;
   31238: result <= 12'b000100101011;
   31239: result <= 12'b000100101011;
   31240: result <= 12'b000100101010;
   31241: result <= 12'b000100101010;
   31242: result <= 12'b000100101010;
   31243: result <= 12'b000100101010;
   31244: result <= 12'b000100101010;
   31245: result <= 12'b000100101001;
   31246: result <= 12'b000100101001;
   31247: result <= 12'b000100101001;
   31248: result <= 12'b000100101001;
   31249: result <= 12'b000100101001;
   31250: result <= 12'b000100101001;
   31251: result <= 12'b000100101000;
   31252: result <= 12'b000100101000;
   31253: result <= 12'b000100101000;
   31254: result <= 12'b000100101000;
   31255: result <= 12'b000100101000;
   31256: result <= 12'b000100100111;
   31257: result <= 12'b000100100111;
   31258: result <= 12'b000100100111;
   31259: result <= 12'b000100100111;
   31260: result <= 12'b000100100111;
   31261: result <= 12'b000100100110;
   31262: result <= 12'b000100100110;
   31263: result <= 12'b000100100110;
   31264: result <= 12'b000100100110;
   31265: result <= 12'b000100100110;
   31266: result <= 12'b000100100101;
   31267: result <= 12'b000100100101;
   31268: result <= 12'b000100100101;
   31269: result <= 12'b000100100101;
   31270: result <= 12'b000100100101;
   31271: result <= 12'b000100100100;
   31272: result <= 12'b000100100100;
   31273: result <= 12'b000100100100;
   31274: result <= 12'b000100100100;
   31275: result <= 12'b000100100100;
   31276: result <= 12'b000100100011;
   31277: result <= 12'b000100100011;
   31278: result <= 12'b000100100011;
   31279: result <= 12'b000100100011;
   31280: result <= 12'b000100100011;
   31281: result <= 12'b000100100010;
   31282: result <= 12'b000100100010;
   31283: result <= 12'b000100100010;
   31284: result <= 12'b000100100010;
   31285: result <= 12'b000100100010;
   31286: result <= 12'b000100100010;
   31287: result <= 12'b000100100001;
   31288: result <= 12'b000100100001;
   31289: result <= 12'b000100100001;
   31290: result <= 12'b000100100001;
   31291: result <= 12'b000100100001;
   31292: result <= 12'b000100100000;
   31293: result <= 12'b000100100000;
   31294: result <= 12'b000100100000;
   31295: result <= 12'b000100100000;
   31296: result <= 12'b000100100000;
   31297: result <= 12'b000100011111;
   31298: result <= 12'b000100011111;
   31299: result <= 12'b000100011111;
   31300: result <= 12'b000100011111;
   31301: result <= 12'b000100011111;
   31302: result <= 12'b000100011110;
   31303: result <= 12'b000100011110;
   31304: result <= 12'b000100011110;
   31305: result <= 12'b000100011110;
   31306: result <= 12'b000100011110;
   31307: result <= 12'b000100011101;
   31308: result <= 12'b000100011101;
   31309: result <= 12'b000100011101;
   31310: result <= 12'b000100011101;
   31311: result <= 12'b000100011101;
   31312: result <= 12'b000100011100;
   31313: result <= 12'b000100011100;
   31314: result <= 12'b000100011100;
   31315: result <= 12'b000100011100;
   31316: result <= 12'b000100011100;
   31317: result <= 12'b000100011011;
   31318: result <= 12'b000100011011;
   31319: result <= 12'b000100011011;
   31320: result <= 12'b000100011011;
   31321: result <= 12'b000100011011;
   31322: result <= 12'b000100011011;
   31323: result <= 12'b000100011010;
   31324: result <= 12'b000100011010;
   31325: result <= 12'b000100011010;
   31326: result <= 12'b000100011010;
   31327: result <= 12'b000100011010;
   31328: result <= 12'b000100011001;
   31329: result <= 12'b000100011001;
   31330: result <= 12'b000100011001;
   31331: result <= 12'b000100011001;
   31332: result <= 12'b000100011001;
   31333: result <= 12'b000100011000;
   31334: result <= 12'b000100011000;
   31335: result <= 12'b000100011000;
   31336: result <= 12'b000100011000;
   31337: result <= 12'b000100011000;
   31338: result <= 12'b000100010111;
   31339: result <= 12'b000100010111;
   31340: result <= 12'b000100010111;
   31341: result <= 12'b000100010111;
   31342: result <= 12'b000100010111;
   31343: result <= 12'b000100010110;
   31344: result <= 12'b000100010110;
   31345: result <= 12'b000100010110;
   31346: result <= 12'b000100010110;
   31347: result <= 12'b000100010110;
   31348: result <= 12'b000100010101;
   31349: result <= 12'b000100010101;
   31350: result <= 12'b000100010101;
   31351: result <= 12'b000100010101;
   31352: result <= 12'b000100010101;
   31353: result <= 12'b000100010100;
   31354: result <= 12'b000100010100;
   31355: result <= 12'b000100010100;
   31356: result <= 12'b000100010100;
   31357: result <= 12'b000100010100;
   31358: result <= 12'b000100010100;
   31359: result <= 12'b000100010011;
   31360: result <= 12'b000100010011;
   31361: result <= 12'b000100010011;
   31362: result <= 12'b000100010011;
   31363: result <= 12'b000100010011;
   31364: result <= 12'b000100010010;
   31365: result <= 12'b000100010010;
   31366: result <= 12'b000100010010;
   31367: result <= 12'b000100010010;
   31368: result <= 12'b000100010010;
   31369: result <= 12'b000100010001;
   31370: result <= 12'b000100010001;
   31371: result <= 12'b000100010001;
   31372: result <= 12'b000100010001;
   31373: result <= 12'b000100010001;
   31374: result <= 12'b000100010000;
   31375: result <= 12'b000100010000;
   31376: result <= 12'b000100010000;
   31377: result <= 12'b000100010000;
   31378: result <= 12'b000100010000;
   31379: result <= 12'b000100001111;
   31380: result <= 12'b000100001111;
   31381: result <= 12'b000100001111;
   31382: result <= 12'b000100001111;
   31383: result <= 12'b000100001111;
   31384: result <= 12'b000100001110;
   31385: result <= 12'b000100001110;
   31386: result <= 12'b000100001110;
   31387: result <= 12'b000100001110;
   31388: result <= 12'b000100001110;
   31389: result <= 12'b000100001101;
   31390: result <= 12'b000100001101;
   31391: result <= 12'b000100001101;
   31392: result <= 12'b000100001101;
   31393: result <= 12'b000100001101;
   31394: result <= 12'b000100001101;
   31395: result <= 12'b000100001100;
   31396: result <= 12'b000100001100;
   31397: result <= 12'b000100001100;
   31398: result <= 12'b000100001100;
   31399: result <= 12'b000100001100;
   31400: result <= 12'b000100001011;
   31401: result <= 12'b000100001011;
   31402: result <= 12'b000100001011;
   31403: result <= 12'b000100001011;
   31404: result <= 12'b000100001011;
   31405: result <= 12'b000100001010;
   31406: result <= 12'b000100001010;
   31407: result <= 12'b000100001010;
   31408: result <= 12'b000100001010;
   31409: result <= 12'b000100001010;
   31410: result <= 12'b000100001001;
   31411: result <= 12'b000100001001;
   31412: result <= 12'b000100001001;
   31413: result <= 12'b000100001001;
   31414: result <= 12'b000100001001;
   31415: result <= 12'b000100001000;
   31416: result <= 12'b000100001000;
   31417: result <= 12'b000100001000;
   31418: result <= 12'b000100001000;
   31419: result <= 12'b000100001000;
   31420: result <= 12'b000100000111;
   31421: result <= 12'b000100000111;
   31422: result <= 12'b000100000111;
   31423: result <= 12'b000100000111;
   31424: result <= 12'b000100000111;
   31425: result <= 12'b000100000110;
   31426: result <= 12'b000100000110;
   31427: result <= 12'b000100000110;
   31428: result <= 12'b000100000110;
   31429: result <= 12'b000100000110;
   31430: result <= 12'b000100000101;
   31431: result <= 12'b000100000101;
   31432: result <= 12'b000100000101;
   31433: result <= 12'b000100000101;
   31434: result <= 12'b000100000101;
   31435: result <= 12'b000100000101;
   31436: result <= 12'b000100000100;
   31437: result <= 12'b000100000100;
   31438: result <= 12'b000100000100;
   31439: result <= 12'b000100000100;
   31440: result <= 12'b000100000100;
   31441: result <= 12'b000100000011;
   31442: result <= 12'b000100000011;
   31443: result <= 12'b000100000011;
   31444: result <= 12'b000100000011;
   31445: result <= 12'b000100000011;
   31446: result <= 12'b000100000010;
   31447: result <= 12'b000100000010;
   31448: result <= 12'b000100000010;
   31449: result <= 12'b000100000010;
   31450: result <= 12'b000100000010;
   31451: result <= 12'b000100000001;
   31452: result <= 12'b000100000001;
   31453: result <= 12'b000100000001;
   31454: result <= 12'b000100000001;
   31455: result <= 12'b000100000001;
   31456: result <= 12'b000100000000;
   31457: result <= 12'b000100000000;
   31458: result <= 12'b000100000000;
   31459: result <= 12'b000100000000;
   31460: result <= 12'b000100000000;
   31461: result <= 12'b000011111111;
   31462: result <= 12'b000011111111;
   31463: result <= 12'b000011111111;
   31464: result <= 12'b000011111111;
   31465: result <= 12'b000011111111;
   31466: result <= 12'b000011111110;
   31467: result <= 12'b000011111110;
   31468: result <= 12'b000011111110;
   31469: result <= 12'b000011111110;
   31470: result <= 12'b000011111110;
   31471: result <= 12'b000011111110;
   31472: result <= 12'b000011111101;
   31473: result <= 12'b000011111101;
   31474: result <= 12'b000011111101;
   31475: result <= 12'b000011111101;
   31476: result <= 12'b000011111101;
   31477: result <= 12'b000011111100;
   31478: result <= 12'b000011111100;
   31479: result <= 12'b000011111100;
   31480: result <= 12'b000011111100;
   31481: result <= 12'b000011111100;
   31482: result <= 12'b000011111011;
   31483: result <= 12'b000011111011;
   31484: result <= 12'b000011111011;
   31485: result <= 12'b000011111011;
   31486: result <= 12'b000011111011;
   31487: result <= 12'b000011111010;
   31488: result <= 12'b000011111010;
   31489: result <= 12'b000011111010;
   31490: result <= 12'b000011111010;
   31491: result <= 12'b000011111010;
   31492: result <= 12'b000011111001;
   31493: result <= 12'b000011111001;
   31494: result <= 12'b000011111001;
   31495: result <= 12'b000011111001;
   31496: result <= 12'b000011111001;
   31497: result <= 12'b000011111000;
   31498: result <= 12'b000011111000;
   31499: result <= 12'b000011111000;
   31500: result <= 12'b000011111000;
   31501: result <= 12'b000011111000;
   31502: result <= 12'b000011110111;
   31503: result <= 12'b000011110111;
   31504: result <= 12'b000011110111;
   31505: result <= 12'b000011110111;
   31506: result <= 12'b000011110111;
   31507: result <= 12'b000011110110;
   31508: result <= 12'b000011110110;
   31509: result <= 12'b000011110110;
   31510: result <= 12'b000011110110;
   31511: result <= 12'b000011110110;
   31512: result <= 12'b000011110110;
   31513: result <= 12'b000011110101;
   31514: result <= 12'b000011110101;
   31515: result <= 12'b000011110101;
   31516: result <= 12'b000011110101;
   31517: result <= 12'b000011110101;
   31518: result <= 12'b000011110100;
   31519: result <= 12'b000011110100;
   31520: result <= 12'b000011110100;
   31521: result <= 12'b000011110100;
   31522: result <= 12'b000011110100;
   31523: result <= 12'b000011110011;
   31524: result <= 12'b000011110011;
   31525: result <= 12'b000011110011;
   31526: result <= 12'b000011110011;
   31527: result <= 12'b000011110011;
   31528: result <= 12'b000011110010;
   31529: result <= 12'b000011110010;
   31530: result <= 12'b000011110010;
   31531: result <= 12'b000011110010;
   31532: result <= 12'b000011110010;
   31533: result <= 12'b000011110001;
   31534: result <= 12'b000011110001;
   31535: result <= 12'b000011110001;
   31536: result <= 12'b000011110001;
   31537: result <= 12'b000011110001;
   31538: result <= 12'b000011110000;
   31539: result <= 12'b000011110000;
   31540: result <= 12'b000011110000;
   31541: result <= 12'b000011110000;
   31542: result <= 12'b000011110000;
   31543: result <= 12'b000011101111;
   31544: result <= 12'b000011101111;
   31545: result <= 12'b000011101111;
   31546: result <= 12'b000011101111;
   31547: result <= 12'b000011101111;
   31548: result <= 12'b000011101111;
   31549: result <= 12'b000011101110;
   31550: result <= 12'b000011101110;
   31551: result <= 12'b000011101110;
   31552: result <= 12'b000011101110;
   31553: result <= 12'b000011101110;
   31554: result <= 12'b000011101101;
   31555: result <= 12'b000011101101;
   31556: result <= 12'b000011101101;
   31557: result <= 12'b000011101101;
   31558: result <= 12'b000011101101;
   31559: result <= 12'b000011101100;
   31560: result <= 12'b000011101100;
   31561: result <= 12'b000011101100;
   31562: result <= 12'b000011101100;
   31563: result <= 12'b000011101100;
   31564: result <= 12'b000011101011;
   31565: result <= 12'b000011101011;
   31566: result <= 12'b000011101011;
   31567: result <= 12'b000011101011;
   31568: result <= 12'b000011101011;
   31569: result <= 12'b000011101010;
   31570: result <= 12'b000011101010;
   31571: result <= 12'b000011101010;
   31572: result <= 12'b000011101010;
   31573: result <= 12'b000011101010;
   31574: result <= 12'b000011101001;
   31575: result <= 12'b000011101001;
   31576: result <= 12'b000011101001;
   31577: result <= 12'b000011101001;
   31578: result <= 12'b000011101001;
   31579: result <= 12'b000011101000;
   31580: result <= 12'b000011101000;
   31581: result <= 12'b000011101000;
   31582: result <= 12'b000011101000;
   31583: result <= 12'b000011101000;
   31584: result <= 12'b000011100111;
   31585: result <= 12'b000011100111;
   31586: result <= 12'b000011100111;
   31587: result <= 12'b000011100111;
   31588: result <= 12'b000011100111;
   31589: result <= 12'b000011100111;
   31590: result <= 12'b000011100110;
   31591: result <= 12'b000011100110;
   31592: result <= 12'b000011100110;
   31593: result <= 12'b000011100110;
   31594: result <= 12'b000011100110;
   31595: result <= 12'b000011100101;
   31596: result <= 12'b000011100101;
   31597: result <= 12'b000011100101;
   31598: result <= 12'b000011100101;
   31599: result <= 12'b000011100101;
   31600: result <= 12'b000011100100;
   31601: result <= 12'b000011100100;
   31602: result <= 12'b000011100100;
   31603: result <= 12'b000011100100;
   31604: result <= 12'b000011100100;
   31605: result <= 12'b000011100011;
   31606: result <= 12'b000011100011;
   31607: result <= 12'b000011100011;
   31608: result <= 12'b000011100011;
   31609: result <= 12'b000011100011;
   31610: result <= 12'b000011100010;
   31611: result <= 12'b000011100010;
   31612: result <= 12'b000011100010;
   31613: result <= 12'b000011100010;
   31614: result <= 12'b000011100010;
   31615: result <= 12'b000011100001;
   31616: result <= 12'b000011100001;
   31617: result <= 12'b000011100001;
   31618: result <= 12'b000011100001;
   31619: result <= 12'b000011100001;
   31620: result <= 12'b000011100000;
   31621: result <= 12'b000011100000;
   31622: result <= 12'b000011100000;
   31623: result <= 12'b000011100000;
   31624: result <= 12'b000011100000;
   31625: result <= 12'b000011011111;
   31626: result <= 12'b000011011111;
   31627: result <= 12'b000011011111;
   31628: result <= 12'b000011011111;
   31629: result <= 12'b000011011111;
   31630: result <= 12'b000011011111;
   31631: result <= 12'b000011011110;
   31632: result <= 12'b000011011110;
   31633: result <= 12'b000011011110;
   31634: result <= 12'b000011011110;
   31635: result <= 12'b000011011110;
   31636: result <= 12'b000011011101;
   31637: result <= 12'b000011011101;
   31638: result <= 12'b000011011101;
   31639: result <= 12'b000011011101;
   31640: result <= 12'b000011011101;
   31641: result <= 12'b000011011100;
   31642: result <= 12'b000011011100;
   31643: result <= 12'b000011011100;
   31644: result <= 12'b000011011100;
   31645: result <= 12'b000011011100;
   31646: result <= 12'b000011011011;
   31647: result <= 12'b000011011011;
   31648: result <= 12'b000011011011;
   31649: result <= 12'b000011011011;
   31650: result <= 12'b000011011011;
   31651: result <= 12'b000011011010;
   31652: result <= 12'b000011011010;
   31653: result <= 12'b000011011010;
   31654: result <= 12'b000011011010;
   31655: result <= 12'b000011011010;
   31656: result <= 12'b000011011001;
   31657: result <= 12'b000011011001;
   31658: result <= 12'b000011011001;
   31659: result <= 12'b000011011001;
   31660: result <= 12'b000011011001;
   31661: result <= 12'b000011011000;
   31662: result <= 12'b000011011000;
   31663: result <= 12'b000011011000;
   31664: result <= 12'b000011011000;
   31665: result <= 12'b000011011000;
   31666: result <= 12'b000011010111;
   31667: result <= 12'b000011010111;
   31668: result <= 12'b000011010111;
   31669: result <= 12'b000011010111;
   31670: result <= 12'b000011010111;
   31671: result <= 12'b000011010110;
   31672: result <= 12'b000011010110;
   31673: result <= 12'b000011010110;
   31674: result <= 12'b000011010110;
   31675: result <= 12'b000011010110;
   31676: result <= 12'b000011010110;
   31677: result <= 12'b000011010101;
   31678: result <= 12'b000011010101;
   31679: result <= 12'b000011010101;
   31680: result <= 12'b000011010101;
   31681: result <= 12'b000011010101;
   31682: result <= 12'b000011010100;
   31683: result <= 12'b000011010100;
   31684: result <= 12'b000011010100;
   31685: result <= 12'b000011010100;
   31686: result <= 12'b000011010100;
   31687: result <= 12'b000011010011;
   31688: result <= 12'b000011010011;
   31689: result <= 12'b000011010011;
   31690: result <= 12'b000011010011;
   31691: result <= 12'b000011010011;
   31692: result <= 12'b000011010010;
   31693: result <= 12'b000011010010;
   31694: result <= 12'b000011010010;
   31695: result <= 12'b000011010010;
   31696: result <= 12'b000011010010;
   31697: result <= 12'b000011010001;
   31698: result <= 12'b000011010001;
   31699: result <= 12'b000011010001;
   31700: result <= 12'b000011010001;
   31701: result <= 12'b000011010001;
   31702: result <= 12'b000011010000;
   31703: result <= 12'b000011010000;
   31704: result <= 12'b000011010000;
   31705: result <= 12'b000011010000;
   31706: result <= 12'b000011010000;
   31707: result <= 12'b000011001111;
   31708: result <= 12'b000011001111;
   31709: result <= 12'b000011001111;
   31710: result <= 12'b000011001111;
   31711: result <= 12'b000011001111;
   31712: result <= 12'b000011001110;
   31713: result <= 12'b000011001110;
   31714: result <= 12'b000011001110;
   31715: result <= 12'b000011001110;
   31716: result <= 12'b000011001110;
   31717: result <= 12'b000011001110;
   31718: result <= 12'b000011001101;
   31719: result <= 12'b000011001101;
   31720: result <= 12'b000011001101;
   31721: result <= 12'b000011001101;
   31722: result <= 12'b000011001101;
   31723: result <= 12'b000011001100;
   31724: result <= 12'b000011001100;
   31725: result <= 12'b000011001100;
   31726: result <= 12'b000011001100;
   31727: result <= 12'b000011001100;
   31728: result <= 12'b000011001011;
   31729: result <= 12'b000011001011;
   31730: result <= 12'b000011001011;
   31731: result <= 12'b000011001011;
   31732: result <= 12'b000011001011;
   31733: result <= 12'b000011001010;
   31734: result <= 12'b000011001010;
   31735: result <= 12'b000011001010;
   31736: result <= 12'b000011001010;
   31737: result <= 12'b000011001010;
   31738: result <= 12'b000011001001;
   31739: result <= 12'b000011001001;
   31740: result <= 12'b000011001001;
   31741: result <= 12'b000011001001;
   31742: result <= 12'b000011001001;
   31743: result <= 12'b000011001000;
   31744: result <= 12'b000011001000;
   31745: result <= 12'b000011001000;
   31746: result <= 12'b000011001000;
   31747: result <= 12'b000011001000;
   31748: result <= 12'b000011000111;
   31749: result <= 12'b000011000111;
   31750: result <= 12'b000011000111;
   31751: result <= 12'b000011000111;
   31752: result <= 12'b000011000111;
   31753: result <= 12'b000011000110;
   31754: result <= 12'b000011000110;
   31755: result <= 12'b000011000110;
   31756: result <= 12'b000011000110;
   31757: result <= 12'b000011000110;
   31758: result <= 12'b000011000110;
   31759: result <= 12'b000011000101;
   31760: result <= 12'b000011000101;
   31761: result <= 12'b000011000101;
   31762: result <= 12'b000011000101;
   31763: result <= 12'b000011000101;
   31764: result <= 12'b000011000100;
   31765: result <= 12'b000011000100;
   31766: result <= 12'b000011000100;
   31767: result <= 12'b000011000100;
   31768: result <= 12'b000011000100;
   31769: result <= 12'b000011000011;
   31770: result <= 12'b000011000011;
   31771: result <= 12'b000011000011;
   31772: result <= 12'b000011000011;
   31773: result <= 12'b000011000011;
   31774: result <= 12'b000011000010;
   31775: result <= 12'b000011000010;
   31776: result <= 12'b000011000010;
   31777: result <= 12'b000011000010;
   31778: result <= 12'b000011000010;
   31779: result <= 12'b000011000001;
   31780: result <= 12'b000011000001;
   31781: result <= 12'b000011000001;
   31782: result <= 12'b000011000001;
   31783: result <= 12'b000011000001;
   31784: result <= 12'b000011000000;
   31785: result <= 12'b000011000000;
   31786: result <= 12'b000011000000;
   31787: result <= 12'b000011000000;
   31788: result <= 12'b000011000000;
   31789: result <= 12'b000010111111;
   31790: result <= 12'b000010111111;
   31791: result <= 12'b000010111111;
   31792: result <= 12'b000010111111;
   31793: result <= 12'b000010111111;
   31794: result <= 12'b000010111110;
   31795: result <= 12'b000010111110;
   31796: result <= 12'b000010111110;
   31797: result <= 12'b000010111110;
   31798: result <= 12'b000010111110;
   31799: result <= 12'b000010111101;
   31800: result <= 12'b000010111101;
   31801: result <= 12'b000010111101;
   31802: result <= 12'b000010111101;
   31803: result <= 12'b000010111101;
   31804: result <= 12'b000010111101;
   31805: result <= 12'b000010111100;
   31806: result <= 12'b000010111100;
   31807: result <= 12'b000010111100;
   31808: result <= 12'b000010111100;
   31809: result <= 12'b000010111100;
   31810: result <= 12'b000010111011;
   31811: result <= 12'b000010111011;
   31812: result <= 12'b000010111011;
   31813: result <= 12'b000010111011;
   31814: result <= 12'b000010111011;
   31815: result <= 12'b000010111010;
   31816: result <= 12'b000010111010;
   31817: result <= 12'b000010111010;
   31818: result <= 12'b000010111010;
   31819: result <= 12'b000010111010;
   31820: result <= 12'b000010111001;
   31821: result <= 12'b000010111001;
   31822: result <= 12'b000010111001;
   31823: result <= 12'b000010111001;
   31824: result <= 12'b000010111001;
   31825: result <= 12'b000010111000;
   31826: result <= 12'b000010111000;
   31827: result <= 12'b000010111000;
   31828: result <= 12'b000010111000;
   31829: result <= 12'b000010111000;
   31830: result <= 12'b000010110111;
   31831: result <= 12'b000010110111;
   31832: result <= 12'b000010110111;
   31833: result <= 12'b000010110111;
   31834: result <= 12'b000010110111;
   31835: result <= 12'b000010110110;
   31836: result <= 12'b000010110110;
   31837: result <= 12'b000010110110;
   31838: result <= 12'b000010110110;
   31839: result <= 12'b000010110110;
   31840: result <= 12'b000010110101;
   31841: result <= 12'b000010110101;
   31842: result <= 12'b000010110101;
   31843: result <= 12'b000010110101;
   31844: result <= 12'b000010110101;
   31845: result <= 12'b000010110100;
   31846: result <= 12'b000010110100;
   31847: result <= 12'b000010110100;
   31848: result <= 12'b000010110100;
   31849: result <= 12'b000010110100;
   31850: result <= 12'b000010110100;
   31851: result <= 12'b000010110011;
   31852: result <= 12'b000010110011;
   31853: result <= 12'b000010110011;
   31854: result <= 12'b000010110011;
   31855: result <= 12'b000010110011;
   31856: result <= 12'b000010110010;
   31857: result <= 12'b000010110010;
   31858: result <= 12'b000010110010;
   31859: result <= 12'b000010110010;
   31860: result <= 12'b000010110010;
   31861: result <= 12'b000010110001;
   31862: result <= 12'b000010110001;
   31863: result <= 12'b000010110001;
   31864: result <= 12'b000010110001;
   31865: result <= 12'b000010110001;
   31866: result <= 12'b000010110000;
   31867: result <= 12'b000010110000;
   31868: result <= 12'b000010110000;
   31869: result <= 12'b000010110000;
   31870: result <= 12'b000010110000;
   31871: result <= 12'b000010101111;
   31872: result <= 12'b000010101111;
   31873: result <= 12'b000010101111;
   31874: result <= 12'b000010101111;
   31875: result <= 12'b000010101111;
   31876: result <= 12'b000010101110;
   31877: result <= 12'b000010101110;
   31878: result <= 12'b000010101110;
   31879: result <= 12'b000010101110;
   31880: result <= 12'b000010101110;
   31881: result <= 12'b000010101101;
   31882: result <= 12'b000010101101;
   31883: result <= 12'b000010101101;
   31884: result <= 12'b000010101101;
   31885: result <= 12'b000010101101;
   31886: result <= 12'b000010101100;
   31887: result <= 12'b000010101100;
   31888: result <= 12'b000010101100;
   31889: result <= 12'b000010101100;
   31890: result <= 12'b000010101100;
   31891: result <= 12'b000010101011;
   31892: result <= 12'b000010101011;
   31893: result <= 12'b000010101011;
   31894: result <= 12'b000010101011;
   31895: result <= 12'b000010101011;
   31896: result <= 12'b000010101011;
   31897: result <= 12'b000010101010;
   31898: result <= 12'b000010101010;
   31899: result <= 12'b000010101010;
   31900: result <= 12'b000010101010;
   31901: result <= 12'b000010101010;
   31902: result <= 12'b000010101001;
   31903: result <= 12'b000010101001;
   31904: result <= 12'b000010101001;
   31905: result <= 12'b000010101001;
   31906: result <= 12'b000010101001;
   31907: result <= 12'b000010101000;
   31908: result <= 12'b000010101000;
   31909: result <= 12'b000010101000;
   31910: result <= 12'b000010101000;
   31911: result <= 12'b000010101000;
   31912: result <= 12'b000010100111;
   31913: result <= 12'b000010100111;
   31914: result <= 12'b000010100111;
   31915: result <= 12'b000010100111;
   31916: result <= 12'b000010100111;
   31917: result <= 12'b000010100110;
   31918: result <= 12'b000010100110;
   31919: result <= 12'b000010100110;
   31920: result <= 12'b000010100110;
   31921: result <= 12'b000010100110;
   31922: result <= 12'b000010100101;
   31923: result <= 12'b000010100101;
   31924: result <= 12'b000010100101;
   31925: result <= 12'b000010100101;
   31926: result <= 12'b000010100101;
   31927: result <= 12'b000010100100;
   31928: result <= 12'b000010100100;
   31929: result <= 12'b000010100100;
   31930: result <= 12'b000010100100;
   31931: result <= 12'b000010100100;
   31932: result <= 12'b000010100011;
   31933: result <= 12'b000010100011;
   31934: result <= 12'b000010100011;
   31935: result <= 12'b000010100011;
   31936: result <= 12'b000010100011;
   31937: result <= 12'b000010100010;
   31938: result <= 12'b000010100010;
   31939: result <= 12'b000010100010;
   31940: result <= 12'b000010100010;
   31941: result <= 12'b000010100010;
   31942: result <= 12'b000010100010;
   31943: result <= 12'b000010100001;
   31944: result <= 12'b000010100001;
   31945: result <= 12'b000010100001;
   31946: result <= 12'b000010100001;
   31947: result <= 12'b000010100001;
   31948: result <= 12'b000010100000;
   31949: result <= 12'b000010100000;
   31950: result <= 12'b000010100000;
   31951: result <= 12'b000010100000;
   31952: result <= 12'b000010100000;
   31953: result <= 12'b000010011111;
   31954: result <= 12'b000010011111;
   31955: result <= 12'b000010011111;
   31956: result <= 12'b000010011111;
   31957: result <= 12'b000010011111;
   31958: result <= 12'b000010011110;
   31959: result <= 12'b000010011110;
   31960: result <= 12'b000010011110;
   31961: result <= 12'b000010011110;
   31962: result <= 12'b000010011110;
   31963: result <= 12'b000010011101;
   31964: result <= 12'b000010011101;
   31965: result <= 12'b000010011101;
   31966: result <= 12'b000010011101;
   31967: result <= 12'b000010011101;
   31968: result <= 12'b000010011100;
   31969: result <= 12'b000010011100;
   31970: result <= 12'b000010011100;
   31971: result <= 12'b000010011100;
   31972: result <= 12'b000010011100;
   31973: result <= 12'b000010011011;
   31974: result <= 12'b000010011011;
   31975: result <= 12'b000010011011;
   31976: result <= 12'b000010011011;
   31977: result <= 12'b000010011011;
   31978: result <= 12'b000010011010;
   31979: result <= 12'b000010011010;
   31980: result <= 12'b000010011010;
   31981: result <= 12'b000010011010;
   31982: result <= 12'b000010011010;
   31983: result <= 12'b000010011001;
   31984: result <= 12'b000010011001;
   31985: result <= 12'b000010011001;
   31986: result <= 12'b000010011001;
   31987: result <= 12'b000010011001;
   31988: result <= 12'b000010011001;
   31989: result <= 12'b000010011000;
   31990: result <= 12'b000010011000;
   31991: result <= 12'b000010011000;
   31992: result <= 12'b000010011000;
   31993: result <= 12'b000010011000;
   31994: result <= 12'b000010010111;
   31995: result <= 12'b000010010111;
   31996: result <= 12'b000010010111;
   31997: result <= 12'b000010010111;
   31998: result <= 12'b000010010111;
   31999: result <= 12'b000010010110;
   32000: result <= 12'b000010010110;
   32001: result <= 12'b000010010110;
   32002: result <= 12'b000010010110;
   32003: result <= 12'b000010010110;
   32004: result <= 12'b000010010101;
   32005: result <= 12'b000010010101;
   32006: result <= 12'b000010010101;
   32007: result <= 12'b000010010101;
   32008: result <= 12'b000010010101;
   32009: result <= 12'b000010010100;
   32010: result <= 12'b000010010100;
   32011: result <= 12'b000010010100;
   32012: result <= 12'b000010010100;
   32013: result <= 12'b000010010100;
   32014: result <= 12'b000010010011;
   32015: result <= 12'b000010010011;
   32016: result <= 12'b000010010011;
   32017: result <= 12'b000010010011;
   32018: result <= 12'b000010010011;
   32019: result <= 12'b000010010010;
   32020: result <= 12'b000010010010;
   32021: result <= 12'b000010010010;
   32022: result <= 12'b000010010010;
   32023: result <= 12'b000010010010;
   32024: result <= 12'b000010010001;
   32025: result <= 12'b000010010001;
   32026: result <= 12'b000010010001;
   32027: result <= 12'b000010010001;
   32028: result <= 12'b000010010001;
   32029: result <= 12'b000010010000;
   32030: result <= 12'b000010010000;
   32031: result <= 12'b000010010000;
   32032: result <= 12'b000010010000;
   32033: result <= 12'b000010010000;
   32034: result <= 12'b000010010000;
   32035: result <= 12'b000010001111;
   32036: result <= 12'b000010001111;
   32037: result <= 12'b000010001111;
   32038: result <= 12'b000010001111;
   32039: result <= 12'b000010001111;
   32040: result <= 12'b000010001110;
   32041: result <= 12'b000010001110;
   32042: result <= 12'b000010001110;
   32043: result <= 12'b000010001110;
   32044: result <= 12'b000010001110;
   32045: result <= 12'b000010001101;
   32046: result <= 12'b000010001101;
   32047: result <= 12'b000010001101;
   32048: result <= 12'b000010001101;
   32049: result <= 12'b000010001101;
   32050: result <= 12'b000010001100;
   32051: result <= 12'b000010001100;
   32052: result <= 12'b000010001100;
   32053: result <= 12'b000010001100;
   32054: result <= 12'b000010001100;
   32055: result <= 12'b000010001011;
   32056: result <= 12'b000010001011;
   32057: result <= 12'b000010001011;
   32058: result <= 12'b000010001011;
   32059: result <= 12'b000010001011;
   32060: result <= 12'b000010001010;
   32061: result <= 12'b000010001010;
   32062: result <= 12'b000010001010;
   32063: result <= 12'b000010001010;
   32064: result <= 12'b000010001010;
   32065: result <= 12'b000010001001;
   32066: result <= 12'b000010001001;
   32067: result <= 12'b000010001001;
   32068: result <= 12'b000010001001;
   32069: result <= 12'b000010001001;
   32070: result <= 12'b000010001000;
   32071: result <= 12'b000010001000;
   32072: result <= 12'b000010001000;
   32073: result <= 12'b000010001000;
   32074: result <= 12'b000010001000;
   32075: result <= 12'b000010000111;
   32076: result <= 12'b000010000111;
   32077: result <= 12'b000010000111;
   32078: result <= 12'b000010000111;
   32079: result <= 12'b000010000111;
   32080: result <= 12'b000010000110;
   32081: result <= 12'b000010000110;
   32082: result <= 12'b000010000110;
   32083: result <= 12'b000010000110;
   32084: result <= 12'b000010000110;
   32085: result <= 12'b000010000110;
   32086: result <= 12'b000010000101;
   32087: result <= 12'b000010000101;
   32088: result <= 12'b000010000101;
   32089: result <= 12'b000010000101;
   32090: result <= 12'b000010000101;
   32091: result <= 12'b000010000100;
   32092: result <= 12'b000010000100;
   32093: result <= 12'b000010000100;
   32094: result <= 12'b000010000100;
   32095: result <= 12'b000010000100;
   32096: result <= 12'b000010000011;
   32097: result <= 12'b000010000011;
   32098: result <= 12'b000010000011;
   32099: result <= 12'b000010000011;
   32100: result <= 12'b000010000011;
   32101: result <= 12'b000010000010;
   32102: result <= 12'b000010000010;
   32103: result <= 12'b000010000010;
   32104: result <= 12'b000010000010;
   32105: result <= 12'b000010000010;
   32106: result <= 12'b000010000001;
   32107: result <= 12'b000010000001;
   32108: result <= 12'b000010000001;
   32109: result <= 12'b000010000001;
   32110: result <= 12'b000010000001;
   32111: result <= 12'b000010000000;
   32112: result <= 12'b000010000000;
   32113: result <= 12'b000010000000;
   32114: result <= 12'b000010000000;
   32115: result <= 12'b000010000000;
   32116: result <= 12'b000001111111;
   32117: result <= 12'b000001111111;
   32118: result <= 12'b000001111111;
   32119: result <= 12'b000001111111;
   32120: result <= 12'b000001111111;
   32121: result <= 12'b000001111110;
   32122: result <= 12'b000001111110;
   32123: result <= 12'b000001111110;
   32124: result <= 12'b000001111110;
   32125: result <= 12'b000001111110;
   32126: result <= 12'b000001111101;
   32127: result <= 12'b000001111101;
   32128: result <= 12'b000001111101;
   32129: result <= 12'b000001111101;
   32130: result <= 12'b000001111101;
   32131: result <= 12'b000001111100;
   32132: result <= 12'b000001111100;
   32133: result <= 12'b000001111100;
   32134: result <= 12'b000001111100;
   32135: result <= 12'b000001111100;
   32136: result <= 12'b000001111100;
   32137: result <= 12'b000001111011;
   32138: result <= 12'b000001111011;
   32139: result <= 12'b000001111011;
   32140: result <= 12'b000001111011;
   32141: result <= 12'b000001111011;
   32142: result <= 12'b000001111010;
   32143: result <= 12'b000001111010;
   32144: result <= 12'b000001111010;
   32145: result <= 12'b000001111010;
   32146: result <= 12'b000001111010;
   32147: result <= 12'b000001111001;
   32148: result <= 12'b000001111001;
   32149: result <= 12'b000001111001;
   32150: result <= 12'b000001111001;
   32151: result <= 12'b000001111001;
   32152: result <= 12'b000001111000;
   32153: result <= 12'b000001111000;
   32154: result <= 12'b000001111000;
   32155: result <= 12'b000001111000;
   32156: result <= 12'b000001111000;
   32157: result <= 12'b000001110111;
   32158: result <= 12'b000001110111;
   32159: result <= 12'b000001110111;
   32160: result <= 12'b000001110111;
   32161: result <= 12'b000001110111;
   32162: result <= 12'b000001110110;
   32163: result <= 12'b000001110110;
   32164: result <= 12'b000001110110;
   32165: result <= 12'b000001110110;
   32166: result <= 12'b000001110110;
   32167: result <= 12'b000001110101;
   32168: result <= 12'b000001110101;
   32169: result <= 12'b000001110101;
   32170: result <= 12'b000001110101;
   32171: result <= 12'b000001110101;
   32172: result <= 12'b000001110100;
   32173: result <= 12'b000001110100;
   32174: result <= 12'b000001110100;
   32175: result <= 12'b000001110100;
   32176: result <= 12'b000001110100;
   32177: result <= 12'b000001110011;
   32178: result <= 12'b000001110011;
   32179: result <= 12'b000001110011;
   32180: result <= 12'b000001110011;
   32181: result <= 12'b000001110011;
   32182: result <= 12'b000001110011;
   32183: result <= 12'b000001110010;
   32184: result <= 12'b000001110010;
   32185: result <= 12'b000001110010;
   32186: result <= 12'b000001110010;
   32187: result <= 12'b000001110010;
   32188: result <= 12'b000001110001;
   32189: result <= 12'b000001110001;
   32190: result <= 12'b000001110001;
   32191: result <= 12'b000001110001;
   32192: result <= 12'b000001110001;
   32193: result <= 12'b000001110000;
   32194: result <= 12'b000001110000;
   32195: result <= 12'b000001110000;
   32196: result <= 12'b000001110000;
   32197: result <= 12'b000001110000;
   32198: result <= 12'b000001101111;
   32199: result <= 12'b000001101111;
   32200: result <= 12'b000001101111;
   32201: result <= 12'b000001101111;
   32202: result <= 12'b000001101111;
   32203: result <= 12'b000001101110;
   32204: result <= 12'b000001101110;
   32205: result <= 12'b000001101110;
   32206: result <= 12'b000001101110;
   32207: result <= 12'b000001101110;
   32208: result <= 12'b000001101101;
   32209: result <= 12'b000001101101;
   32210: result <= 12'b000001101101;
   32211: result <= 12'b000001101101;
   32212: result <= 12'b000001101101;
   32213: result <= 12'b000001101100;
   32214: result <= 12'b000001101100;
   32215: result <= 12'b000001101100;
   32216: result <= 12'b000001101100;
   32217: result <= 12'b000001101100;
   32218: result <= 12'b000001101011;
   32219: result <= 12'b000001101011;
   32220: result <= 12'b000001101011;
   32221: result <= 12'b000001101011;
   32222: result <= 12'b000001101011;
   32223: result <= 12'b000001101010;
   32224: result <= 12'b000001101010;
   32225: result <= 12'b000001101010;
   32226: result <= 12'b000001101010;
   32227: result <= 12'b000001101010;
   32228: result <= 12'b000001101001;
   32229: result <= 12'b000001101001;
   32230: result <= 12'b000001101001;
   32231: result <= 12'b000001101001;
   32232: result <= 12'b000001101001;
   32233: result <= 12'b000001101001;
   32234: result <= 12'b000001101000;
   32235: result <= 12'b000001101000;
   32236: result <= 12'b000001101000;
   32237: result <= 12'b000001101000;
   32238: result <= 12'b000001101000;
   32239: result <= 12'b000001100111;
   32240: result <= 12'b000001100111;
   32241: result <= 12'b000001100111;
   32242: result <= 12'b000001100111;
   32243: result <= 12'b000001100111;
   32244: result <= 12'b000001100110;
   32245: result <= 12'b000001100110;
   32246: result <= 12'b000001100110;
   32247: result <= 12'b000001100110;
   32248: result <= 12'b000001100110;
   32249: result <= 12'b000001100101;
   32250: result <= 12'b000001100101;
   32251: result <= 12'b000001100101;
   32252: result <= 12'b000001100101;
   32253: result <= 12'b000001100101;
   32254: result <= 12'b000001100100;
   32255: result <= 12'b000001100100;
   32256: result <= 12'b000001100100;
   32257: result <= 12'b000001100100;
   32258: result <= 12'b000001100100;
   32259: result <= 12'b000001100011;
   32260: result <= 12'b000001100011;
   32261: result <= 12'b000001100011;
   32262: result <= 12'b000001100011;
   32263: result <= 12'b000001100011;
   32264: result <= 12'b000001100010;
   32265: result <= 12'b000001100010;
   32266: result <= 12'b000001100010;
   32267: result <= 12'b000001100010;
   32268: result <= 12'b000001100010;
   32269: result <= 12'b000001100001;
   32270: result <= 12'b000001100001;
   32271: result <= 12'b000001100001;
   32272: result <= 12'b000001100001;
   32273: result <= 12'b000001100001;
   32274: result <= 12'b000001100000;
   32275: result <= 12'b000001100000;
   32276: result <= 12'b000001100000;
   32277: result <= 12'b000001100000;
   32278: result <= 12'b000001100000;
   32279: result <= 12'b000001011111;
   32280: result <= 12'b000001011111;
   32281: result <= 12'b000001011111;
   32282: result <= 12'b000001011111;
   32283: result <= 12'b000001011111;
   32284: result <= 12'b000001011110;
   32285: result <= 12'b000001011110;
   32286: result <= 12'b000001011110;
   32287: result <= 12'b000001011110;
   32288: result <= 12'b000001011110;
   32289: result <= 12'b000001011110;
   32290: result <= 12'b000001011101;
   32291: result <= 12'b000001011101;
   32292: result <= 12'b000001011101;
   32293: result <= 12'b000001011101;
   32294: result <= 12'b000001011101;
   32295: result <= 12'b000001011100;
   32296: result <= 12'b000001011100;
   32297: result <= 12'b000001011100;
   32298: result <= 12'b000001011100;
   32299: result <= 12'b000001011100;
   32300: result <= 12'b000001011011;
   32301: result <= 12'b000001011011;
   32302: result <= 12'b000001011011;
   32303: result <= 12'b000001011011;
   32304: result <= 12'b000001011011;
   32305: result <= 12'b000001011010;
   32306: result <= 12'b000001011010;
   32307: result <= 12'b000001011010;
   32308: result <= 12'b000001011010;
   32309: result <= 12'b000001011010;
   32310: result <= 12'b000001011001;
   32311: result <= 12'b000001011001;
   32312: result <= 12'b000001011001;
   32313: result <= 12'b000001011001;
   32314: result <= 12'b000001011001;
   32315: result <= 12'b000001011000;
   32316: result <= 12'b000001011000;
   32317: result <= 12'b000001011000;
   32318: result <= 12'b000001011000;
   32319: result <= 12'b000001011000;
   32320: result <= 12'b000001010111;
   32321: result <= 12'b000001010111;
   32322: result <= 12'b000001010111;
   32323: result <= 12'b000001010111;
   32324: result <= 12'b000001010111;
   32325: result <= 12'b000001010110;
   32326: result <= 12'b000001010110;
   32327: result <= 12'b000001010110;
   32328: result <= 12'b000001010110;
   32329: result <= 12'b000001010110;
   32330: result <= 12'b000001010101;
   32331: result <= 12'b000001010101;
   32332: result <= 12'b000001010101;
   32333: result <= 12'b000001010101;
   32334: result <= 12'b000001010101;
   32335: result <= 12'b000001010100;
   32336: result <= 12'b000001010100;
   32337: result <= 12'b000001010100;
   32338: result <= 12'b000001010100;
   32339: result <= 12'b000001010100;
   32340: result <= 12'b000001010100;
   32341: result <= 12'b000001010011;
   32342: result <= 12'b000001010011;
   32343: result <= 12'b000001010011;
   32344: result <= 12'b000001010011;
   32345: result <= 12'b000001010011;
   32346: result <= 12'b000001010010;
   32347: result <= 12'b000001010010;
   32348: result <= 12'b000001010010;
   32349: result <= 12'b000001010010;
   32350: result <= 12'b000001010010;
   32351: result <= 12'b000001010001;
   32352: result <= 12'b000001010001;
   32353: result <= 12'b000001010001;
   32354: result <= 12'b000001010001;
   32355: result <= 12'b000001010001;
   32356: result <= 12'b000001010000;
   32357: result <= 12'b000001010000;
   32358: result <= 12'b000001010000;
   32359: result <= 12'b000001010000;
   32360: result <= 12'b000001010000;
   32361: result <= 12'b000001001111;
   32362: result <= 12'b000001001111;
   32363: result <= 12'b000001001111;
   32364: result <= 12'b000001001111;
   32365: result <= 12'b000001001111;
   32366: result <= 12'b000001001110;
   32367: result <= 12'b000001001110;
   32368: result <= 12'b000001001110;
   32369: result <= 12'b000001001110;
   32370: result <= 12'b000001001110;
   32371: result <= 12'b000001001101;
   32372: result <= 12'b000001001101;
   32373: result <= 12'b000001001101;
   32374: result <= 12'b000001001101;
   32375: result <= 12'b000001001101;
   32376: result <= 12'b000001001100;
   32377: result <= 12'b000001001100;
   32378: result <= 12'b000001001100;
   32379: result <= 12'b000001001100;
   32380: result <= 12'b000001001100;
   32381: result <= 12'b000001001011;
   32382: result <= 12'b000001001011;
   32383: result <= 12'b000001001011;
   32384: result <= 12'b000001001011;
   32385: result <= 12'b000001001011;
   32386: result <= 12'b000001001010;
   32387: result <= 12'b000001001010;
   32388: result <= 12'b000001001010;
   32389: result <= 12'b000001001010;
   32390: result <= 12'b000001001010;
   32391: result <= 12'b000001001010;
   32392: result <= 12'b000001001001;
   32393: result <= 12'b000001001001;
   32394: result <= 12'b000001001001;
   32395: result <= 12'b000001001001;
   32396: result <= 12'b000001001001;
   32397: result <= 12'b000001001000;
   32398: result <= 12'b000001001000;
   32399: result <= 12'b000001001000;
   32400: result <= 12'b000001001000;
   32401: result <= 12'b000001001000;
   32402: result <= 12'b000001000111;
   32403: result <= 12'b000001000111;
   32404: result <= 12'b000001000111;
   32405: result <= 12'b000001000111;
   32406: result <= 12'b000001000111;
   32407: result <= 12'b000001000110;
   32408: result <= 12'b000001000110;
   32409: result <= 12'b000001000110;
   32410: result <= 12'b000001000110;
   32411: result <= 12'b000001000110;
   32412: result <= 12'b000001000101;
   32413: result <= 12'b000001000101;
   32414: result <= 12'b000001000101;
   32415: result <= 12'b000001000101;
   32416: result <= 12'b000001000101;
   32417: result <= 12'b000001000100;
   32418: result <= 12'b000001000100;
   32419: result <= 12'b000001000100;
   32420: result <= 12'b000001000100;
   32421: result <= 12'b000001000100;
   32422: result <= 12'b000001000011;
   32423: result <= 12'b000001000011;
   32424: result <= 12'b000001000011;
   32425: result <= 12'b000001000011;
   32426: result <= 12'b000001000011;
   32427: result <= 12'b000001000010;
   32428: result <= 12'b000001000010;
   32429: result <= 12'b000001000010;
   32430: result <= 12'b000001000010;
   32431: result <= 12'b000001000010;
   32432: result <= 12'b000001000001;
   32433: result <= 12'b000001000001;
   32434: result <= 12'b000001000001;
   32435: result <= 12'b000001000001;
   32436: result <= 12'b000001000001;
   32437: result <= 12'b000001000000;
   32438: result <= 12'b000001000000;
   32439: result <= 12'b000001000000;
   32440: result <= 12'b000001000000;
   32441: result <= 12'b000001000000;
   32442: result <= 12'b000000111111;
   32443: result <= 12'b000000111111;
   32444: result <= 12'b000000111111;
   32445: result <= 12'b000000111111;
   32446: result <= 12'b000000111111;
   32447: result <= 12'b000000111111;
   32448: result <= 12'b000000111110;
   32449: result <= 12'b000000111110;
   32450: result <= 12'b000000111110;
   32451: result <= 12'b000000111110;
   32452: result <= 12'b000000111110;
   32453: result <= 12'b000000111101;
   32454: result <= 12'b000000111101;
   32455: result <= 12'b000000111101;
   32456: result <= 12'b000000111101;
   32457: result <= 12'b000000111101;
   32458: result <= 12'b000000111100;
   32459: result <= 12'b000000111100;
   32460: result <= 12'b000000111100;
   32461: result <= 12'b000000111100;
   32462: result <= 12'b000000111100;
   32463: result <= 12'b000000111011;
   32464: result <= 12'b000000111011;
   32465: result <= 12'b000000111011;
   32466: result <= 12'b000000111011;
   32467: result <= 12'b000000111011;
   32468: result <= 12'b000000111010;
   32469: result <= 12'b000000111010;
   32470: result <= 12'b000000111010;
   32471: result <= 12'b000000111010;
   32472: result <= 12'b000000111010;
   32473: result <= 12'b000000111001;
   32474: result <= 12'b000000111001;
   32475: result <= 12'b000000111001;
   32476: result <= 12'b000000111001;
   32477: result <= 12'b000000111001;
   32478: result <= 12'b000000111000;
   32479: result <= 12'b000000111000;
   32480: result <= 12'b000000111000;
   32481: result <= 12'b000000111000;
   32482: result <= 12'b000000111000;
   32483: result <= 12'b000000110111;
   32484: result <= 12'b000000110111;
   32485: result <= 12'b000000110111;
   32486: result <= 12'b000000110111;
   32487: result <= 12'b000000110111;
   32488: result <= 12'b000000110110;
   32489: result <= 12'b000000110110;
   32490: result <= 12'b000000110110;
   32491: result <= 12'b000000110110;
   32492: result <= 12'b000000110110;
   32493: result <= 12'b000000110101;
   32494: result <= 12'b000000110101;
   32495: result <= 12'b000000110101;
   32496: result <= 12'b000000110101;
   32497: result <= 12'b000000110101;
   32498: result <= 12'b000000110101;
   32499: result <= 12'b000000110100;
   32500: result <= 12'b000000110100;
   32501: result <= 12'b000000110100;
   32502: result <= 12'b000000110100;
   32503: result <= 12'b000000110100;
   32504: result <= 12'b000000110011;
   32505: result <= 12'b000000110011;
   32506: result <= 12'b000000110011;
   32507: result <= 12'b000000110011;
   32508: result <= 12'b000000110011;
   32509: result <= 12'b000000110010;
   32510: result <= 12'b000000110010;
   32511: result <= 12'b000000110010;
   32512: result <= 12'b000000110010;
   32513: result <= 12'b000000110010;
   32514: result <= 12'b000000110001;
   32515: result <= 12'b000000110001;
   32516: result <= 12'b000000110001;
   32517: result <= 12'b000000110001;
   32518: result <= 12'b000000110001;
   32519: result <= 12'b000000110000;
   32520: result <= 12'b000000110000;
   32521: result <= 12'b000000110000;
   32522: result <= 12'b000000110000;
   32523: result <= 12'b000000110000;
   32524: result <= 12'b000000101111;
   32525: result <= 12'b000000101111;
   32526: result <= 12'b000000101111;
   32527: result <= 12'b000000101111;
   32528: result <= 12'b000000101111;
   32529: result <= 12'b000000101110;
   32530: result <= 12'b000000101110;
   32531: result <= 12'b000000101110;
   32532: result <= 12'b000000101110;
   32533: result <= 12'b000000101110;
   32534: result <= 12'b000000101101;
   32535: result <= 12'b000000101101;
   32536: result <= 12'b000000101101;
   32537: result <= 12'b000000101101;
   32538: result <= 12'b000000101101;
   32539: result <= 12'b000000101100;
   32540: result <= 12'b000000101100;
   32541: result <= 12'b000000101100;
   32542: result <= 12'b000000101100;
   32543: result <= 12'b000000101100;
   32544: result <= 12'b000000101011;
   32545: result <= 12'b000000101011;
   32546: result <= 12'b000000101011;
   32547: result <= 12'b000000101011;
   32548: result <= 12'b000000101011;
   32549: result <= 12'b000000101010;
   32550: result <= 12'b000000101010;
   32551: result <= 12'b000000101010;
   32552: result <= 12'b000000101010;
   32553: result <= 12'b000000101010;
   32554: result <= 12'b000000101010;
   32555: result <= 12'b000000101001;
   32556: result <= 12'b000000101001;
   32557: result <= 12'b000000101001;
   32558: result <= 12'b000000101001;
   32559: result <= 12'b000000101001;
   32560: result <= 12'b000000101000;
   32561: result <= 12'b000000101000;
   32562: result <= 12'b000000101000;
   32563: result <= 12'b000000101000;
   32564: result <= 12'b000000101000;
   32565: result <= 12'b000000100111;
   32566: result <= 12'b000000100111;
   32567: result <= 12'b000000100111;
   32568: result <= 12'b000000100111;
   32569: result <= 12'b000000100111;
   32570: result <= 12'b000000100110;
   32571: result <= 12'b000000100110;
   32572: result <= 12'b000000100110;
   32573: result <= 12'b000000100110;
   32574: result <= 12'b000000100110;
   32575: result <= 12'b000000100101;
   32576: result <= 12'b000000100101;
   32577: result <= 12'b000000100101;
   32578: result <= 12'b000000100101;
   32579: result <= 12'b000000100101;
   32580: result <= 12'b000000100100;
   32581: result <= 12'b000000100100;
   32582: result <= 12'b000000100100;
   32583: result <= 12'b000000100100;
   32584: result <= 12'b000000100100;
   32585: result <= 12'b000000100011;
   32586: result <= 12'b000000100011;
   32587: result <= 12'b000000100011;
   32588: result <= 12'b000000100011;
   32589: result <= 12'b000000100011;
   32590: result <= 12'b000000100010;
   32591: result <= 12'b000000100010;
   32592: result <= 12'b000000100010;
   32593: result <= 12'b000000100010;
   32594: result <= 12'b000000100010;
   32595: result <= 12'b000000100001;
   32596: result <= 12'b000000100001;
   32597: result <= 12'b000000100001;
   32598: result <= 12'b000000100001;
   32599: result <= 12'b000000100001;
   32600: result <= 12'b000000100000;
   32601: result <= 12'b000000100000;
   32602: result <= 12'b000000100000;
   32603: result <= 12'b000000100000;
   32604: result <= 12'b000000100000;
   32605: result <= 12'b000000100000;
   32606: result <= 12'b000000011111;
   32607: result <= 12'b000000011111;
   32608: result <= 12'b000000011111;
   32609: result <= 12'b000000011111;
   32610: result <= 12'b000000011111;
   32611: result <= 12'b000000011110;
   32612: result <= 12'b000000011110;
   32613: result <= 12'b000000011110;
   32614: result <= 12'b000000011110;
   32615: result <= 12'b000000011110;
   32616: result <= 12'b000000011101;
   32617: result <= 12'b000000011101;
   32618: result <= 12'b000000011101;
   32619: result <= 12'b000000011101;
   32620: result <= 12'b000000011101;
   32621: result <= 12'b000000011100;
   32622: result <= 12'b000000011100;
   32623: result <= 12'b000000011100;
   32624: result <= 12'b000000011100;
   32625: result <= 12'b000000011100;
   32626: result <= 12'b000000011011;
   32627: result <= 12'b000000011011;
   32628: result <= 12'b000000011011;
   32629: result <= 12'b000000011011;
   32630: result <= 12'b000000011011;
   32631: result <= 12'b000000011010;
   32632: result <= 12'b000000011010;
   32633: result <= 12'b000000011010;
   32634: result <= 12'b000000011010;
   32635: result <= 12'b000000011010;
   32636: result <= 12'b000000011001;
   32637: result <= 12'b000000011001;
   32638: result <= 12'b000000011001;
   32639: result <= 12'b000000011001;
   32640: result <= 12'b000000011001;
   32641: result <= 12'b000000011000;
   32642: result <= 12'b000000011000;
   32643: result <= 12'b000000011000;
   32644: result <= 12'b000000011000;
   32645: result <= 12'b000000011000;
   32646: result <= 12'b000000010111;
   32647: result <= 12'b000000010111;
   32648: result <= 12'b000000010111;
   32649: result <= 12'b000000010111;
   32650: result <= 12'b000000010111;
   32651: result <= 12'b000000010110;
   32652: result <= 12'b000000010110;
   32653: result <= 12'b000000010110;
   32654: result <= 12'b000000010110;
   32655: result <= 12'b000000010110;
   32656: result <= 12'b000000010101;
   32657: result <= 12'b000000010101;
   32658: result <= 12'b000000010101;
   32659: result <= 12'b000000010101;
   32660: result <= 12'b000000010101;
   32661: result <= 12'b000000010101;
   32662: result <= 12'b000000010100;
   32663: result <= 12'b000000010100;
   32664: result <= 12'b000000010100;
   32665: result <= 12'b000000010100;
   32666: result <= 12'b000000010100;
   32667: result <= 12'b000000010011;
   32668: result <= 12'b000000010011;
   32669: result <= 12'b000000010011;
   32670: result <= 12'b000000010011;
   32671: result <= 12'b000000010011;
   32672: result <= 12'b000000010010;
   32673: result <= 12'b000000010010;
   32674: result <= 12'b000000010010;
   32675: result <= 12'b000000010010;
   32676: result <= 12'b000000010010;
   32677: result <= 12'b000000010001;
   32678: result <= 12'b000000010001;
   32679: result <= 12'b000000010001;
   32680: result <= 12'b000000010001;
   32681: result <= 12'b000000010001;
   32682: result <= 12'b000000010000;
   32683: result <= 12'b000000010000;
   32684: result <= 12'b000000010000;
   32685: result <= 12'b000000010000;
   32686: result <= 12'b000000010000;
   32687: result <= 12'b000000001111;
   32688: result <= 12'b000000001111;
   32689: result <= 12'b000000001111;
   32690: result <= 12'b000000001111;
   32691: result <= 12'b000000001111;
   32692: result <= 12'b000000001110;
   32693: result <= 12'b000000001110;
   32694: result <= 12'b000000001110;
   32695: result <= 12'b000000001110;
   32696: result <= 12'b000000001110;
   32697: result <= 12'b000000001101;
   32698: result <= 12'b000000001101;
   32699: result <= 12'b000000001101;
   32700: result <= 12'b000000001101;
   32701: result <= 12'b000000001101;
   32702: result <= 12'b000000001100;
   32703: result <= 12'b000000001100;
   32704: result <= 12'b000000001100;
   32705: result <= 12'b000000001100;
   32706: result <= 12'b000000001100;
   32707: result <= 12'b000000001011;
   32708: result <= 12'b000000001011;
   32709: result <= 12'b000000001011;
   32710: result <= 12'b000000001011;
   32711: result <= 12'b000000001011;
   32712: result <= 12'b000000001010;
   32713: result <= 12'b000000001010;
   32714: result <= 12'b000000001010;
   32715: result <= 12'b000000001010;
   32716: result <= 12'b000000001010;
   32717: result <= 12'b000000001010;
   32718: result <= 12'b000000001001;
   32719: result <= 12'b000000001001;
   32720: result <= 12'b000000001001;
   32721: result <= 12'b000000001001;
   32722: result <= 12'b000000001001;
   32723: result <= 12'b000000001000;
   32724: result <= 12'b000000001000;
   32725: result <= 12'b000000001000;
   32726: result <= 12'b000000001000;
   32727: result <= 12'b000000001000;
   32728: result <= 12'b000000000111;
   32729: result <= 12'b000000000111;
   32730: result <= 12'b000000000111;
   32731: result <= 12'b000000000111;
   32732: result <= 12'b000000000111;
   32733: result <= 12'b000000000110;
   32734: result <= 12'b000000000110;
   32735: result <= 12'b000000000110;
   32736: result <= 12'b000000000110;
   32737: result <= 12'b000000000110;
   32738: result <= 12'b000000000101;
   32739: result <= 12'b000000000101;
   32740: result <= 12'b000000000101;
   32741: result <= 12'b000000000101;
   32742: result <= 12'b000000000101;
   32743: result <= 12'b000000000100;
   32744: result <= 12'b000000000100;
   32745: result <= 12'b000000000100;
   32746: result <= 12'b000000000100;
   32747: result <= 12'b000000000100;
   32748: result <= 12'b000000000011;
   32749: result <= 12'b000000000011;
   32750: result <= 12'b000000000011;
   32751: result <= 12'b000000000011;
   32752: result <= 12'b000000000011;
   32753: result <= 12'b000000000010;
   32754: result <= 12'b000000000010;
   32755: result <= 12'b000000000010;
   32756: result <= 12'b000000000010;
   32757: result <= 12'b000000000010;
   32758: result <= 12'b000000000001;
   32759: result <= 12'b000000000001;
   32760: result <= 12'b000000000001;
   32761: result <= 12'b000000000001;
   32762: result <= 12'b000000000001;
   32763: result <= 12'b000000000000;
   32764: result <= 12'b000000000000;
   32765: result <= 12'b000000000000;
   32766: result <= 12'b000000000000;
   32767: result <= 12'b000000000000;
   32768: result <= 12'b000000000000;
   32769: result <= 12'b000000000000;
   32770: result <= 12'b000000000000;
   32771: result <= 12'b000000000000;
   32772: result <= 12'b000000000000;
   32773: result <= 12'b000000000000;
   32774: result <= 12'b111111111111;
   32775: result <= 12'b111111111111;
   32776: result <= 12'b111111111111;
   32777: result <= 12'b111111111111;
   32778: result <= 12'b111111111111;
   32779: result <= 12'b111111111110;
   32780: result <= 12'b111111111110;
   32781: result <= 12'b111111111110;
   32782: result <= 12'b111111111110;
   32783: result <= 12'b111111111110;
   32784: result <= 12'b111111111111;
   32785: result <= 12'b111111111111;
   32786: result <= 12'b111111111111;
   32787: result <= 12'b111111111111;
   32788: result <= 12'b111111111111;
   32789: result <= 12'b111111111100;
   32790: result <= 12'b111111111100;
   32791: result <= 12'b111111111100;
   32792: result <= 12'b111111111100;
   32793: result <= 12'b111111111100;
   32794: result <= 12'b111111111101;
   32795: result <= 12'b111111111101;
   32796: result <= 12'b111111111101;
   32797: result <= 12'b111111111101;
   32798: result <= 12'b111111111101;
   32799: result <= 12'b111111111110;
   32800: result <= 12'b111111111110;
   32801: result <= 12'b111111111110;
   32802: result <= 12'b111111111110;
   32803: result <= 12'b111111111110;
   32804: result <= 12'b111111111111;
   32805: result <= 12'b111111111111;
   32806: result <= 12'b111111111111;
   32807: result <= 12'b111111111111;
   32808: result <= 12'b111111111111;
   32809: result <= 12'b111111111000;
   32810: result <= 12'b111111111000;
   32811: result <= 12'b111111111000;
   32812: result <= 12'b111111111000;
   32813: result <= 12'b111111111000;
   32814: result <= 12'b111111111001;
   32815: result <= 12'b111111111001;
   32816: result <= 12'b111111111001;
   32817: result <= 12'b111111111001;
   32818: result <= 12'b111111111001;
   32819: result <= 12'b111111111010;
   32820: result <= 12'b111111111010;
   32821: result <= 12'b111111111010;
   32822: result <= 12'b111111111010;
   32823: result <= 12'b111111111010;
   32824: result <= 12'b111111111010;
   32825: result <= 12'b111111111011;
   32826: result <= 12'b111111111011;
   32827: result <= 12'b111111111011;
   32828: result <= 12'b111111111011;
   32829: result <= 12'b111111111011;
   32830: result <= 12'b111111111100;
   32831: result <= 12'b111111111100;
   32832: result <= 12'b111111111100;
   32833: result <= 12'b111111111100;
   32834: result <= 12'b111111111100;
   32835: result <= 12'b111111111101;
   32836: result <= 12'b111111111101;
   32837: result <= 12'b111111111101;
   32838: result <= 12'b111111111101;
   32839: result <= 12'b111111111101;
   32840: result <= 12'b111111111110;
   32841: result <= 12'b111111111110;
   32842: result <= 12'b111111111110;
   32843: result <= 12'b111111111110;
   32844: result <= 12'b111111111110;
   32845: result <= 12'b111111111111;
   32846: result <= 12'b111111111111;
   32847: result <= 12'b111111111111;
   32848: result <= 12'b111111111111;
   32849: result <= 12'b111111111111;
   32850: result <= 12'b111111110000;
   32851: result <= 12'b111111110000;
   32852: result <= 12'b111111110000;
   32853: result <= 12'b111111110000;
   32854: result <= 12'b111111110000;
   32855: result <= 12'b111111110001;
   32856: result <= 12'b111111110001;
   32857: result <= 12'b111111110001;
   32858: result <= 12'b111111110001;
   32859: result <= 12'b111111110001;
   32860: result <= 12'b111111110010;
   32861: result <= 12'b111111110010;
   32862: result <= 12'b111111110010;
   32863: result <= 12'b111111110010;
   32864: result <= 12'b111111110010;
   32865: result <= 12'b111111110011;
   32866: result <= 12'b111111110011;
   32867: result <= 12'b111111110011;
   32868: result <= 12'b111111110011;
   32869: result <= 12'b111111110011;
   32870: result <= 12'b111111110100;
   32871: result <= 12'b111111110100;
   32872: result <= 12'b111111110100;
   32873: result <= 12'b111111110100;
   32874: result <= 12'b111111110100;
   32875: result <= 12'b111111110101;
   32876: result <= 12'b111111110101;
   32877: result <= 12'b111111110101;
   32878: result <= 12'b111111110101;
   32879: result <= 12'b111111110101;
   32880: result <= 12'b111111110101;
   32881: result <= 12'b111111110110;
   32882: result <= 12'b111111110110;
   32883: result <= 12'b111111110110;
   32884: result <= 12'b111111110110;
   32885: result <= 12'b111111110110;
   32886: result <= 12'b111111110111;
   32887: result <= 12'b111111110111;
   32888: result <= 12'b111111110111;
   32889: result <= 12'b111111110111;
   32890: result <= 12'b111111110111;
   32891: result <= 12'b111111111000;
   32892: result <= 12'b111111111000;
   32893: result <= 12'b111111111000;
   32894: result <= 12'b111111111000;
   32895: result <= 12'b111111111000;
   32896: result <= 12'b111111111001;
   32897: result <= 12'b111111111001;
   32898: result <= 12'b111111111001;
   32899: result <= 12'b111111111001;
   32900: result <= 12'b111111111001;
   32901: result <= 12'b111111111010;
   32902: result <= 12'b111111111010;
   32903: result <= 12'b111111111010;
   32904: result <= 12'b111111111010;
   32905: result <= 12'b111111111010;
   32906: result <= 12'b111111111011;
   32907: result <= 12'b111111111011;
   32908: result <= 12'b111111111011;
   32909: result <= 12'b111111111011;
   32910: result <= 12'b111111111011;
   32911: result <= 12'b111111111100;
   32912: result <= 12'b111111111100;
   32913: result <= 12'b111111111100;
   32914: result <= 12'b111111111100;
   32915: result <= 12'b111111111100;
   32916: result <= 12'b111111111101;
   32917: result <= 12'b111111111101;
   32918: result <= 12'b111111111101;
   32919: result <= 12'b111111111101;
   32920: result <= 12'b111111111101;
   32921: result <= 12'b111111111110;
   32922: result <= 12'b111111111110;
   32923: result <= 12'b111111111110;
   32924: result <= 12'b111111111110;
   32925: result <= 12'b111111111110;
   32926: result <= 12'b111111111111;
   32927: result <= 12'b111111111111;
   32928: result <= 12'b111111111111;
   32929: result <= 12'b111111111111;
   32930: result <= 12'b111111111111;
   32931: result <= 12'b111111100000;
   32932: result <= 12'b111111100000;
   32933: result <= 12'b111111100000;
   32934: result <= 12'b111111100000;
   32935: result <= 12'b111111100000;
   32936: result <= 12'b111111100000;
   32937: result <= 12'b111111100001;
   32938: result <= 12'b111111100001;
   32939: result <= 12'b111111100001;
   32940: result <= 12'b111111100001;
   32941: result <= 12'b111111100001;
   32942: result <= 12'b111111100010;
   32943: result <= 12'b111111100010;
   32944: result <= 12'b111111100010;
   32945: result <= 12'b111111100010;
   32946: result <= 12'b111111100010;
   32947: result <= 12'b111111100011;
   32948: result <= 12'b111111100011;
   32949: result <= 12'b111111100011;
   32950: result <= 12'b111111100011;
   32951: result <= 12'b111111100011;
   32952: result <= 12'b111111100100;
   32953: result <= 12'b111111100100;
   32954: result <= 12'b111111100100;
   32955: result <= 12'b111111100100;
   32956: result <= 12'b111111100100;
   32957: result <= 12'b111111100101;
   32958: result <= 12'b111111100101;
   32959: result <= 12'b111111100101;
   32960: result <= 12'b111111100101;
   32961: result <= 12'b111111100101;
   32962: result <= 12'b111111100110;
   32963: result <= 12'b111111100110;
   32964: result <= 12'b111111100110;
   32965: result <= 12'b111111100110;
   32966: result <= 12'b111111100110;
   32967: result <= 12'b111111100111;
   32968: result <= 12'b111111100111;
   32969: result <= 12'b111111100111;
   32970: result <= 12'b111111100111;
   32971: result <= 12'b111111100111;
   32972: result <= 12'b111111101000;
   32973: result <= 12'b111111101000;
   32974: result <= 12'b111111101000;
   32975: result <= 12'b111111101000;
   32976: result <= 12'b111111101000;
   32977: result <= 12'b111111101001;
   32978: result <= 12'b111111101001;
   32979: result <= 12'b111111101001;
   32980: result <= 12'b111111101001;
   32981: result <= 12'b111111101001;
   32982: result <= 12'b111111101010;
   32983: result <= 12'b111111101010;
   32984: result <= 12'b111111101010;
   32985: result <= 12'b111111101010;
   32986: result <= 12'b111111101010;
   32987: result <= 12'b111111101010;
   32988: result <= 12'b111111101011;
   32989: result <= 12'b111111101011;
   32990: result <= 12'b111111101011;
   32991: result <= 12'b111111101011;
   32992: result <= 12'b111111101011;
   32993: result <= 12'b111111101100;
   32994: result <= 12'b111111101100;
   32995: result <= 12'b111111101100;
   32996: result <= 12'b111111101100;
   32997: result <= 12'b111111101100;
   32998: result <= 12'b111111101101;
   32999: result <= 12'b111111101101;
   33000: result <= 12'b111111101101;
   33001: result <= 12'b111111101101;
   33002: result <= 12'b111111101101;
   33003: result <= 12'b111111101110;
   33004: result <= 12'b111111101110;
   33005: result <= 12'b111111101110;
   33006: result <= 12'b111111101110;
   33007: result <= 12'b111111101110;
   33008: result <= 12'b111111101111;
   33009: result <= 12'b111111101111;
   33010: result <= 12'b111111101111;
   33011: result <= 12'b111111101111;
   33012: result <= 12'b111111101111;
   33013: result <= 12'b111111110000;
   33014: result <= 12'b111111110000;
   33015: result <= 12'b111111110000;
   33016: result <= 12'b111111110000;
   33017: result <= 12'b111111110000;
   33018: result <= 12'b111111110001;
   33019: result <= 12'b111111110001;
   33020: result <= 12'b111111110001;
   33021: result <= 12'b111111110001;
   33022: result <= 12'b111111110001;
   33023: result <= 12'b111111110010;
   33024: result <= 12'b111111110010;
   33025: result <= 12'b111111110010;
   33026: result <= 12'b111111110010;
   33027: result <= 12'b111111110010;
   33028: result <= 12'b111111110011;
   33029: result <= 12'b111111110011;
   33030: result <= 12'b111111110011;
   33031: result <= 12'b111111110011;
   33032: result <= 12'b111111110011;
   33033: result <= 12'b111111110100;
   33034: result <= 12'b111111110100;
   33035: result <= 12'b111111110100;
   33036: result <= 12'b111111110100;
   33037: result <= 12'b111111110100;
   33038: result <= 12'b111111110101;
   33039: result <= 12'b111111110101;
   33040: result <= 12'b111111110101;
   33041: result <= 12'b111111110101;
   33042: result <= 12'b111111110101;
   33043: result <= 12'b111111110101;
   33044: result <= 12'b111111110110;
   33045: result <= 12'b111111110110;
   33046: result <= 12'b111111110110;
   33047: result <= 12'b111111110110;
   33048: result <= 12'b111111110110;
   33049: result <= 12'b111111110111;
   33050: result <= 12'b111111110111;
   33051: result <= 12'b111111110111;
   33052: result <= 12'b111111110111;
   33053: result <= 12'b111111110111;
   33054: result <= 12'b111111111000;
   33055: result <= 12'b111111111000;
   33056: result <= 12'b111111111000;
   33057: result <= 12'b111111111000;
   33058: result <= 12'b111111111000;
   33059: result <= 12'b111111111001;
   33060: result <= 12'b111111111001;
   33061: result <= 12'b111111111001;
   33062: result <= 12'b111111111001;
   33063: result <= 12'b111111111001;
   33064: result <= 12'b111111111010;
   33065: result <= 12'b111111111010;
   33066: result <= 12'b111111111010;
   33067: result <= 12'b111111111010;
   33068: result <= 12'b111111111010;
   33069: result <= 12'b111111111011;
   33070: result <= 12'b111111111011;
   33071: result <= 12'b111111111011;
   33072: result <= 12'b111111111011;
   33073: result <= 12'b111111111011;
   33074: result <= 12'b111111111100;
   33075: result <= 12'b111111111100;
   33076: result <= 12'b111111111100;
   33077: result <= 12'b111111111100;
   33078: result <= 12'b111111111100;
   33079: result <= 12'b111111111101;
   33080: result <= 12'b111111111101;
   33081: result <= 12'b111111111101;
   33082: result <= 12'b111111111101;
   33083: result <= 12'b111111111101;
   33084: result <= 12'b111111111110;
   33085: result <= 12'b111111111110;
   33086: result <= 12'b111111111110;
   33087: result <= 12'b111111111110;
   33088: result <= 12'b111111111110;
   33089: result <= 12'b111111111111;
   33090: result <= 12'b111111111111;
   33091: result <= 12'b111111111111;
   33092: result <= 12'b111111111111;
   33093: result <= 12'b111111111111;
   33094: result <= 12'b111111111111;
   33095: result <= 12'b111111000000;
   33096: result <= 12'b111111000000;
   33097: result <= 12'b111111000000;
   33098: result <= 12'b111111000000;
   33099: result <= 12'b111111000000;
   33100: result <= 12'b111111000001;
   33101: result <= 12'b111111000001;
   33102: result <= 12'b111111000001;
   33103: result <= 12'b111111000001;
   33104: result <= 12'b111111000001;
   33105: result <= 12'b111111000010;
   33106: result <= 12'b111111000010;
   33107: result <= 12'b111111000010;
   33108: result <= 12'b111111000010;
   33109: result <= 12'b111111000010;
   33110: result <= 12'b111111000011;
   33111: result <= 12'b111111000011;
   33112: result <= 12'b111111000011;
   33113: result <= 12'b111111000011;
   33114: result <= 12'b111111000011;
   33115: result <= 12'b111111000100;
   33116: result <= 12'b111111000100;
   33117: result <= 12'b111111000100;
   33118: result <= 12'b111111000100;
   33119: result <= 12'b111111000100;
   33120: result <= 12'b111111000101;
   33121: result <= 12'b111111000101;
   33122: result <= 12'b111111000101;
   33123: result <= 12'b111111000101;
   33124: result <= 12'b111111000101;
   33125: result <= 12'b111111000110;
   33126: result <= 12'b111111000110;
   33127: result <= 12'b111111000110;
   33128: result <= 12'b111111000110;
   33129: result <= 12'b111111000110;
   33130: result <= 12'b111111000111;
   33131: result <= 12'b111111000111;
   33132: result <= 12'b111111000111;
   33133: result <= 12'b111111000111;
   33134: result <= 12'b111111000111;
   33135: result <= 12'b111111001000;
   33136: result <= 12'b111111001000;
   33137: result <= 12'b111111001000;
   33138: result <= 12'b111111001000;
   33139: result <= 12'b111111001000;
   33140: result <= 12'b111111001001;
   33141: result <= 12'b111111001001;
   33142: result <= 12'b111111001001;
   33143: result <= 12'b111111001001;
   33144: result <= 12'b111111001001;
   33145: result <= 12'b111111001010;
   33146: result <= 12'b111111001010;
   33147: result <= 12'b111111001010;
   33148: result <= 12'b111111001010;
   33149: result <= 12'b111111001010;
   33150: result <= 12'b111111001010;
   33151: result <= 12'b111111001011;
   33152: result <= 12'b111111001011;
   33153: result <= 12'b111111001011;
   33154: result <= 12'b111111001011;
   33155: result <= 12'b111111001011;
   33156: result <= 12'b111111001100;
   33157: result <= 12'b111111001100;
   33158: result <= 12'b111111001100;
   33159: result <= 12'b111111001100;
   33160: result <= 12'b111111001100;
   33161: result <= 12'b111111001101;
   33162: result <= 12'b111111001101;
   33163: result <= 12'b111111001101;
   33164: result <= 12'b111111001101;
   33165: result <= 12'b111111001101;
   33166: result <= 12'b111111001110;
   33167: result <= 12'b111111001110;
   33168: result <= 12'b111111001110;
   33169: result <= 12'b111111001110;
   33170: result <= 12'b111111001110;
   33171: result <= 12'b111111001111;
   33172: result <= 12'b111111001111;
   33173: result <= 12'b111111001111;
   33174: result <= 12'b111111001111;
   33175: result <= 12'b111111001111;
   33176: result <= 12'b111111010000;
   33177: result <= 12'b111111010000;
   33178: result <= 12'b111111010000;
   33179: result <= 12'b111111010000;
   33180: result <= 12'b111111010000;
   33181: result <= 12'b111111010001;
   33182: result <= 12'b111111010001;
   33183: result <= 12'b111111010001;
   33184: result <= 12'b111111010001;
   33185: result <= 12'b111111010001;
   33186: result <= 12'b111111010010;
   33187: result <= 12'b111111010010;
   33188: result <= 12'b111111010010;
   33189: result <= 12'b111111010010;
   33190: result <= 12'b111111010010;
   33191: result <= 12'b111111010011;
   33192: result <= 12'b111111010011;
   33193: result <= 12'b111111010011;
   33194: result <= 12'b111111010011;
   33195: result <= 12'b111111010011;
   33196: result <= 12'b111111010100;
   33197: result <= 12'b111111010100;
   33198: result <= 12'b111111010100;
   33199: result <= 12'b111111010100;
   33200: result <= 12'b111111010100;
   33201: result <= 12'b111111010100;
   33202: result <= 12'b111111010101;
   33203: result <= 12'b111111010101;
   33204: result <= 12'b111111010101;
   33205: result <= 12'b111111010101;
   33206: result <= 12'b111111010101;
   33207: result <= 12'b111111010110;
   33208: result <= 12'b111111010110;
   33209: result <= 12'b111111010110;
   33210: result <= 12'b111111010110;
   33211: result <= 12'b111111010110;
   33212: result <= 12'b111111010111;
   33213: result <= 12'b111111010111;
   33214: result <= 12'b111111010111;
   33215: result <= 12'b111111010111;
   33216: result <= 12'b111111010111;
   33217: result <= 12'b111111011000;
   33218: result <= 12'b111111011000;
   33219: result <= 12'b111111011000;
   33220: result <= 12'b111111011000;
   33221: result <= 12'b111111011000;
   33222: result <= 12'b111111011001;
   33223: result <= 12'b111111011001;
   33224: result <= 12'b111111011001;
   33225: result <= 12'b111111011001;
   33226: result <= 12'b111111011001;
   33227: result <= 12'b111111011010;
   33228: result <= 12'b111111011010;
   33229: result <= 12'b111111011010;
   33230: result <= 12'b111111011010;
   33231: result <= 12'b111111011010;
   33232: result <= 12'b111111011011;
   33233: result <= 12'b111111011011;
   33234: result <= 12'b111111011011;
   33235: result <= 12'b111111011011;
   33236: result <= 12'b111111011011;
   33237: result <= 12'b111111011100;
   33238: result <= 12'b111111011100;
   33239: result <= 12'b111111011100;
   33240: result <= 12'b111111011100;
   33241: result <= 12'b111111011100;
   33242: result <= 12'b111111011101;
   33243: result <= 12'b111111011101;
   33244: result <= 12'b111111011101;
   33245: result <= 12'b111111011101;
   33246: result <= 12'b111111011101;
   33247: result <= 12'b111111011110;
   33248: result <= 12'b111111011110;
   33249: result <= 12'b111111011110;
   33250: result <= 12'b111111011110;
   33251: result <= 12'b111111011110;
   33252: result <= 12'b111111011110;
   33253: result <= 12'b111111011111;
   33254: result <= 12'b111111011111;
   33255: result <= 12'b111111011111;
   33256: result <= 12'b111111011111;
   33257: result <= 12'b111111011111;
   33258: result <= 12'b111111100000;
   33259: result <= 12'b111111100000;
   33260: result <= 12'b111111100000;
   33261: result <= 12'b111111100000;
   33262: result <= 12'b111111100000;
   33263: result <= 12'b111111100001;
   33264: result <= 12'b111111100001;
   33265: result <= 12'b111111100001;
   33266: result <= 12'b111111100001;
   33267: result <= 12'b111111100001;
   33268: result <= 12'b111111100010;
   33269: result <= 12'b111111100010;
   33270: result <= 12'b111111100010;
   33271: result <= 12'b111111100010;
   33272: result <= 12'b111111100010;
   33273: result <= 12'b111111100011;
   33274: result <= 12'b111111100011;
   33275: result <= 12'b111111100011;
   33276: result <= 12'b111111100011;
   33277: result <= 12'b111111100011;
   33278: result <= 12'b111111100100;
   33279: result <= 12'b111111100100;
   33280: result <= 12'b111111100100;
   33281: result <= 12'b111111100100;
   33282: result <= 12'b111111100100;
   33283: result <= 12'b111111100101;
   33284: result <= 12'b111111100101;
   33285: result <= 12'b111111100101;
   33286: result <= 12'b111111100101;
   33287: result <= 12'b111111100101;
   33288: result <= 12'b111111100110;
   33289: result <= 12'b111111100110;
   33290: result <= 12'b111111100110;
   33291: result <= 12'b111111100110;
   33292: result <= 12'b111111100110;
   33293: result <= 12'b111111100111;
   33294: result <= 12'b111111100111;
   33295: result <= 12'b111111100111;
   33296: result <= 12'b111111100111;
   33297: result <= 12'b111111100111;
   33298: result <= 12'b111111101000;
   33299: result <= 12'b111111101000;
   33300: result <= 12'b111111101000;
   33301: result <= 12'b111111101000;
   33302: result <= 12'b111111101000;
   33303: result <= 12'b111111101001;
   33304: result <= 12'b111111101001;
   33305: result <= 12'b111111101001;
   33306: result <= 12'b111111101001;
   33307: result <= 12'b111111101001;
   33308: result <= 12'b111111101001;
   33309: result <= 12'b111111101010;
   33310: result <= 12'b111111101010;
   33311: result <= 12'b111111101010;
   33312: result <= 12'b111111101010;
   33313: result <= 12'b111111101010;
   33314: result <= 12'b111111101011;
   33315: result <= 12'b111111101011;
   33316: result <= 12'b111111101011;
   33317: result <= 12'b111111101011;
   33318: result <= 12'b111111101011;
   33319: result <= 12'b111111101100;
   33320: result <= 12'b111111101100;
   33321: result <= 12'b111111101100;
   33322: result <= 12'b111111101100;
   33323: result <= 12'b111111101100;
   33324: result <= 12'b111111101101;
   33325: result <= 12'b111111101101;
   33326: result <= 12'b111111101101;
   33327: result <= 12'b111111101101;
   33328: result <= 12'b111111101101;
   33329: result <= 12'b111111101110;
   33330: result <= 12'b111111101110;
   33331: result <= 12'b111111101110;
   33332: result <= 12'b111111101110;
   33333: result <= 12'b111111101110;
   33334: result <= 12'b111111101111;
   33335: result <= 12'b111111101111;
   33336: result <= 12'b111111101111;
   33337: result <= 12'b111111101111;
   33338: result <= 12'b111111101111;
   33339: result <= 12'b111111110000;
   33340: result <= 12'b111111110000;
   33341: result <= 12'b111111110000;
   33342: result <= 12'b111111110000;
   33343: result <= 12'b111111110000;
   33344: result <= 12'b111111110001;
   33345: result <= 12'b111111110001;
   33346: result <= 12'b111111110001;
   33347: result <= 12'b111111110001;
   33348: result <= 12'b111111110001;
   33349: result <= 12'b111111110010;
   33350: result <= 12'b111111110010;
   33351: result <= 12'b111111110010;
   33352: result <= 12'b111111110010;
   33353: result <= 12'b111111110010;
   33354: result <= 12'b111111110011;
   33355: result <= 12'b111111110011;
   33356: result <= 12'b111111110011;
   33357: result <= 12'b111111110011;
   33358: result <= 12'b111111110011;
   33359: result <= 12'b111111110011;
   33360: result <= 12'b111111110100;
   33361: result <= 12'b111111110100;
   33362: result <= 12'b111111110100;
   33363: result <= 12'b111111110100;
   33364: result <= 12'b111111110100;
   33365: result <= 12'b111111110101;
   33366: result <= 12'b111111110101;
   33367: result <= 12'b111111110101;
   33368: result <= 12'b111111110101;
   33369: result <= 12'b111111110101;
   33370: result <= 12'b111111110110;
   33371: result <= 12'b111111110110;
   33372: result <= 12'b111111110110;
   33373: result <= 12'b111111110110;
   33374: result <= 12'b111111110110;
   33375: result <= 12'b111111110111;
   33376: result <= 12'b111111110111;
   33377: result <= 12'b111111110111;
   33378: result <= 12'b111111110111;
   33379: result <= 12'b111111110111;
   33380: result <= 12'b111111111000;
   33381: result <= 12'b111111111000;
   33382: result <= 12'b111111111000;
   33383: result <= 12'b111111111000;
   33384: result <= 12'b111111111000;
   33385: result <= 12'b111111111001;
   33386: result <= 12'b111111111001;
   33387: result <= 12'b111111111001;
   33388: result <= 12'b111111111001;
   33389: result <= 12'b111111111001;
   33390: result <= 12'b111111111010;
   33391: result <= 12'b111111111010;
   33392: result <= 12'b111111111010;
   33393: result <= 12'b111111111010;
   33394: result <= 12'b111111111010;
   33395: result <= 12'b111111111011;
   33396: result <= 12'b111111111011;
   33397: result <= 12'b111111111011;
   33398: result <= 12'b111111111011;
   33399: result <= 12'b111111111011;
   33400: result <= 12'b111111111100;
   33401: result <= 12'b111111111100;
   33402: result <= 12'b111111111100;
   33403: result <= 12'b111111111100;
   33404: result <= 12'b111111111100;
   33405: result <= 12'b111111111100;
   33406: result <= 12'b111111111101;
   33407: result <= 12'b111111111101;
   33408: result <= 12'b111111111101;
   33409: result <= 12'b111111111101;
   33410: result <= 12'b111111111101;
   33411: result <= 12'b111111111110;
   33412: result <= 12'b111111111110;
   33413: result <= 12'b111111111110;
   33414: result <= 12'b111111111110;
   33415: result <= 12'b111111111110;
   33416: result <= 12'b111111111111;
   33417: result <= 12'b111111111111;
   33418: result <= 12'b111111111111;
   33419: result <= 12'b111111111111;
   33420: result <= 12'b111111111111;
   33421: result <= 12'b111110000000;
   33422: result <= 12'b111110000000;
   33423: result <= 12'b111110000000;
   33424: result <= 12'b111110000000;
   33425: result <= 12'b111110000000;
   33426: result <= 12'b111110000001;
   33427: result <= 12'b111110000001;
   33428: result <= 12'b111110000001;
   33429: result <= 12'b111110000001;
   33430: result <= 12'b111110000001;
   33431: result <= 12'b111110000010;
   33432: result <= 12'b111110000010;
   33433: result <= 12'b111110000010;
   33434: result <= 12'b111110000010;
   33435: result <= 12'b111110000010;
   33436: result <= 12'b111110000011;
   33437: result <= 12'b111110000011;
   33438: result <= 12'b111110000011;
   33439: result <= 12'b111110000011;
   33440: result <= 12'b111110000011;
   33441: result <= 12'b111110000100;
   33442: result <= 12'b111110000100;
   33443: result <= 12'b111110000100;
   33444: result <= 12'b111110000100;
   33445: result <= 12'b111110000100;
   33446: result <= 12'b111110000101;
   33447: result <= 12'b111110000101;
   33448: result <= 12'b111110000101;
   33449: result <= 12'b111110000101;
   33450: result <= 12'b111110000101;
   33451: result <= 12'b111110000110;
   33452: result <= 12'b111110000110;
   33453: result <= 12'b111110000110;
   33454: result <= 12'b111110000110;
   33455: result <= 12'b111110000110;
   33456: result <= 12'b111110000110;
   33457: result <= 12'b111110000111;
   33458: result <= 12'b111110000111;
   33459: result <= 12'b111110000111;
   33460: result <= 12'b111110000111;
   33461: result <= 12'b111110000111;
   33462: result <= 12'b111110001000;
   33463: result <= 12'b111110001000;
   33464: result <= 12'b111110001000;
   33465: result <= 12'b111110001000;
   33466: result <= 12'b111110001000;
   33467: result <= 12'b111110001001;
   33468: result <= 12'b111110001001;
   33469: result <= 12'b111110001001;
   33470: result <= 12'b111110001001;
   33471: result <= 12'b111110001001;
   33472: result <= 12'b111110001010;
   33473: result <= 12'b111110001010;
   33474: result <= 12'b111110001010;
   33475: result <= 12'b111110001010;
   33476: result <= 12'b111110001010;
   33477: result <= 12'b111110001011;
   33478: result <= 12'b111110001011;
   33479: result <= 12'b111110001011;
   33480: result <= 12'b111110001011;
   33481: result <= 12'b111110001011;
   33482: result <= 12'b111110001100;
   33483: result <= 12'b111110001100;
   33484: result <= 12'b111110001100;
   33485: result <= 12'b111110001100;
   33486: result <= 12'b111110001100;
   33487: result <= 12'b111110001101;
   33488: result <= 12'b111110001101;
   33489: result <= 12'b111110001101;
   33490: result <= 12'b111110001101;
   33491: result <= 12'b111110001101;
   33492: result <= 12'b111110001110;
   33493: result <= 12'b111110001110;
   33494: result <= 12'b111110001110;
   33495: result <= 12'b111110001110;
   33496: result <= 12'b111110001110;
   33497: result <= 12'b111110001111;
   33498: result <= 12'b111110001111;
   33499: result <= 12'b111110001111;
   33500: result <= 12'b111110001111;
   33501: result <= 12'b111110001111;
   33502: result <= 12'b111110010000;
   33503: result <= 12'b111110010000;
   33504: result <= 12'b111110010000;
   33505: result <= 12'b111110010000;
   33506: result <= 12'b111110010000;
   33507: result <= 12'b111110010000;
   33508: result <= 12'b111110010001;
   33509: result <= 12'b111110010001;
   33510: result <= 12'b111110010001;
   33511: result <= 12'b111110010001;
   33512: result <= 12'b111110010001;
   33513: result <= 12'b111110010010;
   33514: result <= 12'b111110010010;
   33515: result <= 12'b111110010010;
   33516: result <= 12'b111110010010;
   33517: result <= 12'b111110010010;
   33518: result <= 12'b111110010011;
   33519: result <= 12'b111110010011;
   33520: result <= 12'b111110010011;
   33521: result <= 12'b111110010011;
   33522: result <= 12'b111110010011;
   33523: result <= 12'b111110010100;
   33524: result <= 12'b111110010100;
   33525: result <= 12'b111110010100;
   33526: result <= 12'b111110010100;
   33527: result <= 12'b111110010100;
   33528: result <= 12'b111110010101;
   33529: result <= 12'b111110010101;
   33530: result <= 12'b111110010101;
   33531: result <= 12'b111110010101;
   33532: result <= 12'b111110010101;
   33533: result <= 12'b111110010110;
   33534: result <= 12'b111110010110;
   33535: result <= 12'b111110010110;
   33536: result <= 12'b111110010110;
   33537: result <= 12'b111110010110;
   33538: result <= 12'b111110010111;
   33539: result <= 12'b111110010111;
   33540: result <= 12'b111110010111;
   33541: result <= 12'b111110010111;
   33542: result <= 12'b111110010111;
   33543: result <= 12'b111110011000;
   33544: result <= 12'b111110011000;
   33545: result <= 12'b111110011000;
   33546: result <= 12'b111110011000;
   33547: result <= 12'b111110011000;
   33548: result <= 12'b111110011001;
   33549: result <= 12'b111110011001;
   33550: result <= 12'b111110011001;
   33551: result <= 12'b111110011001;
   33552: result <= 12'b111110011001;
   33553: result <= 12'b111110011001;
   33554: result <= 12'b111110011010;
   33555: result <= 12'b111110011010;
   33556: result <= 12'b111110011010;
   33557: result <= 12'b111110011010;
   33558: result <= 12'b111110011010;
   33559: result <= 12'b111110011011;
   33560: result <= 12'b111110011011;
   33561: result <= 12'b111110011011;
   33562: result <= 12'b111110011011;
   33563: result <= 12'b111110011011;
   33564: result <= 12'b111110011100;
   33565: result <= 12'b111110011100;
   33566: result <= 12'b111110011100;
   33567: result <= 12'b111110011100;
   33568: result <= 12'b111110011100;
   33569: result <= 12'b111110011101;
   33570: result <= 12'b111110011101;
   33571: result <= 12'b111110011101;
   33572: result <= 12'b111110011101;
   33573: result <= 12'b111110011101;
   33574: result <= 12'b111110011110;
   33575: result <= 12'b111110011110;
   33576: result <= 12'b111110011110;
   33577: result <= 12'b111110011110;
   33578: result <= 12'b111110011110;
   33579: result <= 12'b111110011111;
   33580: result <= 12'b111110011111;
   33581: result <= 12'b111110011111;
   33582: result <= 12'b111110011111;
   33583: result <= 12'b111110011111;
   33584: result <= 12'b111110100000;
   33585: result <= 12'b111110100000;
   33586: result <= 12'b111110100000;
   33587: result <= 12'b111110100000;
   33588: result <= 12'b111110100000;
   33589: result <= 12'b111110100001;
   33590: result <= 12'b111110100001;
   33591: result <= 12'b111110100001;
   33592: result <= 12'b111110100001;
   33593: result <= 12'b111110100001;
   33594: result <= 12'b111110100010;
   33595: result <= 12'b111110100010;
   33596: result <= 12'b111110100010;
   33597: result <= 12'b111110100010;
   33598: result <= 12'b111110100010;
   33599: result <= 12'b111110100010;
   33600: result <= 12'b111110100011;
   33601: result <= 12'b111110100011;
   33602: result <= 12'b111110100011;
   33603: result <= 12'b111110100011;
   33604: result <= 12'b111110100011;
   33605: result <= 12'b111110100100;
   33606: result <= 12'b111110100100;
   33607: result <= 12'b111110100100;
   33608: result <= 12'b111110100100;
   33609: result <= 12'b111110100100;
   33610: result <= 12'b111110100101;
   33611: result <= 12'b111110100101;
   33612: result <= 12'b111110100101;
   33613: result <= 12'b111110100101;
   33614: result <= 12'b111110100101;
   33615: result <= 12'b111110100110;
   33616: result <= 12'b111110100110;
   33617: result <= 12'b111110100110;
   33618: result <= 12'b111110100110;
   33619: result <= 12'b111110100110;
   33620: result <= 12'b111110100111;
   33621: result <= 12'b111110100111;
   33622: result <= 12'b111110100111;
   33623: result <= 12'b111110100111;
   33624: result <= 12'b111110100111;
   33625: result <= 12'b111110101000;
   33626: result <= 12'b111110101000;
   33627: result <= 12'b111110101000;
   33628: result <= 12'b111110101000;
   33629: result <= 12'b111110101000;
   33630: result <= 12'b111110101001;
   33631: result <= 12'b111110101001;
   33632: result <= 12'b111110101001;
   33633: result <= 12'b111110101001;
   33634: result <= 12'b111110101001;
   33635: result <= 12'b111110101010;
   33636: result <= 12'b111110101010;
   33637: result <= 12'b111110101010;
   33638: result <= 12'b111110101010;
   33639: result <= 12'b111110101010;
   33640: result <= 12'b111110101011;
   33641: result <= 12'b111110101011;
   33642: result <= 12'b111110101011;
   33643: result <= 12'b111110101011;
   33644: result <= 12'b111110101011;
   33645: result <= 12'b111110101011;
   33646: result <= 12'b111110101100;
   33647: result <= 12'b111110101100;
   33648: result <= 12'b111110101100;
   33649: result <= 12'b111110101100;
   33650: result <= 12'b111110101100;
   33651: result <= 12'b111110101101;
   33652: result <= 12'b111110101101;
   33653: result <= 12'b111110101101;
   33654: result <= 12'b111110101101;
   33655: result <= 12'b111110101101;
   33656: result <= 12'b111110101110;
   33657: result <= 12'b111110101110;
   33658: result <= 12'b111110101110;
   33659: result <= 12'b111110101110;
   33660: result <= 12'b111110101110;
   33661: result <= 12'b111110101111;
   33662: result <= 12'b111110101111;
   33663: result <= 12'b111110101111;
   33664: result <= 12'b111110101111;
   33665: result <= 12'b111110101111;
   33666: result <= 12'b111110110000;
   33667: result <= 12'b111110110000;
   33668: result <= 12'b111110110000;
   33669: result <= 12'b111110110000;
   33670: result <= 12'b111110110000;
   33671: result <= 12'b111110110001;
   33672: result <= 12'b111110110001;
   33673: result <= 12'b111110110001;
   33674: result <= 12'b111110110001;
   33675: result <= 12'b111110110001;
   33676: result <= 12'b111110110010;
   33677: result <= 12'b111110110010;
   33678: result <= 12'b111110110010;
   33679: result <= 12'b111110110010;
   33680: result <= 12'b111110110010;
   33681: result <= 12'b111110110011;
   33682: result <= 12'b111110110011;
   33683: result <= 12'b111110110011;
   33684: result <= 12'b111110110011;
   33685: result <= 12'b111110110011;
   33686: result <= 12'b111110110100;
   33687: result <= 12'b111110110100;
   33688: result <= 12'b111110110100;
   33689: result <= 12'b111110110100;
   33690: result <= 12'b111110110100;
   33691: result <= 12'b111110110100;
   33692: result <= 12'b111110110101;
   33693: result <= 12'b111110110101;
   33694: result <= 12'b111110110101;
   33695: result <= 12'b111110110101;
   33696: result <= 12'b111110110101;
   33697: result <= 12'b111110110110;
   33698: result <= 12'b111110110110;
   33699: result <= 12'b111110110110;
   33700: result <= 12'b111110110110;
   33701: result <= 12'b111110110110;
   33702: result <= 12'b111110110111;
   33703: result <= 12'b111110110111;
   33704: result <= 12'b111110110111;
   33705: result <= 12'b111110110111;
   33706: result <= 12'b111110110111;
   33707: result <= 12'b111110111000;
   33708: result <= 12'b111110111000;
   33709: result <= 12'b111110111000;
   33710: result <= 12'b111110111000;
   33711: result <= 12'b111110111000;
   33712: result <= 12'b111110111001;
   33713: result <= 12'b111110111001;
   33714: result <= 12'b111110111001;
   33715: result <= 12'b111110111001;
   33716: result <= 12'b111110111001;
   33717: result <= 12'b111110111010;
   33718: result <= 12'b111110111010;
   33719: result <= 12'b111110111010;
   33720: result <= 12'b111110111010;
   33721: result <= 12'b111110111010;
   33722: result <= 12'b111110111011;
   33723: result <= 12'b111110111011;
   33724: result <= 12'b111110111011;
   33725: result <= 12'b111110111011;
   33726: result <= 12'b111110111011;
   33727: result <= 12'b111110111100;
   33728: result <= 12'b111110111100;
   33729: result <= 12'b111110111100;
   33730: result <= 12'b111110111100;
   33731: result <= 12'b111110111100;
   33732: result <= 12'b111110111101;
   33733: result <= 12'b111110111101;
   33734: result <= 12'b111110111101;
   33735: result <= 12'b111110111101;
   33736: result <= 12'b111110111101;
   33737: result <= 12'b111110111101;
   33738: result <= 12'b111110111110;
   33739: result <= 12'b111110111110;
   33740: result <= 12'b111110111110;
   33741: result <= 12'b111110111110;
   33742: result <= 12'b111110111110;
   33743: result <= 12'b111110111111;
   33744: result <= 12'b111110111111;
   33745: result <= 12'b111110111111;
   33746: result <= 12'b111110111111;
   33747: result <= 12'b111110111111;
   33748: result <= 12'b111111000000;
   33749: result <= 12'b111111000000;
   33750: result <= 12'b111111000000;
   33751: result <= 12'b111111000000;
   33752: result <= 12'b111111000000;
   33753: result <= 12'b111111000001;
   33754: result <= 12'b111111000001;
   33755: result <= 12'b111111000001;
   33756: result <= 12'b111111000001;
   33757: result <= 12'b111111000001;
   33758: result <= 12'b111111000010;
   33759: result <= 12'b111111000010;
   33760: result <= 12'b111111000010;
   33761: result <= 12'b111111000010;
   33762: result <= 12'b111111000010;
   33763: result <= 12'b111111000011;
   33764: result <= 12'b111111000011;
   33765: result <= 12'b111111000011;
   33766: result <= 12'b111111000011;
   33767: result <= 12'b111111000011;
   33768: result <= 12'b111111000100;
   33769: result <= 12'b111111000100;
   33770: result <= 12'b111111000100;
   33771: result <= 12'b111111000100;
   33772: result <= 12'b111111000100;
   33773: result <= 12'b111111000101;
   33774: result <= 12'b111111000101;
   33775: result <= 12'b111111000101;
   33776: result <= 12'b111111000101;
   33777: result <= 12'b111111000101;
   33778: result <= 12'b111111000110;
   33779: result <= 12'b111111000110;
   33780: result <= 12'b111111000110;
   33781: result <= 12'b111111000110;
   33782: result <= 12'b111111000110;
   33783: result <= 12'b111111000110;
   33784: result <= 12'b111111000111;
   33785: result <= 12'b111111000111;
   33786: result <= 12'b111111000111;
   33787: result <= 12'b111111000111;
   33788: result <= 12'b111111000111;
   33789: result <= 12'b111111001000;
   33790: result <= 12'b111111001000;
   33791: result <= 12'b111111001000;
   33792: result <= 12'b111111001000;
   33793: result <= 12'b111111001000;
   33794: result <= 12'b111111001001;
   33795: result <= 12'b111111001001;
   33796: result <= 12'b111111001001;
   33797: result <= 12'b111111001001;
   33798: result <= 12'b111111001001;
   33799: result <= 12'b111111001010;
   33800: result <= 12'b111111001010;
   33801: result <= 12'b111111001010;
   33802: result <= 12'b111111001010;
   33803: result <= 12'b111111001010;
   33804: result <= 12'b111111001011;
   33805: result <= 12'b111111001011;
   33806: result <= 12'b111111001011;
   33807: result <= 12'b111111001011;
   33808: result <= 12'b111111001011;
   33809: result <= 12'b111111001100;
   33810: result <= 12'b111111001100;
   33811: result <= 12'b111111001100;
   33812: result <= 12'b111111001100;
   33813: result <= 12'b111111001100;
   33814: result <= 12'b111111001101;
   33815: result <= 12'b111111001101;
   33816: result <= 12'b111111001101;
   33817: result <= 12'b111111001101;
   33818: result <= 12'b111111001101;
   33819: result <= 12'b111111001110;
   33820: result <= 12'b111111001110;
   33821: result <= 12'b111111001110;
   33822: result <= 12'b111111001110;
   33823: result <= 12'b111111001110;
   33824: result <= 12'b111111001110;
   33825: result <= 12'b111111001111;
   33826: result <= 12'b111111001111;
   33827: result <= 12'b111111001111;
   33828: result <= 12'b111111001111;
   33829: result <= 12'b111111001111;
   33830: result <= 12'b111111010000;
   33831: result <= 12'b111111010000;
   33832: result <= 12'b111111010000;
   33833: result <= 12'b111111010000;
   33834: result <= 12'b111111010000;
   33835: result <= 12'b111111010001;
   33836: result <= 12'b111111010001;
   33837: result <= 12'b111111010001;
   33838: result <= 12'b111111010001;
   33839: result <= 12'b111111010001;
   33840: result <= 12'b111111010010;
   33841: result <= 12'b111111010010;
   33842: result <= 12'b111111010010;
   33843: result <= 12'b111111010010;
   33844: result <= 12'b111111010010;
   33845: result <= 12'b111111010011;
   33846: result <= 12'b111111010011;
   33847: result <= 12'b111111010011;
   33848: result <= 12'b111111010011;
   33849: result <= 12'b111111010011;
   33850: result <= 12'b111111010100;
   33851: result <= 12'b111111010100;
   33852: result <= 12'b111111010100;
   33853: result <= 12'b111111010100;
   33854: result <= 12'b111111010100;
   33855: result <= 12'b111111010101;
   33856: result <= 12'b111111010101;
   33857: result <= 12'b111111010101;
   33858: result <= 12'b111111010101;
   33859: result <= 12'b111111010101;
   33860: result <= 12'b111111010110;
   33861: result <= 12'b111111010110;
   33862: result <= 12'b111111010110;
   33863: result <= 12'b111111010110;
   33864: result <= 12'b111111010110;
   33865: result <= 12'b111111010110;
   33866: result <= 12'b111111010111;
   33867: result <= 12'b111111010111;
   33868: result <= 12'b111111010111;
   33869: result <= 12'b111111010111;
   33870: result <= 12'b111111010111;
   33871: result <= 12'b111111011000;
   33872: result <= 12'b111111011000;
   33873: result <= 12'b111111011000;
   33874: result <= 12'b111111011000;
   33875: result <= 12'b111111011000;
   33876: result <= 12'b111111011001;
   33877: result <= 12'b111111011001;
   33878: result <= 12'b111111011001;
   33879: result <= 12'b111111011001;
   33880: result <= 12'b111111011001;
   33881: result <= 12'b111111011010;
   33882: result <= 12'b111111011010;
   33883: result <= 12'b111111011010;
   33884: result <= 12'b111111011010;
   33885: result <= 12'b111111011010;
   33886: result <= 12'b111111011011;
   33887: result <= 12'b111111011011;
   33888: result <= 12'b111111011011;
   33889: result <= 12'b111111011011;
   33890: result <= 12'b111111011011;
   33891: result <= 12'b111111011100;
   33892: result <= 12'b111111011100;
   33893: result <= 12'b111111011100;
   33894: result <= 12'b111111011100;
   33895: result <= 12'b111111011100;
   33896: result <= 12'b111111011101;
   33897: result <= 12'b111111011101;
   33898: result <= 12'b111111011101;
   33899: result <= 12'b111111011101;
   33900: result <= 12'b111111011101;
   33901: result <= 12'b111111011110;
   33902: result <= 12'b111111011110;
   33903: result <= 12'b111111011110;
   33904: result <= 12'b111111011110;
   33905: result <= 12'b111111011110;
   33906: result <= 12'b111111011111;
   33907: result <= 12'b111111011111;
   33908: result <= 12'b111111011111;
   33909: result <= 12'b111111011111;
   33910: result <= 12'b111111011111;
   33911: result <= 12'b111111011111;
   33912: result <= 12'b111111100000;
   33913: result <= 12'b111111100000;
   33914: result <= 12'b111111100000;
   33915: result <= 12'b111111100000;
   33916: result <= 12'b111111100000;
   33917: result <= 12'b111111100001;
   33918: result <= 12'b111111100001;
   33919: result <= 12'b111111100001;
   33920: result <= 12'b111111100001;
   33921: result <= 12'b111111100001;
   33922: result <= 12'b111111100010;
   33923: result <= 12'b111111100010;
   33924: result <= 12'b111111100010;
   33925: result <= 12'b111111100010;
   33926: result <= 12'b111111100010;
   33927: result <= 12'b111111100011;
   33928: result <= 12'b111111100011;
   33929: result <= 12'b111111100011;
   33930: result <= 12'b111111100011;
   33931: result <= 12'b111111100011;
   33932: result <= 12'b111111100100;
   33933: result <= 12'b111111100100;
   33934: result <= 12'b111111100100;
   33935: result <= 12'b111111100100;
   33936: result <= 12'b111111100100;
   33937: result <= 12'b111111100101;
   33938: result <= 12'b111111100101;
   33939: result <= 12'b111111100101;
   33940: result <= 12'b111111100101;
   33941: result <= 12'b111111100101;
   33942: result <= 12'b111111100110;
   33943: result <= 12'b111111100110;
   33944: result <= 12'b111111100110;
   33945: result <= 12'b111111100110;
   33946: result <= 12'b111111100110;
   33947: result <= 12'b111111100111;
   33948: result <= 12'b111111100111;
   33949: result <= 12'b111111100111;
   33950: result <= 12'b111111100111;
   33951: result <= 12'b111111100111;
   33952: result <= 12'b111111100111;
   33953: result <= 12'b111111101000;
   33954: result <= 12'b111111101000;
   33955: result <= 12'b111111101000;
   33956: result <= 12'b111111101000;
   33957: result <= 12'b111111101000;
   33958: result <= 12'b111111101001;
   33959: result <= 12'b111111101001;
   33960: result <= 12'b111111101001;
   33961: result <= 12'b111111101001;
   33962: result <= 12'b111111101001;
   33963: result <= 12'b111111101010;
   33964: result <= 12'b111111101010;
   33965: result <= 12'b111111101010;
   33966: result <= 12'b111111101010;
   33967: result <= 12'b111111101010;
   33968: result <= 12'b111111101011;
   33969: result <= 12'b111111101011;
   33970: result <= 12'b111111101011;
   33971: result <= 12'b111111101011;
   33972: result <= 12'b111111101011;
   33973: result <= 12'b111111101100;
   33974: result <= 12'b111111101100;
   33975: result <= 12'b111111101100;
   33976: result <= 12'b111111101100;
   33977: result <= 12'b111111101100;
   33978: result <= 12'b111111101101;
   33979: result <= 12'b111111101101;
   33980: result <= 12'b111111101101;
   33981: result <= 12'b111111101101;
   33982: result <= 12'b111111101101;
   33983: result <= 12'b111111101110;
   33984: result <= 12'b111111101110;
   33985: result <= 12'b111111101110;
   33986: result <= 12'b111111101110;
   33987: result <= 12'b111111101110;
   33988: result <= 12'b111111101111;
   33989: result <= 12'b111111101111;
   33990: result <= 12'b111111101111;
   33991: result <= 12'b111111101111;
   33992: result <= 12'b111111101111;
   33993: result <= 12'b111111101111;
   33994: result <= 12'b111111110000;
   33995: result <= 12'b111111110000;
   33996: result <= 12'b111111110000;
   33997: result <= 12'b111111110000;
   33998: result <= 12'b111111110000;
   33999: result <= 12'b111111110001;
   34000: result <= 12'b111111110001;
   34001: result <= 12'b111111110001;
   34002: result <= 12'b111111110001;
   34003: result <= 12'b111111110001;
   34004: result <= 12'b111111110010;
   34005: result <= 12'b111111110010;
   34006: result <= 12'b111111110010;
   34007: result <= 12'b111111110010;
   34008: result <= 12'b111111110010;
   34009: result <= 12'b111111110011;
   34010: result <= 12'b111111110011;
   34011: result <= 12'b111111110011;
   34012: result <= 12'b111111110011;
   34013: result <= 12'b111111110011;
   34014: result <= 12'b111111110100;
   34015: result <= 12'b111111110100;
   34016: result <= 12'b111111110100;
   34017: result <= 12'b111111110100;
   34018: result <= 12'b111111110100;
   34019: result <= 12'b111111110101;
   34020: result <= 12'b111111110101;
   34021: result <= 12'b111111110101;
   34022: result <= 12'b111111110101;
   34023: result <= 12'b111111110101;
   34024: result <= 12'b111111110110;
   34025: result <= 12'b111111110110;
   34026: result <= 12'b111111110110;
   34027: result <= 12'b111111110110;
   34028: result <= 12'b111111110110;
   34029: result <= 12'b111111110110;
   34030: result <= 12'b111111110111;
   34031: result <= 12'b111111110111;
   34032: result <= 12'b111111110111;
   34033: result <= 12'b111111110111;
   34034: result <= 12'b111111110111;
   34035: result <= 12'b111111111000;
   34036: result <= 12'b111111111000;
   34037: result <= 12'b111111111000;
   34038: result <= 12'b111111111000;
   34039: result <= 12'b111111111000;
   34040: result <= 12'b111111111001;
   34041: result <= 12'b111111111001;
   34042: result <= 12'b111111111001;
   34043: result <= 12'b111111111001;
   34044: result <= 12'b111111111001;
   34045: result <= 12'b111111111010;
   34046: result <= 12'b111111111010;
   34047: result <= 12'b111111111010;
   34048: result <= 12'b111111111010;
   34049: result <= 12'b111111111010;
   34050: result <= 12'b111111111011;
   34051: result <= 12'b111111111011;
   34052: result <= 12'b111111111011;
   34053: result <= 12'b111111111011;
   34054: result <= 12'b111111111011;
   34055: result <= 12'b111111111100;
   34056: result <= 12'b111111111100;
   34057: result <= 12'b111111111100;
   34058: result <= 12'b111111111100;
   34059: result <= 12'b111111111100;
   34060: result <= 12'b111111111101;
   34061: result <= 12'b111111111101;
   34062: result <= 12'b111111111101;
   34063: result <= 12'b111111111101;
   34064: result <= 12'b111111111101;
   34065: result <= 12'b111111111110;
   34066: result <= 12'b111111111110;
   34067: result <= 12'b111111111110;
   34068: result <= 12'b111111111110;
   34069: result <= 12'b111111111110;
   34070: result <= 12'b111111111110;
   34071: result <= 12'b111111111111;
   34072: result <= 12'b111111111111;
   34073: result <= 12'b111111111111;
   34074: result <= 12'b111111111111;
   34075: result <= 12'b111111111111;
   34076: result <= 12'b111100000000;
   34077: result <= 12'b111100000000;
   34078: result <= 12'b111100000000;
   34079: result <= 12'b111100000000;
   34080: result <= 12'b111100000000;
   34081: result <= 12'b111100000001;
   34082: result <= 12'b111100000001;
   34083: result <= 12'b111100000001;
   34084: result <= 12'b111100000001;
   34085: result <= 12'b111100000001;
   34086: result <= 12'b111100000010;
   34087: result <= 12'b111100000010;
   34088: result <= 12'b111100000010;
   34089: result <= 12'b111100000010;
   34090: result <= 12'b111100000010;
   34091: result <= 12'b111100000011;
   34092: result <= 12'b111100000011;
   34093: result <= 12'b111100000011;
   34094: result <= 12'b111100000011;
   34095: result <= 12'b111100000011;
   34096: result <= 12'b111100000100;
   34097: result <= 12'b111100000100;
   34098: result <= 12'b111100000100;
   34099: result <= 12'b111100000100;
   34100: result <= 12'b111100000100;
   34101: result <= 12'b111100000101;
   34102: result <= 12'b111100000101;
   34103: result <= 12'b111100000101;
   34104: result <= 12'b111100000101;
   34105: result <= 12'b111100000101;
   34106: result <= 12'b111100000101;
   34107: result <= 12'b111100000110;
   34108: result <= 12'b111100000110;
   34109: result <= 12'b111100000110;
   34110: result <= 12'b111100000110;
   34111: result <= 12'b111100000110;
   34112: result <= 12'b111100000111;
   34113: result <= 12'b111100000111;
   34114: result <= 12'b111100000111;
   34115: result <= 12'b111100000111;
   34116: result <= 12'b111100000111;
   34117: result <= 12'b111100001000;
   34118: result <= 12'b111100001000;
   34119: result <= 12'b111100001000;
   34120: result <= 12'b111100001000;
   34121: result <= 12'b111100001000;
   34122: result <= 12'b111100001001;
   34123: result <= 12'b111100001001;
   34124: result <= 12'b111100001001;
   34125: result <= 12'b111100001001;
   34126: result <= 12'b111100001001;
   34127: result <= 12'b111100001010;
   34128: result <= 12'b111100001010;
   34129: result <= 12'b111100001010;
   34130: result <= 12'b111100001010;
   34131: result <= 12'b111100001010;
   34132: result <= 12'b111100001011;
   34133: result <= 12'b111100001011;
   34134: result <= 12'b111100001011;
   34135: result <= 12'b111100001011;
   34136: result <= 12'b111100001011;
   34137: result <= 12'b111100001100;
   34138: result <= 12'b111100001100;
   34139: result <= 12'b111100001100;
   34140: result <= 12'b111100001100;
   34141: result <= 12'b111100001100;
   34142: result <= 12'b111100001101;
   34143: result <= 12'b111100001101;
   34144: result <= 12'b111100001101;
   34145: result <= 12'b111100001101;
   34146: result <= 12'b111100001101;
   34147: result <= 12'b111100001101;
   34148: result <= 12'b111100001110;
   34149: result <= 12'b111100001110;
   34150: result <= 12'b111100001110;
   34151: result <= 12'b111100001110;
   34152: result <= 12'b111100001110;
   34153: result <= 12'b111100001111;
   34154: result <= 12'b111100001111;
   34155: result <= 12'b111100001111;
   34156: result <= 12'b111100001111;
   34157: result <= 12'b111100001111;
   34158: result <= 12'b111100010000;
   34159: result <= 12'b111100010000;
   34160: result <= 12'b111100010000;
   34161: result <= 12'b111100010000;
   34162: result <= 12'b111100010000;
   34163: result <= 12'b111100010001;
   34164: result <= 12'b111100010001;
   34165: result <= 12'b111100010001;
   34166: result <= 12'b111100010001;
   34167: result <= 12'b111100010001;
   34168: result <= 12'b111100010010;
   34169: result <= 12'b111100010010;
   34170: result <= 12'b111100010010;
   34171: result <= 12'b111100010010;
   34172: result <= 12'b111100010010;
   34173: result <= 12'b111100010011;
   34174: result <= 12'b111100010011;
   34175: result <= 12'b111100010011;
   34176: result <= 12'b111100010011;
   34177: result <= 12'b111100010011;
   34178: result <= 12'b111100010100;
   34179: result <= 12'b111100010100;
   34180: result <= 12'b111100010100;
   34181: result <= 12'b111100010100;
   34182: result <= 12'b111100010100;
   34183: result <= 12'b111100010100;
   34184: result <= 12'b111100010101;
   34185: result <= 12'b111100010101;
   34186: result <= 12'b111100010101;
   34187: result <= 12'b111100010101;
   34188: result <= 12'b111100010101;
   34189: result <= 12'b111100010110;
   34190: result <= 12'b111100010110;
   34191: result <= 12'b111100010110;
   34192: result <= 12'b111100010110;
   34193: result <= 12'b111100010110;
   34194: result <= 12'b111100010111;
   34195: result <= 12'b111100010111;
   34196: result <= 12'b111100010111;
   34197: result <= 12'b111100010111;
   34198: result <= 12'b111100010111;
   34199: result <= 12'b111100011000;
   34200: result <= 12'b111100011000;
   34201: result <= 12'b111100011000;
   34202: result <= 12'b111100011000;
   34203: result <= 12'b111100011000;
   34204: result <= 12'b111100011001;
   34205: result <= 12'b111100011001;
   34206: result <= 12'b111100011001;
   34207: result <= 12'b111100011001;
   34208: result <= 12'b111100011001;
   34209: result <= 12'b111100011010;
   34210: result <= 12'b111100011010;
   34211: result <= 12'b111100011010;
   34212: result <= 12'b111100011010;
   34213: result <= 12'b111100011010;
   34214: result <= 12'b111100011011;
   34215: result <= 12'b111100011011;
   34216: result <= 12'b111100011011;
   34217: result <= 12'b111100011011;
   34218: result <= 12'b111100011011;
   34219: result <= 12'b111100011011;
   34220: result <= 12'b111100011100;
   34221: result <= 12'b111100011100;
   34222: result <= 12'b111100011100;
   34223: result <= 12'b111100011100;
   34224: result <= 12'b111100011100;
   34225: result <= 12'b111100011101;
   34226: result <= 12'b111100011101;
   34227: result <= 12'b111100011101;
   34228: result <= 12'b111100011101;
   34229: result <= 12'b111100011101;
   34230: result <= 12'b111100011110;
   34231: result <= 12'b111100011110;
   34232: result <= 12'b111100011110;
   34233: result <= 12'b111100011110;
   34234: result <= 12'b111100011110;
   34235: result <= 12'b111100011111;
   34236: result <= 12'b111100011111;
   34237: result <= 12'b111100011111;
   34238: result <= 12'b111100011111;
   34239: result <= 12'b111100011111;
   34240: result <= 12'b111100100000;
   34241: result <= 12'b111100100000;
   34242: result <= 12'b111100100000;
   34243: result <= 12'b111100100000;
   34244: result <= 12'b111100100000;
   34245: result <= 12'b111100100001;
   34246: result <= 12'b111100100001;
   34247: result <= 12'b111100100001;
   34248: result <= 12'b111100100001;
   34249: result <= 12'b111100100001;
   34250: result <= 12'b111100100010;
   34251: result <= 12'b111100100010;
   34252: result <= 12'b111100100010;
   34253: result <= 12'b111100100010;
   34254: result <= 12'b111100100010;
   34255: result <= 12'b111100100010;
   34256: result <= 12'b111100100011;
   34257: result <= 12'b111100100011;
   34258: result <= 12'b111100100011;
   34259: result <= 12'b111100100011;
   34260: result <= 12'b111100100011;
   34261: result <= 12'b111100100100;
   34262: result <= 12'b111100100100;
   34263: result <= 12'b111100100100;
   34264: result <= 12'b111100100100;
   34265: result <= 12'b111100100100;
   34266: result <= 12'b111100100101;
   34267: result <= 12'b111100100101;
   34268: result <= 12'b111100100101;
   34269: result <= 12'b111100100101;
   34270: result <= 12'b111100100101;
   34271: result <= 12'b111100100110;
   34272: result <= 12'b111100100110;
   34273: result <= 12'b111100100110;
   34274: result <= 12'b111100100110;
   34275: result <= 12'b111100100110;
   34276: result <= 12'b111100100111;
   34277: result <= 12'b111100100111;
   34278: result <= 12'b111100100111;
   34279: result <= 12'b111100100111;
   34280: result <= 12'b111100100111;
   34281: result <= 12'b111100101000;
   34282: result <= 12'b111100101000;
   34283: result <= 12'b111100101000;
   34284: result <= 12'b111100101000;
   34285: result <= 12'b111100101000;
   34286: result <= 12'b111100101001;
   34287: result <= 12'b111100101001;
   34288: result <= 12'b111100101001;
   34289: result <= 12'b111100101001;
   34290: result <= 12'b111100101001;
   34291: result <= 12'b111100101001;
   34292: result <= 12'b111100101010;
   34293: result <= 12'b111100101010;
   34294: result <= 12'b111100101010;
   34295: result <= 12'b111100101010;
   34296: result <= 12'b111100101010;
   34297: result <= 12'b111100101011;
   34298: result <= 12'b111100101011;
   34299: result <= 12'b111100101011;
   34300: result <= 12'b111100101011;
   34301: result <= 12'b111100101011;
   34302: result <= 12'b111100101100;
   34303: result <= 12'b111100101100;
   34304: result <= 12'b111100101100;
   34305: result <= 12'b111100101100;
   34306: result <= 12'b111100101100;
   34307: result <= 12'b111100101101;
   34308: result <= 12'b111100101101;
   34309: result <= 12'b111100101101;
   34310: result <= 12'b111100101101;
   34311: result <= 12'b111100101101;
   34312: result <= 12'b111100101110;
   34313: result <= 12'b111100101110;
   34314: result <= 12'b111100101110;
   34315: result <= 12'b111100101110;
   34316: result <= 12'b111100101110;
   34317: result <= 12'b111100101111;
   34318: result <= 12'b111100101111;
   34319: result <= 12'b111100101111;
   34320: result <= 12'b111100101111;
   34321: result <= 12'b111100101111;
   34322: result <= 12'b111100101111;
   34323: result <= 12'b111100110000;
   34324: result <= 12'b111100110000;
   34325: result <= 12'b111100110000;
   34326: result <= 12'b111100110000;
   34327: result <= 12'b111100110000;
   34328: result <= 12'b111100110001;
   34329: result <= 12'b111100110001;
   34330: result <= 12'b111100110001;
   34331: result <= 12'b111100110001;
   34332: result <= 12'b111100110001;
   34333: result <= 12'b111100110010;
   34334: result <= 12'b111100110010;
   34335: result <= 12'b111100110010;
   34336: result <= 12'b111100110010;
   34337: result <= 12'b111100110010;
   34338: result <= 12'b111100110011;
   34339: result <= 12'b111100110011;
   34340: result <= 12'b111100110011;
   34341: result <= 12'b111100110011;
   34342: result <= 12'b111100110011;
   34343: result <= 12'b111100110100;
   34344: result <= 12'b111100110100;
   34345: result <= 12'b111100110100;
   34346: result <= 12'b111100110100;
   34347: result <= 12'b111100110100;
   34348: result <= 12'b111100110101;
   34349: result <= 12'b111100110101;
   34350: result <= 12'b111100110101;
   34351: result <= 12'b111100110101;
   34352: result <= 12'b111100110101;
   34353: result <= 12'b111100110110;
   34354: result <= 12'b111100110110;
   34355: result <= 12'b111100110110;
   34356: result <= 12'b111100110110;
   34357: result <= 12'b111100110110;
   34358: result <= 12'b111100110110;
   34359: result <= 12'b111100110111;
   34360: result <= 12'b111100110111;
   34361: result <= 12'b111100110111;
   34362: result <= 12'b111100110111;
   34363: result <= 12'b111100110111;
   34364: result <= 12'b111100111000;
   34365: result <= 12'b111100111000;
   34366: result <= 12'b111100111000;
   34367: result <= 12'b111100111000;
   34368: result <= 12'b111100111000;
   34369: result <= 12'b111100111001;
   34370: result <= 12'b111100111001;
   34371: result <= 12'b111100111001;
   34372: result <= 12'b111100111001;
   34373: result <= 12'b111100111001;
   34374: result <= 12'b111100111010;
   34375: result <= 12'b111100111010;
   34376: result <= 12'b111100111010;
   34377: result <= 12'b111100111010;
   34378: result <= 12'b111100111010;
   34379: result <= 12'b111100111011;
   34380: result <= 12'b111100111011;
   34381: result <= 12'b111100111011;
   34382: result <= 12'b111100111011;
   34383: result <= 12'b111100111011;
   34384: result <= 12'b111100111100;
   34385: result <= 12'b111100111100;
   34386: result <= 12'b111100111100;
   34387: result <= 12'b111100111100;
   34388: result <= 12'b111100111100;
   34389: result <= 12'b111100111101;
   34390: result <= 12'b111100111101;
   34391: result <= 12'b111100111101;
   34392: result <= 12'b111100111101;
   34393: result <= 12'b111100111101;
   34394: result <= 12'b111100111101;
   34395: result <= 12'b111100111110;
   34396: result <= 12'b111100111110;
   34397: result <= 12'b111100111110;
   34398: result <= 12'b111100111110;
   34399: result <= 12'b111100111110;
   34400: result <= 12'b111100111111;
   34401: result <= 12'b111100111111;
   34402: result <= 12'b111100111111;
   34403: result <= 12'b111100111111;
   34404: result <= 12'b111100111111;
   34405: result <= 12'b111101000000;
   34406: result <= 12'b111101000000;
   34407: result <= 12'b111101000000;
   34408: result <= 12'b111101000000;
   34409: result <= 12'b111101000000;
   34410: result <= 12'b111101000001;
   34411: result <= 12'b111101000001;
   34412: result <= 12'b111101000001;
   34413: result <= 12'b111101000001;
   34414: result <= 12'b111101000001;
   34415: result <= 12'b111101000010;
   34416: result <= 12'b111101000010;
   34417: result <= 12'b111101000010;
   34418: result <= 12'b111101000010;
   34419: result <= 12'b111101000010;
   34420: result <= 12'b111101000011;
   34421: result <= 12'b111101000011;
   34422: result <= 12'b111101000011;
   34423: result <= 12'b111101000011;
   34424: result <= 12'b111101000011;
   34425: result <= 12'b111101000011;
   34426: result <= 12'b111101000100;
   34427: result <= 12'b111101000100;
   34428: result <= 12'b111101000100;
   34429: result <= 12'b111101000100;
   34430: result <= 12'b111101000100;
   34431: result <= 12'b111101000101;
   34432: result <= 12'b111101000101;
   34433: result <= 12'b111101000101;
   34434: result <= 12'b111101000101;
   34435: result <= 12'b111101000101;
   34436: result <= 12'b111101000110;
   34437: result <= 12'b111101000110;
   34438: result <= 12'b111101000110;
   34439: result <= 12'b111101000110;
   34440: result <= 12'b111101000110;
   34441: result <= 12'b111101000111;
   34442: result <= 12'b111101000111;
   34443: result <= 12'b111101000111;
   34444: result <= 12'b111101000111;
   34445: result <= 12'b111101000111;
   34446: result <= 12'b111101001000;
   34447: result <= 12'b111101001000;
   34448: result <= 12'b111101001000;
   34449: result <= 12'b111101001000;
   34450: result <= 12'b111101001000;
   34451: result <= 12'b111101001001;
   34452: result <= 12'b111101001001;
   34453: result <= 12'b111101001001;
   34454: result <= 12'b111101001001;
   34455: result <= 12'b111101001001;
   34456: result <= 12'b111101001001;
   34457: result <= 12'b111101001010;
   34458: result <= 12'b111101001010;
   34459: result <= 12'b111101001010;
   34460: result <= 12'b111101001010;
   34461: result <= 12'b111101001010;
   34462: result <= 12'b111101001011;
   34463: result <= 12'b111101001011;
   34464: result <= 12'b111101001011;
   34465: result <= 12'b111101001011;
   34466: result <= 12'b111101001011;
   34467: result <= 12'b111101001100;
   34468: result <= 12'b111101001100;
   34469: result <= 12'b111101001100;
   34470: result <= 12'b111101001100;
   34471: result <= 12'b111101001100;
   34472: result <= 12'b111101001101;
   34473: result <= 12'b111101001101;
   34474: result <= 12'b111101001101;
   34475: result <= 12'b111101001101;
   34476: result <= 12'b111101001101;
   34477: result <= 12'b111101001110;
   34478: result <= 12'b111101001110;
   34479: result <= 12'b111101001110;
   34480: result <= 12'b111101001110;
   34481: result <= 12'b111101001110;
   34482: result <= 12'b111101001111;
   34483: result <= 12'b111101001111;
   34484: result <= 12'b111101001111;
   34485: result <= 12'b111101001111;
   34486: result <= 12'b111101001111;
   34487: result <= 12'b111101001111;
   34488: result <= 12'b111101010000;
   34489: result <= 12'b111101010000;
   34490: result <= 12'b111101010000;
   34491: result <= 12'b111101010000;
   34492: result <= 12'b111101010000;
   34493: result <= 12'b111101010001;
   34494: result <= 12'b111101010001;
   34495: result <= 12'b111101010001;
   34496: result <= 12'b111101010001;
   34497: result <= 12'b111101010001;
   34498: result <= 12'b111101010010;
   34499: result <= 12'b111101010010;
   34500: result <= 12'b111101010010;
   34501: result <= 12'b111101010010;
   34502: result <= 12'b111101010010;
   34503: result <= 12'b111101010011;
   34504: result <= 12'b111101010011;
   34505: result <= 12'b111101010011;
   34506: result <= 12'b111101010011;
   34507: result <= 12'b111101010011;
   34508: result <= 12'b111101010100;
   34509: result <= 12'b111101010100;
   34510: result <= 12'b111101010100;
   34511: result <= 12'b111101010100;
   34512: result <= 12'b111101010100;
   34513: result <= 12'b111101010101;
   34514: result <= 12'b111101010101;
   34515: result <= 12'b111101010101;
   34516: result <= 12'b111101010101;
   34517: result <= 12'b111101010101;
   34518: result <= 12'b111101010110;
   34519: result <= 12'b111101010110;
   34520: result <= 12'b111101010110;
   34521: result <= 12'b111101010110;
   34522: result <= 12'b111101010110;
   34523: result <= 12'b111101010110;
   34524: result <= 12'b111101010111;
   34525: result <= 12'b111101010111;
   34526: result <= 12'b111101010111;
   34527: result <= 12'b111101010111;
   34528: result <= 12'b111101010111;
   34529: result <= 12'b111101011000;
   34530: result <= 12'b111101011000;
   34531: result <= 12'b111101011000;
   34532: result <= 12'b111101011000;
   34533: result <= 12'b111101011000;
   34534: result <= 12'b111101011001;
   34535: result <= 12'b111101011001;
   34536: result <= 12'b111101011001;
   34537: result <= 12'b111101011001;
   34538: result <= 12'b111101011001;
   34539: result <= 12'b111101011010;
   34540: result <= 12'b111101011010;
   34541: result <= 12'b111101011010;
   34542: result <= 12'b111101011010;
   34543: result <= 12'b111101011010;
   34544: result <= 12'b111101011011;
   34545: result <= 12'b111101011011;
   34546: result <= 12'b111101011011;
   34547: result <= 12'b111101011011;
   34548: result <= 12'b111101011011;
   34549: result <= 12'b111101011100;
   34550: result <= 12'b111101011100;
   34551: result <= 12'b111101011100;
   34552: result <= 12'b111101011100;
   34553: result <= 12'b111101011100;
   34554: result <= 12'b111101011100;
   34555: result <= 12'b111101011101;
   34556: result <= 12'b111101011101;
   34557: result <= 12'b111101011101;
   34558: result <= 12'b111101011101;
   34559: result <= 12'b111101011101;
   34560: result <= 12'b111101011110;
   34561: result <= 12'b111101011110;
   34562: result <= 12'b111101011110;
   34563: result <= 12'b111101011110;
   34564: result <= 12'b111101011110;
   34565: result <= 12'b111101011111;
   34566: result <= 12'b111101011111;
   34567: result <= 12'b111101011111;
   34568: result <= 12'b111101011111;
   34569: result <= 12'b111101011111;
   34570: result <= 12'b111101100000;
   34571: result <= 12'b111101100000;
   34572: result <= 12'b111101100000;
   34573: result <= 12'b111101100000;
   34574: result <= 12'b111101100000;
   34575: result <= 12'b111101100001;
   34576: result <= 12'b111101100001;
   34577: result <= 12'b111101100001;
   34578: result <= 12'b111101100001;
   34579: result <= 12'b111101100001;
   34580: result <= 12'b111101100001;
   34581: result <= 12'b111101100010;
   34582: result <= 12'b111101100010;
   34583: result <= 12'b111101100010;
   34584: result <= 12'b111101100010;
   34585: result <= 12'b111101100010;
   34586: result <= 12'b111101100011;
   34587: result <= 12'b111101100011;
   34588: result <= 12'b111101100011;
   34589: result <= 12'b111101100011;
   34590: result <= 12'b111101100011;
   34591: result <= 12'b111101100100;
   34592: result <= 12'b111101100100;
   34593: result <= 12'b111101100100;
   34594: result <= 12'b111101100100;
   34595: result <= 12'b111101100100;
   34596: result <= 12'b111101100101;
   34597: result <= 12'b111101100101;
   34598: result <= 12'b111101100101;
   34599: result <= 12'b111101100101;
   34600: result <= 12'b111101100101;
   34601: result <= 12'b111101100110;
   34602: result <= 12'b111101100110;
   34603: result <= 12'b111101100110;
   34604: result <= 12'b111101100110;
   34605: result <= 12'b111101100110;
   34606: result <= 12'b111101100111;
   34607: result <= 12'b111101100111;
   34608: result <= 12'b111101100111;
   34609: result <= 12'b111101100111;
   34610: result <= 12'b111101100111;
   34611: result <= 12'b111101100111;
   34612: result <= 12'b111101101000;
   34613: result <= 12'b111101101000;
   34614: result <= 12'b111101101000;
   34615: result <= 12'b111101101000;
   34616: result <= 12'b111101101000;
   34617: result <= 12'b111101101001;
   34618: result <= 12'b111101101001;
   34619: result <= 12'b111101101001;
   34620: result <= 12'b111101101001;
   34621: result <= 12'b111101101001;
   34622: result <= 12'b111101101010;
   34623: result <= 12'b111101101010;
   34624: result <= 12'b111101101010;
   34625: result <= 12'b111101101010;
   34626: result <= 12'b111101101010;
   34627: result <= 12'b111101101011;
   34628: result <= 12'b111101101011;
   34629: result <= 12'b111101101011;
   34630: result <= 12'b111101101011;
   34631: result <= 12'b111101101011;
   34632: result <= 12'b111101101100;
   34633: result <= 12'b111101101100;
   34634: result <= 12'b111101101100;
   34635: result <= 12'b111101101100;
   34636: result <= 12'b111101101100;
   34637: result <= 12'b111101101101;
   34638: result <= 12'b111101101101;
   34639: result <= 12'b111101101101;
   34640: result <= 12'b111101101101;
   34641: result <= 12'b111101101101;
   34642: result <= 12'b111101101101;
   34643: result <= 12'b111101101110;
   34644: result <= 12'b111101101110;
   34645: result <= 12'b111101101110;
   34646: result <= 12'b111101101110;
   34647: result <= 12'b111101101110;
   34648: result <= 12'b111101101111;
   34649: result <= 12'b111101101111;
   34650: result <= 12'b111101101111;
   34651: result <= 12'b111101101111;
   34652: result <= 12'b111101101111;
   34653: result <= 12'b111101110000;
   34654: result <= 12'b111101110000;
   34655: result <= 12'b111101110000;
   34656: result <= 12'b111101110000;
   34657: result <= 12'b111101110000;
   34658: result <= 12'b111101110001;
   34659: result <= 12'b111101110001;
   34660: result <= 12'b111101110001;
   34661: result <= 12'b111101110001;
   34662: result <= 12'b111101110001;
   34663: result <= 12'b111101110010;
   34664: result <= 12'b111101110010;
   34665: result <= 12'b111101110010;
   34666: result <= 12'b111101110010;
   34667: result <= 12'b111101110010;
   34668: result <= 12'b111101110011;
   34669: result <= 12'b111101110011;
   34670: result <= 12'b111101110011;
   34671: result <= 12'b111101110011;
   34672: result <= 12'b111101110011;
   34673: result <= 12'b111101110011;
   34674: result <= 12'b111101110100;
   34675: result <= 12'b111101110100;
   34676: result <= 12'b111101110100;
   34677: result <= 12'b111101110100;
   34678: result <= 12'b111101110100;
   34679: result <= 12'b111101110101;
   34680: result <= 12'b111101110101;
   34681: result <= 12'b111101110101;
   34682: result <= 12'b111101110101;
   34683: result <= 12'b111101110101;
   34684: result <= 12'b111101110110;
   34685: result <= 12'b111101110110;
   34686: result <= 12'b111101110110;
   34687: result <= 12'b111101110110;
   34688: result <= 12'b111101110110;
   34689: result <= 12'b111101110111;
   34690: result <= 12'b111101110111;
   34691: result <= 12'b111101110111;
   34692: result <= 12'b111101110111;
   34693: result <= 12'b111101110111;
   34694: result <= 12'b111101111000;
   34695: result <= 12'b111101111000;
   34696: result <= 12'b111101111000;
   34697: result <= 12'b111101111000;
   34698: result <= 12'b111101111000;
   34699: result <= 12'b111101111000;
   34700: result <= 12'b111101111001;
   34701: result <= 12'b111101111001;
   34702: result <= 12'b111101111001;
   34703: result <= 12'b111101111001;
   34704: result <= 12'b111101111001;
   34705: result <= 12'b111101111010;
   34706: result <= 12'b111101111010;
   34707: result <= 12'b111101111010;
   34708: result <= 12'b111101111010;
   34709: result <= 12'b111101111010;
   34710: result <= 12'b111101111011;
   34711: result <= 12'b111101111011;
   34712: result <= 12'b111101111011;
   34713: result <= 12'b111101111011;
   34714: result <= 12'b111101111011;
   34715: result <= 12'b111101111100;
   34716: result <= 12'b111101111100;
   34717: result <= 12'b111101111100;
   34718: result <= 12'b111101111100;
   34719: result <= 12'b111101111100;
   34720: result <= 12'b111101111101;
   34721: result <= 12'b111101111101;
   34722: result <= 12'b111101111101;
   34723: result <= 12'b111101111101;
   34724: result <= 12'b111101111101;
   34725: result <= 12'b111101111110;
   34726: result <= 12'b111101111110;
   34727: result <= 12'b111101111110;
   34728: result <= 12'b111101111110;
   34729: result <= 12'b111101111110;
   34730: result <= 12'b111101111110;
   34731: result <= 12'b111101111111;
   34732: result <= 12'b111101111111;
   34733: result <= 12'b111101111111;
   34734: result <= 12'b111101111111;
   34735: result <= 12'b111101111111;
   34736: result <= 12'b111110000000;
   34737: result <= 12'b111110000000;
   34738: result <= 12'b111110000000;
   34739: result <= 12'b111110000000;
   34740: result <= 12'b111110000000;
   34741: result <= 12'b111110000001;
   34742: result <= 12'b111110000001;
   34743: result <= 12'b111110000001;
   34744: result <= 12'b111110000001;
   34745: result <= 12'b111110000001;
   34746: result <= 12'b111110000010;
   34747: result <= 12'b111110000010;
   34748: result <= 12'b111110000010;
   34749: result <= 12'b111110000010;
   34750: result <= 12'b111110000010;
   34751: result <= 12'b111110000011;
   34752: result <= 12'b111110000011;
   34753: result <= 12'b111110000011;
   34754: result <= 12'b111110000011;
   34755: result <= 12'b111110000011;
   34756: result <= 12'b111110000011;
   34757: result <= 12'b111110000100;
   34758: result <= 12'b111110000100;
   34759: result <= 12'b111110000100;
   34760: result <= 12'b111110000100;
   34761: result <= 12'b111110000100;
   34762: result <= 12'b111110000101;
   34763: result <= 12'b111110000101;
   34764: result <= 12'b111110000101;
   34765: result <= 12'b111110000101;
   34766: result <= 12'b111110000101;
   34767: result <= 12'b111110000110;
   34768: result <= 12'b111110000110;
   34769: result <= 12'b111110000110;
   34770: result <= 12'b111110000110;
   34771: result <= 12'b111110000110;
   34772: result <= 12'b111110000111;
   34773: result <= 12'b111110000111;
   34774: result <= 12'b111110000111;
   34775: result <= 12'b111110000111;
   34776: result <= 12'b111110000111;
   34777: result <= 12'b111110001000;
   34778: result <= 12'b111110001000;
   34779: result <= 12'b111110001000;
   34780: result <= 12'b111110001000;
   34781: result <= 12'b111110001000;
   34782: result <= 12'b111110001000;
   34783: result <= 12'b111110001001;
   34784: result <= 12'b111110001001;
   34785: result <= 12'b111110001001;
   34786: result <= 12'b111110001001;
   34787: result <= 12'b111110001001;
   34788: result <= 12'b111110001010;
   34789: result <= 12'b111110001010;
   34790: result <= 12'b111110001010;
   34791: result <= 12'b111110001010;
   34792: result <= 12'b111110001010;
   34793: result <= 12'b111110001011;
   34794: result <= 12'b111110001011;
   34795: result <= 12'b111110001011;
   34796: result <= 12'b111110001011;
   34797: result <= 12'b111110001011;
   34798: result <= 12'b111110001100;
   34799: result <= 12'b111110001100;
   34800: result <= 12'b111110001100;
   34801: result <= 12'b111110001100;
   34802: result <= 12'b111110001100;
   34803: result <= 12'b111110001101;
   34804: result <= 12'b111110001101;
   34805: result <= 12'b111110001101;
   34806: result <= 12'b111110001101;
   34807: result <= 12'b111110001101;
   34808: result <= 12'b111110001110;
   34809: result <= 12'b111110001110;
   34810: result <= 12'b111110001110;
   34811: result <= 12'b111110001110;
   34812: result <= 12'b111110001110;
   34813: result <= 12'b111110001110;
   34814: result <= 12'b111110001111;
   34815: result <= 12'b111110001111;
   34816: result <= 12'b111110001111;
   34817: result <= 12'b111110001111;
   34818: result <= 12'b111110001111;
   34819: result <= 12'b111110010000;
   34820: result <= 12'b111110010000;
   34821: result <= 12'b111110010000;
   34822: result <= 12'b111110010000;
   34823: result <= 12'b111110010000;
   34824: result <= 12'b111110010001;
   34825: result <= 12'b111110010001;
   34826: result <= 12'b111110010001;
   34827: result <= 12'b111110010001;
   34828: result <= 12'b111110010001;
   34829: result <= 12'b111110010010;
   34830: result <= 12'b111110010010;
   34831: result <= 12'b111110010010;
   34832: result <= 12'b111110010010;
   34833: result <= 12'b111110010010;
   34834: result <= 12'b111110010011;
   34835: result <= 12'b111110010011;
   34836: result <= 12'b111110010011;
   34837: result <= 12'b111110010011;
   34838: result <= 12'b111110010011;
   34839: result <= 12'b111110010011;
   34840: result <= 12'b111110010100;
   34841: result <= 12'b111110010100;
   34842: result <= 12'b111110010100;
   34843: result <= 12'b111110010100;
   34844: result <= 12'b111110010100;
   34845: result <= 12'b111110010101;
   34846: result <= 12'b111110010101;
   34847: result <= 12'b111110010101;
   34848: result <= 12'b111110010101;
   34849: result <= 12'b111110010101;
   34850: result <= 12'b111110010110;
   34851: result <= 12'b111110010110;
   34852: result <= 12'b111110010110;
   34853: result <= 12'b111110010110;
   34854: result <= 12'b111110010110;
   34855: result <= 12'b111110010111;
   34856: result <= 12'b111110010111;
   34857: result <= 12'b111110010111;
   34858: result <= 12'b111110010111;
   34859: result <= 12'b111110010111;
   34860: result <= 12'b111110011000;
   34861: result <= 12'b111110011000;
   34862: result <= 12'b111110011000;
   34863: result <= 12'b111110011000;
   34864: result <= 12'b111110011000;
   34865: result <= 12'b111110011000;
   34866: result <= 12'b111110011001;
   34867: result <= 12'b111110011001;
   34868: result <= 12'b111110011001;
   34869: result <= 12'b111110011001;
   34870: result <= 12'b111110011001;
   34871: result <= 12'b111110011010;
   34872: result <= 12'b111110011010;
   34873: result <= 12'b111110011010;
   34874: result <= 12'b111110011010;
   34875: result <= 12'b111110011010;
   34876: result <= 12'b111110011011;
   34877: result <= 12'b111110011011;
   34878: result <= 12'b111110011011;
   34879: result <= 12'b111110011011;
   34880: result <= 12'b111110011011;
   34881: result <= 12'b111110011100;
   34882: result <= 12'b111110011100;
   34883: result <= 12'b111110011100;
   34884: result <= 12'b111110011100;
   34885: result <= 12'b111110011100;
   34886: result <= 12'b111110011101;
   34887: result <= 12'b111110011101;
   34888: result <= 12'b111110011101;
   34889: result <= 12'b111110011101;
   34890: result <= 12'b111110011101;
   34891: result <= 12'b111110011101;
   34892: result <= 12'b111110011110;
   34893: result <= 12'b111110011110;
   34894: result <= 12'b111110011110;
   34895: result <= 12'b111110011110;
   34896: result <= 12'b111110011110;
   34897: result <= 12'b111110011111;
   34898: result <= 12'b111110011111;
   34899: result <= 12'b111110011111;
   34900: result <= 12'b111110011111;
   34901: result <= 12'b111110011111;
   34902: result <= 12'b111110100000;
   34903: result <= 12'b111110100000;
   34904: result <= 12'b111110100000;
   34905: result <= 12'b111110100000;
   34906: result <= 12'b111110100000;
   34907: result <= 12'b111110100001;
   34908: result <= 12'b111110100001;
   34909: result <= 12'b111110100001;
   34910: result <= 12'b111110100001;
   34911: result <= 12'b111110100001;
   34912: result <= 12'b111110100010;
   34913: result <= 12'b111110100010;
   34914: result <= 12'b111110100010;
   34915: result <= 12'b111110100010;
   34916: result <= 12'b111110100010;
   34917: result <= 12'b111110100010;
   34918: result <= 12'b111110100011;
   34919: result <= 12'b111110100011;
   34920: result <= 12'b111110100011;
   34921: result <= 12'b111110100011;
   34922: result <= 12'b111110100011;
   34923: result <= 12'b111110100100;
   34924: result <= 12'b111110100100;
   34925: result <= 12'b111110100100;
   34926: result <= 12'b111110100100;
   34927: result <= 12'b111110100100;
   34928: result <= 12'b111110100101;
   34929: result <= 12'b111110100101;
   34930: result <= 12'b111110100101;
   34931: result <= 12'b111110100101;
   34932: result <= 12'b111110100101;
   34933: result <= 12'b111110100110;
   34934: result <= 12'b111110100110;
   34935: result <= 12'b111110100110;
   34936: result <= 12'b111110100110;
   34937: result <= 12'b111110100110;
   34938: result <= 12'b111110100111;
   34939: result <= 12'b111110100111;
   34940: result <= 12'b111110100111;
   34941: result <= 12'b111110100111;
   34942: result <= 12'b111110100111;
   34943: result <= 12'b111110100111;
   34944: result <= 12'b111110101000;
   34945: result <= 12'b111110101000;
   34946: result <= 12'b111110101000;
   34947: result <= 12'b111110101000;
   34948: result <= 12'b111110101000;
   34949: result <= 12'b111110101001;
   34950: result <= 12'b111110101001;
   34951: result <= 12'b111110101001;
   34952: result <= 12'b111110101001;
   34953: result <= 12'b111110101001;
   34954: result <= 12'b111110101010;
   34955: result <= 12'b111110101010;
   34956: result <= 12'b111110101010;
   34957: result <= 12'b111110101010;
   34958: result <= 12'b111110101010;
   34959: result <= 12'b111110101011;
   34960: result <= 12'b111110101011;
   34961: result <= 12'b111110101011;
   34962: result <= 12'b111110101011;
   34963: result <= 12'b111110101011;
   34964: result <= 12'b111110101100;
   34965: result <= 12'b111110101100;
   34966: result <= 12'b111110101100;
   34967: result <= 12'b111110101100;
   34968: result <= 12'b111110101100;
   34969: result <= 12'b111110101100;
   34970: result <= 12'b111110101101;
   34971: result <= 12'b111110101101;
   34972: result <= 12'b111110101101;
   34973: result <= 12'b111110101101;
   34974: result <= 12'b111110101101;
   34975: result <= 12'b111110101110;
   34976: result <= 12'b111110101110;
   34977: result <= 12'b111110101110;
   34978: result <= 12'b111110101110;
   34979: result <= 12'b111110101110;
   34980: result <= 12'b111110101111;
   34981: result <= 12'b111110101111;
   34982: result <= 12'b111110101111;
   34983: result <= 12'b111110101111;
   34984: result <= 12'b111110101111;
   34985: result <= 12'b111110110000;
   34986: result <= 12'b111110110000;
   34987: result <= 12'b111110110000;
   34988: result <= 12'b111110110000;
   34989: result <= 12'b111110110000;
   34990: result <= 12'b111110110000;
   34991: result <= 12'b111110110001;
   34992: result <= 12'b111110110001;
   34993: result <= 12'b111110110001;
   34994: result <= 12'b111110110001;
   34995: result <= 12'b111110110001;
   34996: result <= 12'b111110110010;
   34997: result <= 12'b111110110010;
   34998: result <= 12'b111110110010;
   34999: result <= 12'b111110110010;
   35000: result <= 12'b111110110010;
   35001: result <= 12'b111110110011;
   35002: result <= 12'b111110110011;
   35003: result <= 12'b111110110011;
   35004: result <= 12'b111110110011;
   35005: result <= 12'b111110110011;
   35006: result <= 12'b111110110100;
   35007: result <= 12'b111110110100;
   35008: result <= 12'b111110110100;
   35009: result <= 12'b111110110100;
   35010: result <= 12'b111110110100;
   35011: result <= 12'b111110110101;
   35012: result <= 12'b111110110101;
   35013: result <= 12'b111110110101;
   35014: result <= 12'b111110110101;
   35015: result <= 12'b111110110101;
   35016: result <= 12'b111110110101;
   35017: result <= 12'b111110110110;
   35018: result <= 12'b111110110110;
   35019: result <= 12'b111110110110;
   35020: result <= 12'b111110110110;
   35021: result <= 12'b111110110110;
   35022: result <= 12'b111110110111;
   35023: result <= 12'b111110110111;
   35024: result <= 12'b111110110111;
   35025: result <= 12'b111110110111;
   35026: result <= 12'b111110110111;
   35027: result <= 12'b111110111000;
   35028: result <= 12'b111110111000;
   35029: result <= 12'b111110111000;
   35030: result <= 12'b111110111000;
   35031: result <= 12'b111110111000;
   35032: result <= 12'b111110111001;
   35033: result <= 12'b111110111001;
   35034: result <= 12'b111110111001;
   35035: result <= 12'b111110111001;
   35036: result <= 12'b111110111001;
   35037: result <= 12'b111110111010;
   35038: result <= 12'b111110111010;
   35039: result <= 12'b111110111010;
   35040: result <= 12'b111110111010;
   35041: result <= 12'b111110111010;
   35042: result <= 12'b111110111010;
   35043: result <= 12'b111110111011;
   35044: result <= 12'b111110111011;
   35045: result <= 12'b111110111011;
   35046: result <= 12'b111110111011;
   35047: result <= 12'b111110111011;
   35048: result <= 12'b111110111100;
   35049: result <= 12'b111110111100;
   35050: result <= 12'b111110111100;
   35051: result <= 12'b111110111100;
   35052: result <= 12'b111110111100;
   35053: result <= 12'b111110111101;
   35054: result <= 12'b111110111101;
   35055: result <= 12'b111110111101;
   35056: result <= 12'b111110111101;
   35057: result <= 12'b111110111101;
   35058: result <= 12'b111110111110;
   35059: result <= 12'b111110111110;
   35060: result <= 12'b111110111110;
   35061: result <= 12'b111110111110;
   35062: result <= 12'b111110111110;
   35063: result <= 12'b111110111110;
   35064: result <= 12'b111110111111;
   35065: result <= 12'b111110111111;
   35066: result <= 12'b111110111111;
   35067: result <= 12'b111110111111;
   35068: result <= 12'b111110111111;
   35069: result <= 12'b111111000000;
   35070: result <= 12'b111111000000;
   35071: result <= 12'b111111000000;
   35072: result <= 12'b111111000000;
   35073: result <= 12'b111111000000;
   35074: result <= 12'b111111000001;
   35075: result <= 12'b111111000001;
   35076: result <= 12'b111111000001;
   35077: result <= 12'b111111000001;
   35078: result <= 12'b111111000001;
   35079: result <= 12'b111111000010;
   35080: result <= 12'b111111000010;
   35081: result <= 12'b111111000010;
   35082: result <= 12'b111111000010;
   35083: result <= 12'b111111000010;
   35084: result <= 12'b111111000011;
   35085: result <= 12'b111111000011;
   35086: result <= 12'b111111000011;
   35087: result <= 12'b111111000011;
   35088: result <= 12'b111111000011;
   35089: result <= 12'b111111000011;
   35090: result <= 12'b111111000100;
   35091: result <= 12'b111111000100;
   35092: result <= 12'b111111000100;
   35093: result <= 12'b111111000100;
   35094: result <= 12'b111111000100;
   35095: result <= 12'b111111000101;
   35096: result <= 12'b111111000101;
   35097: result <= 12'b111111000101;
   35098: result <= 12'b111111000101;
   35099: result <= 12'b111111000101;
   35100: result <= 12'b111111000110;
   35101: result <= 12'b111111000110;
   35102: result <= 12'b111111000110;
   35103: result <= 12'b111111000110;
   35104: result <= 12'b111111000110;
   35105: result <= 12'b111111000111;
   35106: result <= 12'b111111000111;
   35107: result <= 12'b111111000111;
   35108: result <= 12'b111111000111;
   35109: result <= 12'b111111000111;
   35110: result <= 12'b111111000111;
   35111: result <= 12'b111111001000;
   35112: result <= 12'b111111001000;
   35113: result <= 12'b111111001000;
   35114: result <= 12'b111111001000;
   35115: result <= 12'b111111001000;
   35116: result <= 12'b111111001001;
   35117: result <= 12'b111111001001;
   35118: result <= 12'b111111001001;
   35119: result <= 12'b111111001001;
   35120: result <= 12'b111111001001;
   35121: result <= 12'b111111001010;
   35122: result <= 12'b111111001010;
   35123: result <= 12'b111111001010;
   35124: result <= 12'b111111001010;
   35125: result <= 12'b111111001010;
   35126: result <= 12'b111111001011;
   35127: result <= 12'b111111001011;
   35128: result <= 12'b111111001011;
   35129: result <= 12'b111111001011;
   35130: result <= 12'b111111001011;
   35131: result <= 12'b111111001100;
   35132: result <= 12'b111111001100;
   35133: result <= 12'b111111001100;
   35134: result <= 12'b111111001100;
   35135: result <= 12'b111111001100;
   35136: result <= 12'b111111001100;
   35137: result <= 12'b111111001101;
   35138: result <= 12'b111111001101;
   35139: result <= 12'b111111001101;
   35140: result <= 12'b111111001101;
   35141: result <= 12'b111111001101;
   35142: result <= 12'b111111001110;
   35143: result <= 12'b111111001110;
   35144: result <= 12'b111111001110;
   35145: result <= 12'b111111001110;
   35146: result <= 12'b111111001110;
   35147: result <= 12'b111111001111;
   35148: result <= 12'b111111001111;
   35149: result <= 12'b111111001111;
   35150: result <= 12'b111111001111;
   35151: result <= 12'b111111001111;
   35152: result <= 12'b111111010000;
   35153: result <= 12'b111111010000;
   35154: result <= 12'b111111010000;
   35155: result <= 12'b111111010000;
   35156: result <= 12'b111111010000;
   35157: result <= 12'b111111010000;
   35158: result <= 12'b111111010001;
   35159: result <= 12'b111111010001;
   35160: result <= 12'b111111010001;
   35161: result <= 12'b111111010001;
   35162: result <= 12'b111111010001;
   35163: result <= 12'b111111010010;
   35164: result <= 12'b111111010010;
   35165: result <= 12'b111111010010;
   35166: result <= 12'b111111010010;
   35167: result <= 12'b111111010010;
   35168: result <= 12'b111111010011;
   35169: result <= 12'b111111010011;
   35170: result <= 12'b111111010011;
   35171: result <= 12'b111111010011;
   35172: result <= 12'b111111010011;
   35173: result <= 12'b111111010100;
   35174: result <= 12'b111111010100;
   35175: result <= 12'b111111010100;
   35176: result <= 12'b111111010100;
   35177: result <= 12'b111111010100;
   35178: result <= 12'b111111010101;
   35179: result <= 12'b111111010101;
   35180: result <= 12'b111111010101;
   35181: result <= 12'b111111010101;
   35182: result <= 12'b111111010101;
   35183: result <= 12'b111111010101;
   35184: result <= 12'b111111010110;
   35185: result <= 12'b111111010110;
   35186: result <= 12'b111111010110;
   35187: result <= 12'b111111010110;
   35188: result <= 12'b111111010110;
   35189: result <= 12'b111111010111;
   35190: result <= 12'b111111010111;
   35191: result <= 12'b111111010111;
   35192: result <= 12'b111111010111;
   35193: result <= 12'b111111010111;
   35194: result <= 12'b111111011000;
   35195: result <= 12'b111111011000;
   35196: result <= 12'b111111011000;
   35197: result <= 12'b111111011000;
   35198: result <= 12'b111111011000;
   35199: result <= 12'b111111011001;
   35200: result <= 12'b111111011001;
   35201: result <= 12'b111111011001;
   35202: result <= 12'b111111011001;
   35203: result <= 12'b111111011001;
   35204: result <= 12'b111111011001;
   35205: result <= 12'b111111011010;
   35206: result <= 12'b111111011010;
   35207: result <= 12'b111111011010;
   35208: result <= 12'b111111011010;
   35209: result <= 12'b111111011010;
   35210: result <= 12'b111111011011;
   35211: result <= 12'b111111011011;
   35212: result <= 12'b111111011011;
   35213: result <= 12'b111111011011;
   35214: result <= 12'b111111011011;
   35215: result <= 12'b111111011100;
   35216: result <= 12'b111111011100;
   35217: result <= 12'b111111011100;
   35218: result <= 12'b111111011100;
   35219: result <= 12'b111111011100;
   35220: result <= 12'b111111011101;
   35221: result <= 12'b111111011101;
   35222: result <= 12'b111111011101;
   35223: result <= 12'b111111011101;
   35224: result <= 12'b111111011101;
   35225: result <= 12'b111111011101;
   35226: result <= 12'b111111011110;
   35227: result <= 12'b111111011110;
   35228: result <= 12'b111111011110;
   35229: result <= 12'b111111011110;
   35230: result <= 12'b111111011110;
   35231: result <= 12'b111111011111;
   35232: result <= 12'b111111011111;
   35233: result <= 12'b111111011111;
   35234: result <= 12'b111111011111;
   35235: result <= 12'b111111011111;
   35236: result <= 12'b111111100000;
   35237: result <= 12'b111111100000;
   35238: result <= 12'b111111100000;
   35239: result <= 12'b111111100000;
   35240: result <= 12'b111111100000;
   35241: result <= 12'b111111100001;
   35242: result <= 12'b111111100001;
   35243: result <= 12'b111111100001;
   35244: result <= 12'b111111100001;
   35245: result <= 12'b111111100001;
   35246: result <= 12'b111111100001;
   35247: result <= 12'b111111100010;
   35248: result <= 12'b111111100010;
   35249: result <= 12'b111111100010;
   35250: result <= 12'b111111100010;
   35251: result <= 12'b111111100010;
   35252: result <= 12'b111111100011;
   35253: result <= 12'b111111100011;
   35254: result <= 12'b111111100011;
   35255: result <= 12'b111111100011;
   35256: result <= 12'b111111100011;
   35257: result <= 12'b111111100100;
   35258: result <= 12'b111111100100;
   35259: result <= 12'b111111100100;
   35260: result <= 12'b111111100100;
   35261: result <= 12'b111111100100;
   35262: result <= 12'b111111100101;
   35263: result <= 12'b111111100101;
   35264: result <= 12'b111111100101;
   35265: result <= 12'b111111100101;
   35266: result <= 12'b111111100101;
   35267: result <= 12'b111111100101;
   35268: result <= 12'b111111100110;
   35269: result <= 12'b111111100110;
   35270: result <= 12'b111111100110;
   35271: result <= 12'b111111100110;
   35272: result <= 12'b111111100110;
   35273: result <= 12'b111111100111;
   35274: result <= 12'b111111100111;
   35275: result <= 12'b111111100111;
   35276: result <= 12'b111111100111;
   35277: result <= 12'b111111100111;
   35278: result <= 12'b111111101000;
   35279: result <= 12'b111111101000;
   35280: result <= 12'b111111101000;
   35281: result <= 12'b111111101000;
   35282: result <= 12'b111111101000;
   35283: result <= 12'b111111101001;
   35284: result <= 12'b111111101001;
   35285: result <= 12'b111111101001;
   35286: result <= 12'b111111101001;
   35287: result <= 12'b111111101001;
   35288: result <= 12'b111111101010;
   35289: result <= 12'b111111101010;
   35290: result <= 12'b111111101010;
   35291: result <= 12'b111111101010;
   35292: result <= 12'b111111101010;
   35293: result <= 12'b111111101010;
   35294: result <= 12'b111111101011;
   35295: result <= 12'b111111101011;
   35296: result <= 12'b111111101011;
   35297: result <= 12'b111111101011;
   35298: result <= 12'b111111101011;
   35299: result <= 12'b111111101100;
   35300: result <= 12'b111111101100;
   35301: result <= 12'b111111101100;
   35302: result <= 12'b111111101100;
   35303: result <= 12'b111111101100;
   35304: result <= 12'b111111101101;
   35305: result <= 12'b111111101101;
   35306: result <= 12'b111111101101;
   35307: result <= 12'b111111101101;
   35308: result <= 12'b111111101101;
   35309: result <= 12'b111111101110;
   35310: result <= 12'b111111101110;
   35311: result <= 12'b111111101110;
   35312: result <= 12'b111111101110;
   35313: result <= 12'b111111101110;
   35314: result <= 12'b111111101110;
   35315: result <= 12'b111111101111;
   35316: result <= 12'b111111101111;
   35317: result <= 12'b111111101111;
   35318: result <= 12'b111111101111;
   35319: result <= 12'b111111101111;
   35320: result <= 12'b111111110000;
   35321: result <= 12'b111111110000;
   35322: result <= 12'b111111110000;
   35323: result <= 12'b111111110000;
   35324: result <= 12'b111111110000;
   35325: result <= 12'b111111110001;
   35326: result <= 12'b111111110001;
   35327: result <= 12'b111111110001;
   35328: result <= 12'b111111110001;
   35329: result <= 12'b111111110001;
   35330: result <= 12'b111111110010;
   35331: result <= 12'b111111110010;
   35332: result <= 12'b111111110010;
   35333: result <= 12'b111111110010;
   35334: result <= 12'b111111110010;
   35335: result <= 12'b111111110010;
   35336: result <= 12'b111111110011;
   35337: result <= 12'b111111110011;
   35338: result <= 12'b111111110011;
   35339: result <= 12'b111111110011;
   35340: result <= 12'b111111110011;
   35341: result <= 12'b111111110100;
   35342: result <= 12'b111111110100;
   35343: result <= 12'b111111110100;
   35344: result <= 12'b111111110100;
   35345: result <= 12'b111111110100;
   35346: result <= 12'b111111110101;
   35347: result <= 12'b111111110101;
   35348: result <= 12'b111111110101;
   35349: result <= 12'b111111110101;
   35350: result <= 12'b111111110101;
   35351: result <= 12'b111111110110;
   35352: result <= 12'b111111110110;
   35353: result <= 12'b111111110110;
   35354: result <= 12'b111111110110;
   35355: result <= 12'b111111110110;
   35356: result <= 12'b111111110110;
   35357: result <= 12'b111111110111;
   35358: result <= 12'b111111110111;
   35359: result <= 12'b111111110111;
   35360: result <= 12'b111111110111;
   35361: result <= 12'b111111110111;
   35362: result <= 12'b111111111000;
   35363: result <= 12'b111111111000;
   35364: result <= 12'b111111111000;
   35365: result <= 12'b111111111000;
   35366: result <= 12'b111111111000;
   35367: result <= 12'b111111111001;
   35368: result <= 12'b111111111001;
   35369: result <= 12'b111111111001;
   35370: result <= 12'b111111111001;
   35371: result <= 12'b111111111001;
   35372: result <= 12'b111111111001;
   35373: result <= 12'b111111111010;
   35374: result <= 12'b111111111010;
   35375: result <= 12'b111111111010;
   35376: result <= 12'b111111111010;
   35377: result <= 12'b111111111010;
   35378: result <= 12'b111111111011;
   35379: result <= 12'b111111111011;
   35380: result <= 12'b111111111011;
   35381: result <= 12'b111111111011;
   35382: result <= 12'b111111111011;
   35383: result <= 12'b111111111100;
   35384: result <= 12'b111111111100;
   35385: result <= 12'b111111111100;
   35386: result <= 12'b111111111100;
   35387: result <= 12'b111111111100;
   35388: result <= 12'b111111111101;
   35389: result <= 12'b111111111101;
   35390: result <= 12'b111111111101;
   35391: result <= 12'b111111111101;
   35392: result <= 12'b111111111101;
   35393: result <= 12'b111111111101;
   35394: result <= 12'b111111111110;
   35395: result <= 12'b111111111110;
   35396: result <= 12'b111111111110;
   35397: result <= 12'b111111111110;
   35398: result <= 12'b111111111110;
   35399: result <= 12'b111111111111;
   35400: result <= 12'b111111111111;
   35401: result <= 12'b111111111111;
   35402: result <= 12'b111111111111;
   35403: result <= 12'b111111111111;
   35404: result <= 12'b111000000000;
   35405: result <= 12'b111000000000;
   35406: result <= 12'b111000000000;
   35407: result <= 12'b111000000000;
   35408: result <= 12'b111000000000;
   35409: result <= 12'b111000000001;
   35410: result <= 12'b111000000001;
   35411: result <= 12'b111000000001;
   35412: result <= 12'b111000000001;
   35413: result <= 12'b111000000001;
   35414: result <= 12'b111000000001;
   35415: result <= 12'b111000000010;
   35416: result <= 12'b111000000010;
   35417: result <= 12'b111000000010;
   35418: result <= 12'b111000000010;
   35419: result <= 12'b111000000010;
   35420: result <= 12'b111000000011;
   35421: result <= 12'b111000000011;
   35422: result <= 12'b111000000011;
   35423: result <= 12'b111000000011;
   35424: result <= 12'b111000000011;
   35425: result <= 12'b111000000100;
   35426: result <= 12'b111000000100;
   35427: result <= 12'b111000000100;
   35428: result <= 12'b111000000100;
   35429: result <= 12'b111000000100;
   35430: result <= 12'b111000000101;
   35431: result <= 12'b111000000101;
   35432: result <= 12'b111000000101;
   35433: result <= 12'b111000000101;
   35434: result <= 12'b111000000101;
   35435: result <= 12'b111000000101;
   35436: result <= 12'b111000000110;
   35437: result <= 12'b111000000110;
   35438: result <= 12'b111000000110;
   35439: result <= 12'b111000000110;
   35440: result <= 12'b111000000110;
   35441: result <= 12'b111000000111;
   35442: result <= 12'b111000000111;
   35443: result <= 12'b111000000111;
   35444: result <= 12'b111000000111;
   35445: result <= 12'b111000000111;
   35446: result <= 12'b111000001000;
   35447: result <= 12'b111000001000;
   35448: result <= 12'b111000001000;
   35449: result <= 12'b111000001000;
   35450: result <= 12'b111000001000;
   35451: result <= 12'b111000001001;
   35452: result <= 12'b111000001001;
   35453: result <= 12'b111000001001;
   35454: result <= 12'b111000001001;
   35455: result <= 12'b111000001001;
   35456: result <= 12'b111000001001;
   35457: result <= 12'b111000001010;
   35458: result <= 12'b111000001010;
   35459: result <= 12'b111000001010;
   35460: result <= 12'b111000001010;
   35461: result <= 12'b111000001010;
   35462: result <= 12'b111000001011;
   35463: result <= 12'b111000001011;
   35464: result <= 12'b111000001011;
   35465: result <= 12'b111000001011;
   35466: result <= 12'b111000001011;
   35467: result <= 12'b111000001100;
   35468: result <= 12'b111000001100;
   35469: result <= 12'b111000001100;
   35470: result <= 12'b111000001100;
   35471: result <= 12'b111000001100;
   35472: result <= 12'b111000001101;
   35473: result <= 12'b111000001101;
   35474: result <= 12'b111000001101;
   35475: result <= 12'b111000001101;
   35476: result <= 12'b111000001101;
   35477: result <= 12'b111000001101;
   35478: result <= 12'b111000001110;
   35479: result <= 12'b111000001110;
   35480: result <= 12'b111000001110;
   35481: result <= 12'b111000001110;
   35482: result <= 12'b111000001110;
   35483: result <= 12'b111000001111;
   35484: result <= 12'b111000001111;
   35485: result <= 12'b111000001111;
   35486: result <= 12'b111000001111;
   35487: result <= 12'b111000001111;
   35488: result <= 12'b111000010000;
   35489: result <= 12'b111000010000;
   35490: result <= 12'b111000010000;
   35491: result <= 12'b111000010000;
   35492: result <= 12'b111000010000;
   35493: result <= 12'b111000010000;
   35494: result <= 12'b111000010001;
   35495: result <= 12'b111000010001;
   35496: result <= 12'b111000010001;
   35497: result <= 12'b111000010001;
   35498: result <= 12'b111000010001;
   35499: result <= 12'b111000010010;
   35500: result <= 12'b111000010010;
   35501: result <= 12'b111000010010;
   35502: result <= 12'b111000010010;
   35503: result <= 12'b111000010010;
   35504: result <= 12'b111000010011;
   35505: result <= 12'b111000010011;
   35506: result <= 12'b111000010011;
   35507: result <= 12'b111000010011;
   35508: result <= 12'b111000010011;
   35509: result <= 12'b111000010100;
   35510: result <= 12'b111000010100;
   35511: result <= 12'b111000010100;
   35512: result <= 12'b111000010100;
   35513: result <= 12'b111000010100;
   35514: result <= 12'b111000010100;
   35515: result <= 12'b111000010101;
   35516: result <= 12'b111000010101;
   35517: result <= 12'b111000010101;
   35518: result <= 12'b111000010101;
   35519: result <= 12'b111000010101;
   35520: result <= 12'b111000010110;
   35521: result <= 12'b111000010110;
   35522: result <= 12'b111000010110;
   35523: result <= 12'b111000010110;
   35524: result <= 12'b111000010110;
   35525: result <= 12'b111000010111;
   35526: result <= 12'b111000010111;
   35527: result <= 12'b111000010111;
   35528: result <= 12'b111000010111;
   35529: result <= 12'b111000010111;
   35530: result <= 12'b111000011000;
   35531: result <= 12'b111000011000;
   35532: result <= 12'b111000011000;
   35533: result <= 12'b111000011000;
   35534: result <= 12'b111000011000;
   35535: result <= 12'b111000011000;
   35536: result <= 12'b111000011001;
   35537: result <= 12'b111000011001;
   35538: result <= 12'b111000011001;
   35539: result <= 12'b111000011001;
   35540: result <= 12'b111000011001;
   35541: result <= 12'b111000011010;
   35542: result <= 12'b111000011010;
   35543: result <= 12'b111000011010;
   35544: result <= 12'b111000011010;
   35545: result <= 12'b111000011010;
   35546: result <= 12'b111000011011;
   35547: result <= 12'b111000011011;
   35548: result <= 12'b111000011011;
   35549: result <= 12'b111000011011;
   35550: result <= 12'b111000011011;
   35551: result <= 12'b111000011011;
   35552: result <= 12'b111000011100;
   35553: result <= 12'b111000011100;
   35554: result <= 12'b111000011100;
   35555: result <= 12'b111000011100;
   35556: result <= 12'b111000011100;
   35557: result <= 12'b111000011101;
   35558: result <= 12'b111000011101;
   35559: result <= 12'b111000011101;
   35560: result <= 12'b111000011101;
   35561: result <= 12'b111000011101;
   35562: result <= 12'b111000011110;
   35563: result <= 12'b111000011110;
   35564: result <= 12'b111000011110;
   35565: result <= 12'b111000011110;
   35566: result <= 12'b111000011110;
   35567: result <= 12'b111000011111;
   35568: result <= 12'b111000011111;
   35569: result <= 12'b111000011111;
   35570: result <= 12'b111000011111;
   35571: result <= 12'b111000011111;
   35572: result <= 12'b111000011111;
   35573: result <= 12'b111000100000;
   35574: result <= 12'b111000100000;
   35575: result <= 12'b111000100000;
   35576: result <= 12'b111000100000;
   35577: result <= 12'b111000100000;
   35578: result <= 12'b111000100001;
   35579: result <= 12'b111000100001;
   35580: result <= 12'b111000100001;
   35581: result <= 12'b111000100001;
   35582: result <= 12'b111000100001;
   35583: result <= 12'b111000100010;
   35584: result <= 12'b111000100010;
   35585: result <= 12'b111000100010;
   35586: result <= 12'b111000100010;
   35587: result <= 12'b111000100010;
   35588: result <= 12'b111000100010;
   35589: result <= 12'b111000100011;
   35590: result <= 12'b111000100011;
   35591: result <= 12'b111000100011;
   35592: result <= 12'b111000100011;
   35593: result <= 12'b111000100011;
   35594: result <= 12'b111000100100;
   35595: result <= 12'b111000100100;
   35596: result <= 12'b111000100100;
   35597: result <= 12'b111000100100;
   35598: result <= 12'b111000100100;
   35599: result <= 12'b111000100101;
   35600: result <= 12'b111000100101;
   35601: result <= 12'b111000100101;
   35602: result <= 12'b111000100101;
   35603: result <= 12'b111000100101;
   35604: result <= 12'b111000100110;
   35605: result <= 12'b111000100110;
   35606: result <= 12'b111000100110;
   35607: result <= 12'b111000100110;
   35608: result <= 12'b111000100110;
   35609: result <= 12'b111000100110;
   35610: result <= 12'b111000100111;
   35611: result <= 12'b111000100111;
   35612: result <= 12'b111000100111;
   35613: result <= 12'b111000100111;
   35614: result <= 12'b111000100111;
   35615: result <= 12'b111000101000;
   35616: result <= 12'b111000101000;
   35617: result <= 12'b111000101000;
   35618: result <= 12'b111000101000;
   35619: result <= 12'b111000101000;
   35620: result <= 12'b111000101001;
   35621: result <= 12'b111000101001;
   35622: result <= 12'b111000101001;
   35623: result <= 12'b111000101001;
   35624: result <= 12'b111000101001;
   35625: result <= 12'b111000101001;
   35626: result <= 12'b111000101010;
   35627: result <= 12'b111000101010;
   35628: result <= 12'b111000101010;
   35629: result <= 12'b111000101010;
   35630: result <= 12'b111000101010;
   35631: result <= 12'b111000101011;
   35632: result <= 12'b111000101011;
   35633: result <= 12'b111000101011;
   35634: result <= 12'b111000101011;
   35635: result <= 12'b111000101011;
   35636: result <= 12'b111000101100;
   35637: result <= 12'b111000101100;
   35638: result <= 12'b111000101100;
   35639: result <= 12'b111000101100;
   35640: result <= 12'b111000101100;
   35641: result <= 12'b111000101101;
   35642: result <= 12'b111000101101;
   35643: result <= 12'b111000101101;
   35644: result <= 12'b111000101101;
   35645: result <= 12'b111000101101;
   35646: result <= 12'b111000101101;
   35647: result <= 12'b111000101110;
   35648: result <= 12'b111000101110;
   35649: result <= 12'b111000101110;
   35650: result <= 12'b111000101110;
   35651: result <= 12'b111000101110;
   35652: result <= 12'b111000101111;
   35653: result <= 12'b111000101111;
   35654: result <= 12'b111000101111;
   35655: result <= 12'b111000101111;
   35656: result <= 12'b111000101111;
   35657: result <= 12'b111000110000;
   35658: result <= 12'b111000110000;
   35659: result <= 12'b111000110000;
   35660: result <= 12'b111000110000;
   35661: result <= 12'b111000110000;
   35662: result <= 12'b111000110000;
   35663: result <= 12'b111000110001;
   35664: result <= 12'b111000110001;
   35665: result <= 12'b111000110001;
   35666: result <= 12'b111000110001;
   35667: result <= 12'b111000110001;
   35668: result <= 12'b111000110010;
   35669: result <= 12'b111000110010;
   35670: result <= 12'b111000110010;
   35671: result <= 12'b111000110010;
   35672: result <= 12'b111000110010;
   35673: result <= 12'b111000110011;
   35674: result <= 12'b111000110011;
   35675: result <= 12'b111000110011;
   35676: result <= 12'b111000110011;
   35677: result <= 12'b111000110011;
   35678: result <= 12'b111000110011;
   35679: result <= 12'b111000110100;
   35680: result <= 12'b111000110100;
   35681: result <= 12'b111000110100;
   35682: result <= 12'b111000110100;
   35683: result <= 12'b111000110100;
   35684: result <= 12'b111000110101;
   35685: result <= 12'b111000110101;
   35686: result <= 12'b111000110101;
   35687: result <= 12'b111000110101;
   35688: result <= 12'b111000110101;
   35689: result <= 12'b111000110110;
   35690: result <= 12'b111000110110;
   35691: result <= 12'b111000110110;
   35692: result <= 12'b111000110110;
   35693: result <= 12'b111000110110;
   35694: result <= 12'b111000110111;
   35695: result <= 12'b111000110111;
   35696: result <= 12'b111000110111;
   35697: result <= 12'b111000110111;
   35698: result <= 12'b111000110111;
   35699: result <= 12'b111000110111;
   35700: result <= 12'b111000111000;
   35701: result <= 12'b111000111000;
   35702: result <= 12'b111000111000;
   35703: result <= 12'b111000111000;
   35704: result <= 12'b111000111000;
   35705: result <= 12'b111000111001;
   35706: result <= 12'b111000111001;
   35707: result <= 12'b111000111001;
   35708: result <= 12'b111000111001;
   35709: result <= 12'b111000111001;
   35710: result <= 12'b111000111010;
   35711: result <= 12'b111000111010;
   35712: result <= 12'b111000111010;
   35713: result <= 12'b111000111010;
   35714: result <= 12'b111000111010;
   35715: result <= 12'b111000111010;
   35716: result <= 12'b111000111011;
   35717: result <= 12'b111000111011;
   35718: result <= 12'b111000111011;
   35719: result <= 12'b111000111011;
   35720: result <= 12'b111000111011;
   35721: result <= 12'b111000111100;
   35722: result <= 12'b111000111100;
   35723: result <= 12'b111000111100;
   35724: result <= 12'b111000111100;
   35725: result <= 12'b111000111100;
   35726: result <= 12'b111000111101;
   35727: result <= 12'b111000111101;
   35728: result <= 12'b111000111101;
   35729: result <= 12'b111000111101;
   35730: result <= 12'b111000111101;
   35731: result <= 12'b111000111101;
   35732: result <= 12'b111000111110;
   35733: result <= 12'b111000111110;
   35734: result <= 12'b111000111110;
   35735: result <= 12'b111000111110;
   35736: result <= 12'b111000111110;
   35737: result <= 12'b111000111111;
   35738: result <= 12'b111000111111;
   35739: result <= 12'b111000111111;
   35740: result <= 12'b111000111111;
   35741: result <= 12'b111000111111;
   35742: result <= 12'b111001000000;
   35743: result <= 12'b111001000000;
   35744: result <= 12'b111001000000;
   35745: result <= 12'b111001000000;
   35746: result <= 12'b111001000000;
   35747: result <= 12'b111001000001;
   35748: result <= 12'b111001000001;
   35749: result <= 12'b111001000001;
   35750: result <= 12'b111001000001;
   35751: result <= 12'b111001000001;
   35752: result <= 12'b111001000001;
   35753: result <= 12'b111001000010;
   35754: result <= 12'b111001000010;
   35755: result <= 12'b111001000010;
   35756: result <= 12'b111001000010;
   35757: result <= 12'b111001000010;
   35758: result <= 12'b111001000011;
   35759: result <= 12'b111001000011;
   35760: result <= 12'b111001000011;
   35761: result <= 12'b111001000011;
   35762: result <= 12'b111001000011;
   35763: result <= 12'b111001000100;
   35764: result <= 12'b111001000100;
   35765: result <= 12'b111001000100;
   35766: result <= 12'b111001000100;
   35767: result <= 12'b111001000100;
   35768: result <= 12'b111001000100;
   35769: result <= 12'b111001000101;
   35770: result <= 12'b111001000101;
   35771: result <= 12'b111001000101;
   35772: result <= 12'b111001000101;
   35773: result <= 12'b111001000101;
   35774: result <= 12'b111001000110;
   35775: result <= 12'b111001000110;
   35776: result <= 12'b111001000110;
   35777: result <= 12'b111001000110;
   35778: result <= 12'b111001000110;
   35779: result <= 12'b111001000111;
   35780: result <= 12'b111001000111;
   35781: result <= 12'b111001000111;
   35782: result <= 12'b111001000111;
   35783: result <= 12'b111001000111;
   35784: result <= 12'b111001000111;
   35785: result <= 12'b111001001000;
   35786: result <= 12'b111001001000;
   35787: result <= 12'b111001001000;
   35788: result <= 12'b111001001000;
   35789: result <= 12'b111001001000;
   35790: result <= 12'b111001001001;
   35791: result <= 12'b111001001001;
   35792: result <= 12'b111001001001;
   35793: result <= 12'b111001001001;
   35794: result <= 12'b111001001001;
   35795: result <= 12'b111001001010;
   35796: result <= 12'b111001001010;
   35797: result <= 12'b111001001010;
   35798: result <= 12'b111001001010;
   35799: result <= 12'b111001001010;
   35800: result <= 12'b111001001010;
   35801: result <= 12'b111001001011;
   35802: result <= 12'b111001001011;
   35803: result <= 12'b111001001011;
   35804: result <= 12'b111001001011;
   35805: result <= 12'b111001001011;
   35806: result <= 12'b111001001100;
   35807: result <= 12'b111001001100;
   35808: result <= 12'b111001001100;
   35809: result <= 12'b111001001100;
   35810: result <= 12'b111001001100;
   35811: result <= 12'b111001001101;
   35812: result <= 12'b111001001101;
   35813: result <= 12'b111001001101;
   35814: result <= 12'b111001001101;
   35815: result <= 12'b111001001101;
   35816: result <= 12'b111001001101;
   35817: result <= 12'b111001001110;
   35818: result <= 12'b111001001110;
   35819: result <= 12'b111001001110;
   35820: result <= 12'b111001001110;
   35821: result <= 12'b111001001110;
   35822: result <= 12'b111001001111;
   35823: result <= 12'b111001001111;
   35824: result <= 12'b111001001111;
   35825: result <= 12'b111001001111;
   35826: result <= 12'b111001001111;
   35827: result <= 12'b111001010000;
   35828: result <= 12'b111001010000;
   35829: result <= 12'b111001010000;
   35830: result <= 12'b111001010000;
   35831: result <= 12'b111001010000;
   35832: result <= 12'b111001010000;
   35833: result <= 12'b111001010001;
   35834: result <= 12'b111001010001;
   35835: result <= 12'b111001010001;
   35836: result <= 12'b111001010001;
   35837: result <= 12'b111001010001;
   35838: result <= 12'b111001010010;
   35839: result <= 12'b111001010010;
   35840: result <= 12'b111001010010;
   35841: result <= 12'b111001010010;
   35842: result <= 12'b111001010010;
   35843: result <= 12'b111001010011;
   35844: result <= 12'b111001010011;
   35845: result <= 12'b111001010011;
   35846: result <= 12'b111001010011;
   35847: result <= 12'b111001010011;
   35848: result <= 12'b111001010100;
   35849: result <= 12'b111001010100;
   35850: result <= 12'b111001010100;
   35851: result <= 12'b111001010100;
   35852: result <= 12'b111001010100;
   35853: result <= 12'b111001010100;
   35854: result <= 12'b111001010101;
   35855: result <= 12'b111001010101;
   35856: result <= 12'b111001010101;
   35857: result <= 12'b111001010101;
   35858: result <= 12'b111001010101;
   35859: result <= 12'b111001010110;
   35860: result <= 12'b111001010110;
   35861: result <= 12'b111001010110;
   35862: result <= 12'b111001010110;
   35863: result <= 12'b111001010110;
   35864: result <= 12'b111001010111;
   35865: result <= 12'b111001010111;
   35866: result <= 12'b111001010111;
   35867: result <= 12'b111001010111;
   35868: result <= 12'b111001010111;
   35869: result <= 12'b111001010111;
   35870: result <= 12'b111001011000;
   35871: result <= 12'b111001011000;
   35872: result <= 12'b111001011000;
   35873: result <= 12'b111001011000;
   35874: result <= 12'b111001011000;
   35875: result <= 12'b111001011001;
   35876: result <= 12'b111001011001;
   35877: result <= 12'b111001011001;
   35878: result <= 12'b111001011001;
   35879: result <= 12'b111001011001;
   35880: result <= 12'b111001011010;
   35881: result <= 12'b111001011010;
   35882: result <= 12'b111001011010;
   35883: result <= 12'b111001011010;
   35884: result <= 12'b111001011010;
   35885: result <= 12'b111001011010;
   35886: result <= 12'b111001011011;
   35887: result <= 12'b111001011011;
   35888: result <= 12'b111001011011;
   35889: result <= 12'b111001011011;
   35890: result <= 12'b111001011011;
   35891: result <= 12'b111001011100;
   35892: result <= 12'b111001011100;
   35893: result <= 12'b111001011100;
   35894: result <= 12'b111001011100;
   35895: result <= 12'b111001011100;
   35896: result <= 12'b111001011101;
   35897: result <= 12'b111001011101;
   35898: result <= 12'b111001011101;
   35899: result <= 12'b111001011101;
   35900: result <= 12'b111001011101;
   35901: result <= 12'b111001011101;
   35902: result <= 12'b111001011110;
   35903: result <= 12'b111001011110;
   35904: result <= 12'b111001011110;
   35905: result <= 12'b111001011110;
   35906: result <= 12'b111001011110;
   35907: result <= 12'b111001011111;
   35908: result <= 12'b111001011111;
   35909: result <= 12'b111001011111;
   35910: result <= 12'b111001011111;
   35911: result <= 12'b111001011111;
   35912: result <= 12'b111001100000;
   35913: result <= 12'b111001100000;
   35914: result <= 12'b111001100000;
   35915: result <= 12'b111001100000;
   35916: result <= 12'b111001100000;
   35917: result <= 12'b111001100000;
   35918: result <= 12'b111001100001;
   35919: result <= 12'b111001100001;
   35920: result <= 12'b111001100001;
   35921: result <= 12'b111001100001;
   35922: result <= 12'b111001100001;
   35923: result <= 12'b111001100010;
   35924: result <= 12'b111001100010;
   35925: result <= 12'b111001100010;
   35926: result <= 12'b111001100010;
   35927: result <= 12'b111001100010;
   35928: result <= 12'b111001100011;
   35929: result <= 12'b111001100011;
   35930: result <= 12'b111001100011;
   35931: result <= 12'b111001100011;
   35932: result <= 12'b111001100011;
   35933: result <= 12'b111001100011;
   35934: result <= 12'b111001100100;
   35935: result <= 12'b111001100100;
   35936: result <= 12'b111001100100;
   35937: result <= 12'b111001100100;
   35938: result <= 12'b111001100100;
   35939: result <= 12'b111001100101;
   35940: result <= 12'b111001100101;
   35941: result <= 12'b111001100101;
   35942: result <= 12'b111001100101;
   35943: result <= 12'b111001100101;
   35944: result <= 12'b111001100110;
   35945: result <= 12'b111001100110;
   35946: result <= 12'b111001100110;
   35947: result <= 12'b111001100110;
   35948: result <= 12'b111001100110;
   35949: result <= 12'b111001100110;
   35950: result <= 12'b111001100111;
   35951: result <= 12'b111001100111;
   35952: result <= 12'b111001100111;
   35953: result <= 12'b111001100111;
   35954: result <= 12'b111001100111;
   35955: result <= 12'b111001101000;
   35956: result <= 12'b111001101000;
   35957: result <= 12'b111001101000;
   35958: result <= 12'b111001101000;
   35959: result <= 12'b111001101000;
   35960: result <= 12'b111001101001;
   35961: result <= 12'b111001101001;
   35962: result <= 12'b111001101001;
   35963: result <= 12'b111001101001;
   35964: result <= 12'b111001101001;
   35965: result <= 12'b111001101001;
   35966: result <= 12'b111001101010;
   35967: result <= 12'b111001101010;
   35968: result <= 12'b111001101010;
   35969: result <= 12'b111001101010;
   35970: result <= 12'b111001101010;
   35971: result <= 12'b111001101011;
   35972: result <= 12'b111001101011;
   35973: result <= 12'b111001101011;
   35974: result <= 12'b111001101011;
   35975: result <= 12'b111001101011;
   35976: result <= 12'b111001101100;
   35977: result <= 12'b111001101100;
   35978: result <= 12'b111001101100;
   35979: result <= 12'b111001101100;
   35980: result <= 12'b111001101100;
   35981: result <= 12'b111001101100;
   35982: result <= 12'b111001101101;
   35983: result <= 12'b111001101101;
   35984: result <= 12'b111001101101;
   35985: result <= 12'b111001101101;
   35986: result <= 12'b111001101101;
   35987: result <= 12'b111001101110;
   35988: result <= 12'b111001101110;
   35989: result <= 12'b111001101110;
   35990: result <= 12'b111001101110;
   35991: result <= 12'b111001101110;
   35992: result <= 12'b111001101110;
   35993: result <= 12'b111001101111;
   35994: result <= 12'b111001101111;
   35995: result <= 12'b111001101111;
   35996: result <= 12'b111001101111;
   35997: result <= 12'b111001101111;
   35998: result <= 12'b111001110000;
   35999: result <= 12'b111001110000;
   36000: result <= 12'b111001110000;
   36001: result <= 12'b111001110000;
   36002: result <= 12'b111001110000;
   36003: result <= 12'b111001110001;
   36004: result <= 12'b111001110001;
   36005: result <= 12'b111001110001;
   36006: result <= 12'b111001110001;
   36007: result <= 12'b111001110001;
   36008: result <= 12'b111001110001;
   36009: result <= 12'b111001110010;
   36010: result <= 12'b111001110010;
   36011: result <= 12'b111001110010;
   36012: result <= 12'b111001110010;
   36013: result <= 12'b111001110010;
   36014: result <= 12'b111001110011;
   36015: result <= 12'b111001110011;
   36016: result <= 12'b111001110011;
   36017: result <= 12'b111001110011;
   36018: result <= 12'b111001110011;
   36019: result <= 12'b111001110100;
   36020: result <= 12'b111001110100;
   36021: result <= 12'b111001110100;
   36022: result <= 12'b111001110100;
   36023: result <= 12'b111001110100;
   36024: result <= 12'b111001110100;
   36025: result <= 12'b111001110101;
   36026: result <= 12'b111001110101;
   36027: result <= 12'b111001110101;
   36028: result <= 12'b111001110101;
   36029: result <= 12'b111001110101;
   36030: result <= 12'b111001110110;
   36031: result <= 12'b111001110110;
   36032: result <= 12'b111001110110;
   36033: result <= 12'b111001110110;
   36034: result <= 12'b111001110110;
   36035: result <= 12'b111001110111;
   36036: result <= 12'b111001110111;
   36037: result <= 12'b111001110111;
   36038: result <= 12'b111001110111;
   36039: result <= 12'b111001110111;
   36040: result <= 12'b111001110111;
   36041: result <= 12'b111001111000;
   36042: result <= 12'b111001111000;
   36043: result <= 12'b111001111000;
   36044: result <= 12'b111001111000;
   36045: result <= 12'b111001111000;
   36046: result <= 12'b111001111001;
   36047: result <= 12'b111001111001;
   36048: result <= 12'b111001111001;
   36049: result <= 12'b111001111001;
   36050: result <= 12'b111001111001;
   36051: result <= 12'b111001111010;
   36052: result <= 12'b111001111010;
   36053: result <= 12'b111001111010;
   36054: result <= 12'b111001111010;
   36055: result <= 12'b111001111010;
   36056: result <= 12'b111001111010;
   36057: result <= 12'b111001111011;
   36058: result <= 12'b111001111011;
   36059: result <= 12'b111001111011;
   36060: result <= 12'b111001111011;
   36061: result <= 12'b111001111011;
   36062: result <= 12'b111001111100;
   36063: result <= 12'b111001111100;
   36064: result <= 12'b111001111100;
   36065: result <= 12'b111001111100;
   36066: result <= 12'b111001111100;
   36067: result <= 12'b111001111101;
   36068: result <= 12'b111001111101;
   36069: result <= 12'b111001111101;
   36070: result <= 12'b111001111101;
   36071: result <= 12'b111001111101;
   36072: result <= 12'b111001111101;
   36073: result <= 12'b111001111110;
   36074: result <= 12'b111001111110;
   36075: result <= 12'b111001111110;
   36076: result <= 12'b111001111110;
   36077: result <= 12'b111001111110;
   36078: result <= 12'b111001111111;
   36079: result <= 12'b111001111111;
   36080: result <= 12'b111001111111;
   36081: result <= 12'b111001111111;
   36082: result <= 12'b111001111111;
   36083: result <= 12'b111001111111;
   36084: result <= 12'b111010000000;
   36085: result <= 12'b111010000000;
   36086: result <= 12'b111010000000;
   36087: result <= 12'b111010000000;
   36088: result <= 12'b111010000000;
   36089: result <= 12'b111010000001;
   36090: result <= 12'b111010000001;
   36091: result <= 12'b111010000001;
   36092: result <= 12'b111010000001;
   36093: result <= 12'b111010000001;
   36094: result <= 12'b111010000010;
   36095: result <= 12'b111010000010;
   36096: result <= 12'b111010000010;
   36097: result <= 12'b111010000010;
   36098: result <= 12'b111010000010;
   36099: result <= 12'b111010000010;
   36100: result <= 12'b111010000011;
   36101: result <= 12'b111010000011;
   36102: result <= 12'b111010000011;
   36103: result <= 12'b111010000011;
   36104: result <= 12'b111010000011;
   36105: result <= 12'b111010000100;
   36106: result <= 12'b111010000100;
   36107: result <= 12'b111010000100;
   36108: result <= 12'b111010000100;
   36109: result <= 12'b111010000100;
   36110: result <= 12'b111010000101;
   36111: result <= 12'b111010000101;
   36112: result <= 12'b111010000101;
   36113: result <= 12'b111010000101;
   36114: result <= 12'b111010000101;
   36115: result <= 12'b111010000101;
   36116: result <= 12'b111010000110;
   36117: result <= 12'b111010000110;
   36118: result <= 12'b111010000110;
   36119: result <= 12'b111010000110;
   36120: result <= 12'b111010000110;
   36121: result <= 12'b111010000111;
   36122: result <= 12'b111010000111;
   36123: result <= 12'b111010000111;
   36124: result <= 12'b111010000111;
   36125: result <= 12'b111010000111;
   36126: result <= 12'b111010001000;
   36127: result <= 12'b111010001000;
   36128: result <= 12'b111010001000;
   36129: result <= 12'b111010001000;
   36130: result <= 12'b111010001000;
   36131: result <= 12'b111010001000;
   36132: result <= 12'b111010001001;
   36133: result <= 12'b111010001001;
   36134: result <= 12'b111010001001;
   36135: result <= 12'b111010001001;
   36136: result <= 12'b111010001001;
   36137: result <= 12'b111010001010;
   36138: result <= 12'b111010001010;
   36139: result <= 12'b111010001010;
   36140: result <= 12'b111010001010;
   36141: result <= 12'b111010001010;
   36142: result <= 12'b111010001010;
   36143: result <= 12'b111010001011;
   36144: result <= 12'b111010001011;
   36145: result <= 12'b111010001011;
   36146: result <= 12'b111010001011;
   36147: result <= 12'b111010001011;
   36148: result <= 12'b111010001100;
   36149: result <= 12'b111010001100;
   36150: result <= 12'b111010001100;
   36151: result <= 12'b111010001100;
   36152: result <= 12'b111010001100;
   36153: result <= 12'b111010001101;
   36154: result <= 12'b111010001101;
   36155: result <= 12'b111010001101;
   36156: result <= 12'b111010001101;
   36157: result <= 12'b111010001101;
   36158: result <= 12'b111010001101;
   36159: result <= 12'b111010001110;
   36160: result <= 12'b111010001110;
   36161: result <= 12'b111010001110;
   36162: result <= 12'b111010001110;
   36163: result <= 12'b111010001110;
   36164: result <= 12'b111010001111;
   36165: result <= 12'b111010001111;
   36166: result <= 12'b111010001111;
   36167: result <= 12'b111010001111;
   36168: result <= 12'b111010001111;
   36169: result <= 12'b111010010000;
   36170: result <= 12'b111010010000;
   36171: result <= 12'b111010010000;
   36172: result <= 12'b111010010000;
   36173: result <= 12'b111010010000;
   36174: result <= 12'b111010010000;
   36175: result <= 12'b111010010001;
   36176: result <= 12'b111010010001;
   36177: result <= 12'b111010010001;
   36178: result <= 12'b111010010001;
   36179: result <= 12'b111010010001;
   36180: result <= 12'b111010010010;
   36181: result <= 12'b111010010010;
   36182: result <= 12'b111010010010;
   36183: result <= 12'b111010010010;
   36184: result <= 12'b111010010010;
   36185: result <= 12'b111010010010;
   36186: result <= 12'b111010010011;
   36187: result <= 12'b111010010011;
   36188: result <= 12'b111010010011;
   36189: result <= 12'b111010010011;
   36190: result <= 12'b111010010011;
   36191: result <= 12'b111010010100;
   36192: result <= 12'b111010010100;
   36193: result <= 12'b111010010100;
   36194: result <= 12'b111010010100;
   36195: result <= 12'b111010010100;
   36196: result <= 12'b111010010101;
   36197: result <= 12'b111010010101;
   36198: result <= 12'b111010010101;
   36199: result <= 12'b111010010101;
   36200: result <= 12'b111010010101;
   36201: result <= 12'b111010010101;
   36202: result <= 12'b111010010110;
   36203: result <= 12'b111010010110;
   36204: result <= 12'b111010010110;
   36205: result <= 12'b111010010110;
   36206: result <= 12'b111010010110;
   36207: result <= 12'b111010010111;
   36208: result <= 12'b111010010111;
   36209: result <= 12'b111010010111;
   36210: result <= 12'b111010010111;
   36211: result <= 12'b111010010111;
   36212: result <= 12'b111010011000;
   36213: result <= 12'b111010011000;
   36214: result <= 12'b111010011000;
   36215: result <= 12'b111010011000;
   36216: result <= 12'b111010011000;
   36217: result <= 12'b111010011000;
   36218: result <= 12'b111010011001;
   36219: result <= 12'b111010011001;
   36220: result <= 12'b111010011001;
   36221: result <= 12'b111010011001;
   36222: result <= 12'b111010011001;
   36223: result <= 12'b111010011010;
   36224: result <= 12'b111010011010;
   36225: result <= 12'b111010011010;
   36226: result <= 12'b111010011010;
   36227: result <= 12'b111010011010;
   36228: result <= 12'b111010011010;
   36229: result <= 12'b111010011011;
   36230: result <= 12'b111010011011;
   36231: result <= 12'b111010011011;
   36232: result <= 12'b111010011011;
   36233: result <= 12'b111010011011;
   36234: result <= 12'b111010011100;
   36235: result <= 12'b111010011100;
   36236: result <= 12'b111010011100;
   36237: result <= 12'b111010011100;
   36238: result <= 12'b111010011100;
   36239: result <= 12'b111010011101;
   36240: result <= 12'b111010011101;
   36241: result <= 12'b111010011101;
   36242: result <= 12'b111010011101;
   36243: result <= 12'b111010011101;
   36244: result <= 12'b111010011101;
   36245: result <= 12'b111010011110;
   36246: result <= 12'b111010011110;
   36247: result <= 12'b111010011110;
   36248: result <= 12'b111010011110;
   36249: result <= 12'b111010011110;
   36250: result <= 12'b111010011111;
   36251: result <= 12'b111010011111;
   36252: result <= 12'b111010011111;
   36253: result <= 12'b111010011111;
   36254: result <= 12'b111010011111;
   36255: result <= 12'b111010011111;
   36256: result <= 12'b111010100000;
   36257: result <= 12'b111010100000;
   36258: result <= 12'b111010100000;
   36259: result <= 12'b111010100000;
   36260: result <= 12'b111010100000;
   36261: result <= 12'b111010100001;
   36262: result <= 12'b111010100001;
   36263: result <= 12'b111010100001;
   36264: result <= 12'b111010100001;
   36265: result <= 12'b111010100001;
   36266: result <= 12'b111010100010;
   36267: result <= 12'b111010100010;
   36268: result <= 12'b111010100010;
   36269: result <= 12'b111010100010;
   36270: result <= 12'b111010100010;
   36271: result <= 12'b111010100010;
   36272: result <= 12'b111010100011;
   36273: result <= 12'b111010100011;
   36274: result <= 12'b111010100011;
   36275: result <= 12'b111010100011;
   36276: result <= 12'b111010100011;
   36277: result <= 12'b111010100100;
   36278: result <= 12'b111010100100;
   36279: result <= 12'b111010100100;
   36280: result <= 12'b111010100100;
   36281: result <= 12'b111010100100;
   36282: result <= 12'b111010100100;
   36283: result <= 12'b111010100101;
   36284: result <= 12'b111010100101;
   36285: result <= 12'b111010100101;
   36286: result <= 12'b111010100101;
   36287: result <= 12'b111010100101;
   36288: result <= 12'b111010100110;
   36289: result <= 12'b111010100110;
   36290: result <= 12'b111010100110;
   36291: result <= 12'b111010100110;
   36292: result <= 12'b111010100110;
   36293: result <= 12'b111010100111;
   36294: result <= 12'b111010100111;
   36295: result <= 12'b111010100111;
   36296: result <= 12'b111010100111;
   36297: result <= 12'b111010100111;
   36298: result <= 12'b111010100111;
   36299: result <= 12'b111010101000;
   36300: result <= 12'b111010101000;
   36301: result <= 12'b111010101000;
   36302: result <= 12'b111010101000;
   36303: result <= 12'b111010101000;
   36304: result <= 12'b111010101001;
   36305: result <= 12'b111010101001;
   36306: result <= 12'b111010101001;
   36307: result <= 12'b111010101001;
   36308: result <= 12'b111010101001;
   36309: result <= 12'b111010101001;
   36310: result <= 12'b111010101010;
   36311: result <= 12'b111010101010;
   36312: result <= 12'b111010101010;
   36313: result <= 12'b111010101010;
   36314: result <= 12'b111010101010;
   36315: result <= 12'b111010101011;
   36316: result <= 12'b111010101011;
   36317: result <= 12'b111010101011;
   36318: result <= 12'b111010101011;
   36319: result <= 12'b111010101011;
   36320: result <= 12'b111010101100;
   36321: result <= 12'b111010101100;
   36322: result <= 12'b111010101100;
   36323: result <= 12'b111010101100;
   36324: result <= 12'b111010101100;
   36325: result <= 12'b111010101100;
   36326: result <= 12'b111010101101;
   36327: result <= 12'b111010101101;
   36328: result <= 12'b111010101101;
   36329: result <= 12'b111010101101;
   36330: result <= 12'b111010101101;
   36331: result <= 12'b111010101110;
   36332: result <= 12'b111010101110;
   36333: result <= 12'b111010101110;
   36334: result <= 12'b111010101110;
   36335: result <= 12'b111010101110;
   36336: result <= 12'b111010101110;
   36337: result <= 12'b111010101111;
   36338: result <= 12'b111010101111;
   36339: result <= 12'b111010101111;
   36340: result <= 12'b111010101111;
   36341: result <= 12'b111010101111;
   36342: result <= 12'b111010110000;
   36343: result <= 12'b111010110000;
   36344: result <= 12'b111010110000;
   36345: result <= 12'b111010110000;
   36346: result <= 12'b111010110000;
   36347: result <= 12'b111010110001;
   36348: result <= 12'b111010110001;
   36349: result <= 12'b111010110001;
   36350: result <= 12'b111010110001;
   36351: result <= 12'b111010110001;
   36352: result <= 12'b111010110001;
   36353: result <= 12'b111010110010;
   36354: result <= 12'b111010110010;
   36355: result <= 12'b111010110010;
   36356: result <= 12'b111010110010;
   36357: result <= 12'b111010110010;
   36358: result <= 12'b111010110011;
   36359: result <= 12'b111010110011;
   36360: result <= 12'b111010110011;
   36361: result <= 12'b111010110011;
   36362: result <= 12'b111010110011;
   36363: result <= 12'b111010110011;
   36364: result <= 12'b111010110100;
   36365: result <= 12'b111010110100;
   36366: result <= 12'b111010110100;
   36367: result <= 12'b111010110100;
   36368: result <= 12'b111010110100;
   36369: result <= 12'b111010110101;
   36370: result <= 12'b111010110101;
   36371: result <= 12'b111010110101;
   36372: result <= 12'b111010110101;
   36373: result <= 12'b111010110101;
   36374: result <= 12'b111010110110;
   36375: result <= 12'b111010110110;
   36376: result <= 12'b111010110110;
   36377: result <= 12'b111010110110;
   36378: result <= 12'b111010110110;
   36379: result <= 12'b111010110110;
   36380: result <= 12'b111010110111;
   36381: result <= 12'b111010110111;
   36382: result <= 12'b111010110111;
   36383: result <= 12'b111010110111;
   36384: result <= 12'b111010110111;
   36385: result <= 12'b111010111000;
   36386: result <= 12'b111010111000;
   36387: result <= 12'b111010111000;
   36388: result <= 12'b111010111000;
   36389: result <= 12'b111010111000;
   36390: result <= 12'b111010111000;
   36391: result <= 12'b111010111001;
   36392: result <= 12'b111010111001;
   36393: result <= 12'b111010111001;
   36394: result <= 12'b111010111001;
   36395: result <= 12'b111010111001;
   36396: result <= 12'b111010111010;
   36397: result <= 12'b111010111010;
   36398: result <= 12'b111010111010;
   36399: result <= 12'b111010111010;
   36400: result <= 12'b111010111010;
   36401: result <= 12'b111010111011;
   36402: result <= 12'b111010111011;
   36403: result <= 12'b111010111011;
   36404: result <= 12'b111010111011;
   36405: result <= 12'b111010111011;
   36406: result <= 12'b111010111011;
   36407: result <= 12'b111010111100;
   36408: result <= 12'b111010111100;
   36409: result <= 12'b111010111100;
   36410: result <= 12'b111010111100;
   36411: result <= 12'b111010111100;
   36412: result <= 12'b111010111101;
   36413: result <= 12'b111010111101;
   36414: result <= 12'b111010111101;
   36415: result <= 12'b111010111101;
   36416: result <= 12'b111010111101;
   36417: result <= 12'b111010111101;
   36418: result <= 12'b111010111110;
   36419: result <= 12'b111010111110;
   36420: result <= 12'b111010111110;
   36421: result <= 12'b111010111110;
   36422: result <= 12'b111010111110;
   36423: result <= 12'b111010111111;
   36424: result <= 12'b111010111111;
   36425: result <= 12'b111010111111;
   36426: result <= 12'b111010111111;
   36427: result <= 12'b111010111111;
   36428: result <= 12'b111010111111;
   36429: result <= 12'b111011000000;
   36430: result <= 12'b111011000000;
   36431: result <= 12'b111011000000;
   36432: result <= 12'b111011000000;
   36433: result <= 12'b111011000000;
   36434: result <= 12'b111011000001;
   36435: result <= 12'b111011000001;
   36436: result <= 12'b111011000001;
   36437: result <= 12'b111011000001;
   36438: result <= 12'b111011000001;
   36439: result <= 12'b111011000010;
   36440: result <= 12'b111011000010;
   36441: result <= 12'b111011000010;
   36442: result <= 12'b111011000010;
   36443: result <= 12'b111011000010;
   36444: result <= 12'b111011000010;
   36445: result <= 12'b111011000011;
   36446: result <= 12'b111011000011;
   36447: result <= 12'b111011000011;
   36448: result <= 12'b111011000011;
   36449: result <= 12'b111011000011;
   36450: result <= 12'b111011000100;
   36451: result <= 12'b111011000100;
   36452: result <= 12'b111011000100;
   36453: result <= 12'b111011000100;
   36454: result <= 12'b111011000100;
   36455: result <= 12'b111011000100;
   36456: result <= 12'b111011000101;
   36457: result <= 12'b111011000101;
   36458: result <= 12'b111011000101;
   36459: result <= 12'b111011000101;
   36460: result <= 12'b111011000101;
   36461: result <= 12'b111011000110;
   36462: result <= 12'b111011000110;
   36463: result <= 12'b111011000110;
   36464: result <= 12'b111011000110;
   36465: result <= 12'b111011000110;
   36466: result <= 12'b111011000110;
   36467: result <= 12'b111011000111;
   36468: result <= 12'b111011000111;
   36469: result <= 12'b111011000111;
   36470: result <= 12'b111011000111;
   36471: result <= 12'b111011000111;
   36472: result <= 12'b111011001000;
   36473: result <= 12'b111011001000;
   36474: result <= 12'b111011001000;
   36475: result <= 12'b111011001000;
   36476: result <= 12'b111011001000;
   36477: result <= 12'b111011001001;
   36478: result <= 12'b111011001001;
   36479: result <= 12'b111011001001;
   36480: result <= 12'b111011001001;
   36481: result <= 12'b111011001001;
   36482: result <= 12'b111011001001;
   36483: result <= 12'b111011001010;
   36484: result <= 12'b111011001010;
   36485: result <= 12'b111011001010;
   36486: result <= 12'b111011001010;
   36487: result <= 12'b111011001010;
   36488: result <= 12'b111011001011;
   36489: result <= 12'b111011001011;
   36490: result <= 12'b111011001011;
   36491: result <= 12'b111011001011;
   36492: result <= 12'b111011001011;
   36493: result <= 12'b111011001011;
   36494: result <= 12'b111011001100;
   36495: result <= 12'b111011001100;
   36496: result <= 12'b111011001100;
   36497: result <= 12'b111011001100;
   36498: result <= 12'b111011001100;
   36499: result <= 12'b111011001101;
   36500: result <= 12'b111011001101;
   36501: result <= 12'b111011001101;
   36502: result <= 12'b111011001101;
   36503: result <= 12'b111011001101;
   36504: result <= 12'b111011001101;
   36505: result <= 12'b111011001110;
   36506: result <= 12'b111011001110;
   36507: result <= 12'b111011001110;
   36508: result <= 12'b111011001110;
   36509: result <= 12'b111011001110;
   36510: result <= 12'b111011001111;
   36511: result <= 12'b111011001111;
   36512: result <= 12'b111011001111;
   36513: result <= 12'b111011001111;
   36514: result <= 12'b111011001111;
   36515: result <= 12'b111011001111;
   36516: result <= 12'b111011010000;
   36517: result <= 12'b111011010000;
   36518: result <= 12'b111011010000;
   36519: result <= 12'b111011010000;
   36520: result <= 12'b111011010000;
   36521: result <= 12'b111011010001;
   36522: result <= 12'b111011010001;
   36523: result <= 12'b111011010001;
   36524: result <= 12'b111011010001;
   36525: result <= 12'b111011010001;
   36526: result <= 12'b111011010010;
   36527: result <= 12'b111011010010;
   36528: result <= 12'b111011010010;
   36529: result <= 12'b111011010010;
   36530: result <= 12'b111011010010;
   36531: result <= 12'b111011010010;
   36532: result <= 12'b111011010011;
   36533: result <= 12'b111011010011;
   36534: result <= 12'b111011010011;
   36535: result <= 12'b111011010011;
   36536: result <= 12'b111011010011;
   36537: result <= 12'b111011010100;
   36538: result <= 12'b111011010100;
   36539: result <= 12'b111011010100;
   36540: result <= 12'b111011010100;
   36541: result <= 12'b111011010100;
   36542: result <= 12'b111011010100;
   36543: result <= 12'b111011010101;
   36544: result <= 12'b111011010101;
   36545: result <= 12'b111011010101;
   36546: result <= 12'b111011010101;
   36547: result <= 12'b111011010101;
   36548: result <= 12'b111011010110;
   36549: result <= 12'b111011010110;
   36550: result <= 12'b111011010110;
   36551: result <= 12'b111011010110;
   36552: result <= 12'b111011010110;
   36553: result <= 12'b111011010110;
   36554: result <= 12'b111011010111;
   36555: result <= 12'b111011010111;
   36556: result <= 12'b111011010111;
   36557: result <= 12'b111011010111;
   36558: result <= 12'b111011010111;
   36559: result <= 12'b111011011000;
   36560: result <= 12'b111011011000;
   36561: result <= 12'b111011011000;
   36562: result <= 12'b111011011000;
   36563: result <= 12'b111011011000;
   36564: result <= 12'b111011011000;
   36565: result <= 12'b111011011001;
   36566: result <= 12'b111011011001;
   36567: result <= 12'b111011011001;
   36568: result <= 12'b111011011001;
   36569: result <= 12'b111011011001;
   36570: result <= 12'b111011011010;
   36571: result <= 12'b111011011010;
   36572: result <= 12'b111011011010;
   36573: result <= 12'b111011011010;
   36574: result <= 12'b111011011010;
   36575: result <= 12'b111011011011;
   36576: result <= 12'b111011011011;
   36577: result <= 12'b111011011011;
   36578: result <= 12'b111011011011;
   36579: result <= 12'b111011011011;
   36580: result <= 12'b111011011011;
   36581: result <= 12'b111011011100;
   36582: result <= 12'b111011011100;
   36583: result <= 12'b111011011100;
   36584: result <= 12'b111011011100;
   36585: result <= 12'b111011011100;
   36586: result <= 12'b111011011101;
   36587: result <= 12'b111011011101;
   36588: result <= 12'b111011011101;
   36589: result <= 12'b111011011101;
   36590: result <= 12'b111011011101;
   36591: result <= 12'b111011011101;
   36592: result <= 12'b111011011110;
   36593: result <= 12'b111011011110;
   36594: result <= 12'b111011011110;
   36595: result <= 12'b111011011110;
   36596: result <= 12'b111011011110;
   36597: result <= 12'b111011011111;
   36598: result <= 12'b111011011111;
   36599: result <= 12'b111011011111;
   36600: result <= 12'b111011011111;
   36601: result <= 12'b111011011111;
   36602: result <= 12'b111011011111;
   36603: result <= 12'b111011100000;
   36604: result <= 12'b111011100000;
   36605: result <= 12'b111011100000;
   36606: result <= 12'b111011100000;
   36607: result <= 12'b111011100000;
   36608: result <= 12'b111011100001;
   36609: result <= 12'b111011100001;
   36610: result <= 12'b111011100001;
   36611: result <= 12'b111011100001;
   36612: result <= 12'b111011100001;
   36613: result <= 12'b111011100001;
   36614: result <= 12'b111011100010;
   36615: result <= 12'b111011100010;
   36616: result <= 12'b111011100010;
   36617: result <= 12'b111011100010;
   36618: result <= 12'b111011100010;
   36619: result <= 12'b111011100011;
   36620: result <= 12'b111011100011;
   36621: result <= 12'b111011100011;
   36622: result <= 12'b111011100011;
   36623: result <= 12'b111011100011;
   36624: result <= 12'b111011100011;
   36625: result <= 12'b111011100100;
   36626: result <= 12'b111011100100;
   36627: result <= 12'b111011100100;
   36628: result <= 12'b111011100100;
   36629: result <= 12'b111011100100;
   36630: result <= 12'b111011100101;
   36631: result <= 12'b111011100101;
   36632: result <= 12'b111011100101;
   36633: result <= 12'b111011100101;
   36634: result <= 12'b111011100101;
   36635: result <= 12'b111011100110;
   36636: result <= 12'b111011100110;
   36637: result <= 12'b111011100110;
   36638: result <= 12'b111011100110;
   36639: result <= 12'b111011100110;
   36640: result <= 12'b111011100110;
   36641: result <= 12'b111011100111;
   36642: result <= 12'b111011100111;
   36643: result <= 12'b111011100111;
   36644: result <= 12'b111011100111;
   36645: result <= 12'b111011100111;
   36646: result <= 12'b111011101000;
   36647: result <= 12'b111011101000;
   36648: result <= 12'b111011101000;
   36649: result <= 12'b111011101000;
   36650: result <= 12'b111011101000;
   36651: result <= 12'b111011101000;
   36652: result <= 12'b111011101001;
   36653: result <= 12'b111011101001;
   36654: result <= 12'b111011101001;
   36655: result <= 12'b111011101001;
   36656: result <= 12'b111011101001;
   36657: result <= 12'b111011101010;
   36658: result <= 12'b111011101010;
   36659: result <= 12'b111011101010;
   36660: result <= 12'b111011101010;
   36661: result <= 12'b111011101010;
   36662: result <= 12'b111011101010;
   36663: result <= 12'b111011101011;
   36664: result <= 12'b111011101011;
   36665: result <= 12'b111011101011;
   36666: result <= 12'b111011101011;
   36667: result <= 12'b111011101011;
   36668: result <= 12'b111011101100;
   36669: result <= 12'b111011101100;
   36670: result <= 12'b111011101100;
   36671: result <= 12'b111011101100;
   36672: result <= 12'b111011101100;
   36673: result <= 12'b111011101100;
   36674: result <= 12'b111011101101;
   36675: result <= 12'b111011101101;
   36676: result <= 12'b111011101101;
   36677: result <= 12'b111011101101;
   36678: result <= 12'b111011101101;
   36679: result <= 12'b111011101110;
   36680: result <= 12'b111011101110;
   36681: result <= 12'b111011101110;
   36682: result <= 12'b111011101110;
   36683: result <= 12'b111011101110;
   36684: result <= 12'b111011101110;
   36685: result <= 12'b111011101111;
   36686: result <= 12'b111011101111;
   36687: result <= 12'b111011101111;
   36688: result <= 12'b111011101111;
   36689: result <= 12'b111011101111;
   36690: result <= 12'b111011110000;
   36691: result <= 12'b111011110000;
   36692: result <= 12'b111011110000;
   36693: result <= 12'b111011110000;
   36694: result <= 12'b111011110000;
   36695: result <= 12'b111011110000;
   36696: result <= 12'b111011110001;
   36697: result <= 12'b111011110001;
   36698: result <= 12'b111011110001;
   36699: result <= 12'b111011110001;
   36700: result <= 12'b111011110001;
   36701: result <= 12'b111011110010;
   36702: result <= 12'b111011110010;
   36703: result <= 12'b111011110010;
   36704: result <= 12'b111011110010;
   36705: result <= 12'b111011110010;
   36706: result <= 12'b111011110010;
   36707: result <= 12'b111011110011;
   36708: result <= 12'b111011110011;
   36709: result <= 12'b111011110011;
   36710: result <= 12'b111011110011;
   36711: result <= 12'b111011110011;
   36712: result <= 12'b111011110100;
   36713: result <= 12'b111011110100;
   36714: result <= 12'b111011110100;
   36715: result <= 12'b111011110100;
   36716: result <= 12'b111011110100;
   36717: result <= 12'b111011110100;
   36718: result <= 12'b111011110101;
   36719: result <= 12'b111011110101;
   36720: result <= 12'b111011110101;
   36721: result <= 12'b111011110101;
   36722: result <= 12'b111011110101;
   36723: result <= 12'b111011110110;
   36724: result <= 12'b111011110110;
   36725: result <= 12'b111011110110;
   36726: result <= 12'b111011110110;
   36727: result <= 12'b111011110110;
   36728: result <= 12'b111011110110;
   36729: result <= 12'b111011110111;
   36730: result <= 12'b111011110111;
   36731: result <= 12'b111011110111;
   36732: result <= 12'b111011110111;
   36733: result <= 12'b111011110111;
   36734: result <= 12'b111011111000;
   36735: result <= 12'b111011111000;
   36736: result <= 12'b111011111000;
   36737: result <= 12'b111011111000;
   36738: result <= 12'b111011111000;
   36739: result <= 12'b111011111001;
   36740: result <= 12'b111011111001;
   36741: result <= 12'b111011111001;
   36742: result <= 12'b111011111001;
   36743: result <= 12'b111011111001;
   36744: result <= 12'b111011111001;
   36745: result <= 12'b111011111010;
   36746: result <= 12'b111011111010;
   36747: result <= 12'b111011111010;
   36748: result <= 12'b111011111010;
   36749: result <= 12'b111011111010;
   36750: result <= 12'b111011111011;
   36751: result <= 12'b111011111011;
   36752: result <= 12'b111011111011;
   36753: result <= 12'b111011111011;
   36754: result <= 12'b111011111011;
   36755: result <= 12'b111011111011;
   36756: result <= 12'b111011111100;
   36757: result <= 12'b111011111100;
   36758: result <= 12'b111011111100;
   36759: result <= 12'b111011111100;
   36760: result <= 12'b111011111100;
   36761: result <= 12'b111011111101;
   36762: result <= 12'b111011111101;
   36763: result <= 12'b111011111101;
   36764: result <= 12'b111011111101;
   36765: result <= 12'b111011111101;
   36766: result <= 12'b111011111101;
   36767: result <= 12'b111011111110;
   36768: result <= 12'b111011111110;
   36769: result <= 12'b111011111110;
   36770: result <= 12'b111011111110;
   36771: result <= 12'b111011111110;
   36772: result <= 12'b111011111111;
   36773: result <= 12'b111011111111;
   36774: result <= 12'b111011111111;
   36775: result <= 12'b111011111111;
   36776: result <= 12'b111011111111;
   36777: result <= 12'b111011111111;
   36778: result <= 12'b111100000000;
   36779: result <= 12'b111100000000;
   36780: result <= 12'b111100000000;
   36781: result <= 12'b111100000000;
   36782: result <= 12'b111100000000;
   36783: result <= 12'b111100000001;
   36784: result <= 12'b111100000001;
   36785: result <= 12'b111100000001;
   36786: result <= 12'b111100000001;
   36787: result <= 12'b111100000001;
   36788: result <= 12'b111100000001;
   36789: result <= 12'b111100000010;
   36790: result <= 12'b111100000010;
   36791: result <= 12'b111100000010;
   36792: result <= 12'b111100000010;
   36793: result <= 12'b111100000010;
   36794: result <= 12'b111100000011;
   36795: result <= 12'b111100000011;
   36796: result <= 12'b111100000011;
   36797: result <= 12'b111100000011;
   36798: result <= 12'b111100000011;
   36799: result <= 12'b111100000011;
   36800: result <= 12'b111100000100;
   36801: result <= 12'b111100000100;
   36802: result <= 12'b111100000100;
   36803: result <= 12'b111100000100;
   36804: result <= 12'b111100000100;
   36805: result <= 12'b111100000101;
   36806: result <= 12'b111100000101;
   36807: result <= 12'b111100000101;
   36808: result <= 12'b111100000101;
   36809: result <= 12'b111100000101;
   36810: result <= 12'b111100000101;
   36811: result <= 12'b111100000110;
   36812: result <= 12'b111100000110;
   36813: result <= 12'b111100000110;
   36814: result <= 12'b111100000110;
   36815: result <= 12'b111100000110;
   36816: result <= 12'b111100000111;
   36817: result <= 12'b111100000111;
   36818: result <= 12'b111100000111;
   36819: result <= 12'b111100000111;
   36820: result <= 12'b111100000111;
   36821: result <= 12'b111100000111;
   36822: result <= 12'b111100001000;
   36823: result <= 12'b111100001000;
   36824: result <= 12'b111100001000;
   36825: result <= 12'b111100001000;
   36826: result <= 12'b111100001000;
   36827: result <= 12'b111100001001;
   36828: result <= 12'b111100001001;
   36829: result <= 12'b111100001001;
   36830: result <= 12'b111100001001;
   36831: result <= 12'b111100001001;
   36832: result <= 12'b111100001001;
   36833: result <= 12'b111100001010;
   36834: result <= 12'b111100001010;
   36835: result <= 12'b111100001010;
   36836: result <= 12'b111100001010;
   36837: result <= 12'b111100001010;
   36838: result <= 12'b111100001011;
   36839: result <= 12'b111100001011;
   36840: result <= 12'b111100001011;
   36841: result <= 12'b111100001011;
   36842: result <= 12'b111100001011;
   36843: result <= 12'b111100001011;
   36844: result <= 12'b111100001100;
   36845: result <= 12'b111100001100;
   36846: result <= 12'b111100001100;
   36847: result <= 12'b111100001100;
   36848: result <= 12'b111100001100;
   36849: result <= 12'b111100001101;
   36850: result <= 12'b111100001101;
   36851: result <= 12'b111100001101;
   36852: result <= 12'b111100001101;
   36853: result <= 12'b111100001101;
   36854: result <= 12'b111100001101;
   36855: result <= 12'b111100001110;
   36856: result <= 12'b111100001110;
   36857: result <= 12'b111100001110;
   36858: result <= 12'b111100001110;
   36859: result <= 12'b111100001110;
   36860: result <= 12'b111100001111;
   36861: result <= 12'b111100001111;
   36862: result <= 12'b111100001111;
   36863: result <= 12'b111100001111;
   36864: result <= 12'b111100001111;
   36865: result <= 12'b111100001111;
   36866: result <= 12'b111100010000;
   36867: result <= 12'b111100010000;
   36868: result <= 12'b111100010000;
   36869: result <= 12'b111100010000;
   36870: result <= 12'b111100010000;
   36871: result <= 12'b111100010001;
   36872: result <= 12'b111100010001;
   36873: result <= 12'b111100010001;
   36874: result <= 12'b111100010001;
   36875: result <= 12'b111100010001;
   36876: result <= 12'b111100010001;
   36877: result <= 12'b111100010010;
   36878: result <= 12'b111100010010;
   36879: result <= 12'b111100010010;
   36880: result <= 12'b111100010010;
   36881: result <= 12'b111100010010;
   36882: result <= 12'b111100010010;
   36883: result <= 12'b111100010011;
   36884: result <= 12'b111100010011;
   36885: result <= 12'b111100010011;
   36886: result <= 12'b111100010011;
   36887: result <= 12'b111100010011;
   36888: result <= 12'b111100010100;
   36889: result <= 12'b111100010100;
   36890: result <= 12'b111100010100;
   36891: result <= 12'b111100010100;
   36892: result <= 12'b111100010100;
   36893: result <= 12'b111100010100;
   36894: result <= 12'b111100010101;
   36895: result <= 12'b111100010101;
   36896: result <= 12'b111100010101;
   36897: result <= 12'b111100010101;
   36898: result <= 12'b111100010101;
   36899: result <= 12'b111100010110;
   36900: result <= 12'b111100010110;
   36901: result <= 12'b111100010110;
   36902: result <= 12'b111100010110;
   36903: result <= 12'b111100010110;
   36904: result <= 12'b111100010110;
   36905: result <= 12'b111100010111;
   36906: result <= 12'b111100010111;
   36907: result <= 12'b111100010111;
   36908: result <= 12'b111100010111;
   36909: result <= 12'b111100010111;
   36910: result <= 12'b111100011000;
   36911: result <= 12'b111100011000;
   36912: result <= 12'b111100011000;
   36913: result <= 12'b111100011000;
   36914: result <= 12'b111100011000;
   36915: result <= 12'b111100011000;
   36916: result <= 12'b111100011001;
   36917: result <= 12'b111100011001;
   36918: result <= 12'b111100011001;
   36919: result <= 12'b111100011001;
   36920: result <= 12'b111100011001;
   36921: result <= 12'b111100011010;
   36922: result <= 12'b111100011010;
   36923: result <= 12'b111100011010;
   36924: result <= 12'b111100011010;
   36925: result <= 12'b111100011010;
   36926: result <= 12'b111100011010;
   36927: result <= 12'b111100011011;
   36928: result <= 12'b111100011011;
   36929: result <= 12'b111100011011;
   36930: result <= 12'b111100011011;
   36931: result <= 12'b111100011011;
   36932: result <= 12'b111100011100;
   36933: result <= 12'b111100011100;
   36934: result <= 12'b111100011100;
   36935: result <= 12'b111100011100;
   36936: result <= 12'b111100011100;
   36937: result <= 12'b111100011100;
   36938: result <= 12'b111100011101;
   36939: result <= 12'b111100011101;
   36940: result <= 12'b111100011101;
   36941: result <= 12'b111100011101;
   36942: result <= 12'b111100011101;
   36943: result <= 12'b111100011110;
   36944: result <= 12'b111100011110;
   36945: result <= 12'b111100011110;
   36946: result <= 12'b111100011110;
   36947: result <= 12'b111100011110;
   36948: result <= 12'b111100011110;
   36949: result <= 12'b111100011111;
   36950: result <= 12'b111100011111;
   36951: result <= 12'b111100011111;
   36952: result <= 12'b111100011111;
   36953: result <= 12'b111100011111;
   36954: result <= 12'b111100100000;
   36955: result <= 12'b111100100000;
   36956: result <= 12'b111100100000;
   36957: result <= 12'b111100100000;
   36958: result <= 12'b111100100000;
   36959: result <= 12'b111100100000;
   36960: result <= 12'b111100100001;
   36961: result <= 12'b111100100001;
   36962: result <= 12'b111100100001;
   36963: result <= 12'b111100100001;
   36964: result <= 12'b111100100001;
   36965: result <= 12'b111100100010;
   36966: result <= 12'b111100100010;
   36967: result <= 12'b111100100010;
   36968: result <= 12'b111100100010;
   36969: result <= 12'b111100100010;
   36970: result <= 12'b111100100010;
   36971: result <= 12'b111100100011;
   36972: result <= 12'b111100100011;
   36973: result <= 12'b111100100011;
   36974: result <= 12'b111100100011;
   36975: result <= 12'b111100100011;
   36976: result <= 12'b111100100100;
   36977: result <= 12'b111100100100;
   36978: result <= 12'b111100100100;
   36979: result <= 12'b111100100100;
   36980: result <= 12'b111100100100;
   36981: result <= 12'b111100100100;
   36982: result <= 12'b111100100101;
   36983: result <= 12'b111100100101;
   36984: result <= 12'b111100100101;
   36985: result <= 12'b111100100101;
   36986: result <= 12'b111100100101;
   36987: result <= 12'b111100100101;
   36988: result <= 12'b111100100110;
   36989: result <= 12'b111100100110;
   36990: result <= 12'b111100100110;
   36991: result <= 12'b111100100110;
   36992: result <= 12'b111100100110;
   36993: result <= 12'b111100100111;
   36994: result <= 12'b111100100111;
   36995: result <= 12'b111100100111;
   36996: result <= 12'b111100100111;
   36997: result <= 12'b111100100111;
   36998: result <= 12'b111100100111;
   36999: result <= 12'b111100101000;
   37000: result <= 12'b111100101000;
   37001: result <= 12'b111100101000;
   37002: result <= 12'b111100101000;
   37003: result <= 12'b111100101000;
   37004: result <= 12'b111100101001;
   37005: result <= 12'b111100101001;
   37006: result <= 12'b111100101001;
   37007: result <= 12'b111100101001;
   37008: result <= 12'b111100101001;
   37009: result <= 12'b111100101001;
   37010: result <= 12'b111100101010;
   37011: result <= 12'b111100101010;
   37012: result <= 12'b111100101010;
   37013: result <= 12'b111100101010;
   37014: result <= 12'b111100101010;
   37015: result <= 12'b111100101011;
   37016: result <= 12'b111100101011;
   37017: result <= 12'b111100101011;
   37018: result <= 12'b111100101011;
   37019: result <= 12'b111100101011;
   37020: result <= 12'b111100101011;
   37021: result <= 12'b111100101100;
   37022: result <= 12'b111100101100;
   37023: result <= 12'b111100101100;
   37024: result <= 12'b111100101100;
   37025: result <= 12'b111100101100;
   37026: result <= 12'b111100101101;
   37027: result <= 12'b111100101101;
   37028: result <= 12'b111100101101;
   37029: result <= 12'b111100101101;
   37030: result <= 12'b111100101101;
   37031: result <= 12'b111100101101;
   37032: result <= 12'b111100101110;
   37033: result <= 12'b111100101110;
   37034: result <= 12'b111100101110;
   37035: result <= 12'b111100101110;
   37036: result <= 12'b111100101110;
   37037: result <= 12'b111100101111;
   37038: result <= 12'b111100101111;
   37039: result <= 12'b111100101111;
   37040: result <= 12'b111100101111;
   37041: result <= 12'b111100101111;
   37042: result <= 12'b111100101111;
   37043: result <= 12'b111100110000;
   37044: result <= 12'b111100110000;
   37045: result <= 12'b111100110000;
   37046: result <= 12'b111100110000;
   37047: result <= 12'b111100110000;
   37048: result <= 12'b111100110000;
   37049: result <= 12'b111100110001;
   37050: result <= 12'b111100110001;
   37051: result <= 12'b111100110001;
   37052: result <= 12'b111100110001;
   37053: result <= 12'b111100110001;
   37054: result <= 12'b111100110010;
   37055: result <= 12'b111100110010;
   37056: result <= 12'b111100110010;
   37057: result <= 12'b111100110010;
   37058: result <= 12'b111100110010;
   37059: result <= 12'b111100110010;
   37060: result <= 12'b111100110011;
   37061: result <= 12'b111100110011;
   37062: result <= 12'b111100110011;
   37063: result <= 12'b111100110011;
   37064: result <= 12'b111100110011;
   37065: result <= 12'b111100110100;
   37066: result <= 12'b111100110100;
   37067: result <= 12'b111100110100;
   37068: result <= 12'b111100110100;
   37069: result <= 12'b111100110100;
   37070: result <= 12'b111100110100;
   37071: result <= 12'b111100110101;
   37072: result <= 12'b111100110101;
   37073: result <= 12'b111100110101;
   37074: result <= 12'b111100110101;
   37075: result <= 12'b111100110101;
   37076: result <= 12'b111100110110;
   37077: result <= 12'b111100110110;
   37078: result <= 12'b111100110110;
   37079: result <= 12'b111100110110;
   37080: result <= 12'b111100110110;
   37081: result <= 12'b111100110110;
   37082: result <= 12'b111100110111;
   37083: result <= 12'b111100110111;
   37084: result <= 12'b111100110111;
   37085: result <= 12'b111100110111;
   37086: result <= 12'b111100110111;
   37087: result <= 12'b111100111000;
   37088: result <= 12'b111100111000;
   37089: result <= 12'b111100111000;
   37090: result <= 12'b111100111000;
   37091: result <= 12'b111100111000;
   37092: result <= 12'b111100111000;
   37093: result <= 12'b111100111001;
   37094: result <= 12'b111100111001;
   37095: result <= 12'b111100111001;
   37096: result <= 12'b111100111001;
   37097: result <= 12'b111100111001;
   37098: result <= 12'b111100111001;
   37099: result <= 12'b111100111010;
   37100: result <= 12'b111100111010;
   37101: result <= 12'b111100111010;
   37102: result <= 12'b111100111010;
   37103: result <= 12'b111100111010;
   37104: result <= 12'b111100111011;
   37105: result <= 12'b111100111011;
   37106: result <= 12'b111100111011;
   37107: result <= 12'b111100111011;
   37108: result <= 12'b111100111011;
   37109: result <= 12'b111100111011;
   37110: result <= 12'b111100111100;
   37111: result <= 12'b111100111100;
   37112: result <= 12'b111100111100;
   37113: result <= 12'b111100111100;
   37114: result <= 12'b111100111100;
   37115: result <= 12'b111100111101;
   37116: result <= 12'b111100111101;
   37117: result <= 12'b111100111101;
   37118: result <= 12'b111100111101;
   37119: result <= 12'b111100111101;
   37120: result <= 12'b111100111101;
   37121: result <= 12'b111100111110;
   37122: result <= 12'b111100111110;
   37123: result <= 12'b111100111110;
   37124: result <= 12'b111100111110;
   37125: result <= 12'b111100111110;
   37126: result <= 12'b111100111111;
   37127: result <= 12'b111100111111;
   37128: result <= 12'b111100111111;
   37129: result <= 12'b111100111111;
   37130: result <= 12'b111100111111;
   37131: result <= 12'b111100111111;
   37132: result <= 12'b111101000000;
   37133: result <= 12'b111101000000;
   37134: result <= 12'b111101000000;
   37135: result <= 12'b111101000000;
   37136: result <= 12'b111101000000;
   37137: result <= 12'b111101000000;
   37138: result <= 12'b111101000001;
   37139: result <= 12'b111101000001;
   37140: result <= 12'b111101000001;
   37141: result <= 12'b111101000001;
   37142: result <= 12'b111101000001;
   37143: result <= 12'b111101000010;
   37144: result <= 12'b111101000010;
   37145: result <= 12'b111101000010;
   37146: result <= 12'b111101000010;
   37147: result <= 12'b111101000010;
   37148: result <= 12'b111101000010;
   37149: result <= 12'b111101000011;
   37150: result <= 12'b111101000011;
   37151: result <= 12'b111101000011;
   37152: result <= 12'b111101000011;
   37153: result <= 12'b111101000011;
   37154: result <= 12'b111101000100;
   37155: result <= 12'b111101000100;
   37156: result <= 12'b111101000100;
   37157: result <= 12'b111101000100;
   37158: result <= 12'b111101000100;
   37159: result <= 12'b111101000100;
   37160: result <= 12'b111101000101;
   37161: result <= 12'b111101000101;
   37162: result <= 12'b111101000101;
   37163: result <= 12'b111101000101;
   37164: result <= 12'b111101000101;
   37165: result <= 12'b111101000110;
   37166: result <= 12'b111101000110;
   37167: result <= 12'b111101000110;
   37168: result <= 12'b111101000110;
   37169: result <= 12'b111101000110;
   37170: result <= 12'b111101000110;
   37171: result <= 12'b111101000111;
   37172: result <= 12'b111101000111;
   37173: result <= 12'b111101000111;
   37174: result <= 12'b111101000111;
   37175: result <= 12'b111101000111;
   37176: result <= 12'b111101000111;
   37177: result <= 12'b111101001000;
   37178: result <= 12'b111101001000;
   37179: result <= 12'b111101001000;
   37180: result <= 12'b111101001000;
   37181: result <= 12'b111101001000;
   37182: result <= 12'b111101001001;
   37183: result <= 12'b111101001001;
   37184: result <= 12'b111101001001;
   37185: result <= 12'b111101001001;
   37186: result <= 12'b111101001001;
   37187: result <= 12'b111101001001;
   37188: result <= 12'b111101001010;
   37189: result <= 12'b111101001010;
   37190: result <= 12'b111101001010;
   37191: result <= 12'b111101001010;
   37192: result <= 12'b111101001010;
   37193: result <= 12'b111101001011;
   37194: result <= 12'b111101001011;
   37195: result <= 12'b111101001011;
   37196: result <= 12'b111101001011;
   37197: result <= 12'b111101001011;
   37198: result <= 12'b111101001011;
   37199: result <= 12'b111101001100;
   37200: result <= 12'b111101001100;
   37201: result <= 12'b111101001100;
   37202: result <= 12'b111101001100;
   37203: result <= 12'b111101001100;
   37204: result <= 12'b111101001100;
   37205: result <= 12'b111101001101;
   37206: result <= 12'b111101001101;
   37207: result <= 12'b111101001101;
   37208: result <= 12'b111101001101;
   37209: result <= 12'b111101001101;
   37210: result <= 12'b111101001110;
   37211: result <= 12'b111101001110;
   37212: result <= 12'b111101001110;
   37213: result <= 12'b111101001110;
   37214: result <= 12'b111101001110;
   37215: result <= 12'b111101001110;
   37216: result <= 12'b111101001111;
   37217: result <= 12'b111101001111;
   37218: result <= 12'b111101001111;
   37219: result <= 12'b111101001111;
   37220: result <= 12'b111101001111;
   37221: result <= 12'b111101010000;
   37222: result <= 12'b111101010000;
   37223: result <= 12'b111101010000;
   37224: result <= 12'b111101010000;
   37225: result <= 12'b111101010000;
   37226: result <= 12'b111101010000;
   37227: result <= 12'b111101010001;
   37228: result <= 12'b111101010001;
   37229: result <= 12'b111101010001;
   37230: result <= 12'b111101010001;
   37231: result <= 12'b111101010001;
   37232: result <= 12'b111101010001;
   37233: result <= 12'b111101010010;
   37234: result <= 12'b111101010010;
   37235: result <= 12'b111101010010;
   37236: result <= 12'b111101010010;
   37237: result <= 12'b111101010010;
   37238: result <= 12'b111101010011;
   37239: result <= 12'b111101010011;
   37240: result <= 12'b111101010011;
   37241: result <= 12'b111101010011;
   37242: result <= 12'b111101010011;
   37243: result <= 12'b111101010011;
   37244: result <= 12'b111101010100;
   37245: result <= 12'b111101010100;
   37246: result <= 12'b111101010100;
   37247: result <= 12'b111101010100;
   37248: result <= 12'b111101010100;
   37249: result <= 12'b111101010101;
   37250: result <= 12'b111101010101;
   37251: result <= 12'b111101010101;
   37252: result <= 12'b111101010101;
   37253: result <= 12'b111101010101;
   37254: result <= 12'b111101010101;
   37255: result <= 12'b111101010110;
   37256: result <= 12'b111101010110;
   37257: result <= 12'b111101010110;
   37258: result <= 12'b111101010110;
   37259: result <= 12'b111101010110;
   37260: result <= 12'b111101010110;
   37261: result <= 12'b111101010111;
   37262: result <= 12'b111101010111;
   37263: result <= 12'b111101010111;
   37264: result <= 12'b111101010111;
   37265: result <= 12'b111101010111;
   37266: result <= 12'b111101011000;
   37267: result <= 12'b111101011000;
   37268: result <= 12'b111101011000;
   37269: result <= 12'b111101011000;
   37270: result <= 12'b111101011000;
   37271: result <= 12'b111101011000;
   37272: result <= 12'b111101011001;
   37273: result <= 12'b111101011001;
   37274: result <= 12'b111101011001;
   37275: result <= 12'b111101011001;
   37276: result <= 12'b111101011001;
   37277: result <= 12'b111101011010;
   37278: result <= 12'b111101011010;
   37279: result <= 12'b111101011010;
   37280: result <= 12'b111101011010;
   37281: result <= 12'b111101011010;
   37282: result <= 12'b111101011010;
   37283: result <= 12'b111101011011;
   37284: result <= 12'b111101011011;
   37285: result <= 12'b111101011011;
   37286: result <= 12'b111101011011;
   37287: result <= 12'b111101011011;
   37288: result <= 12'b111101011011;
   37289: result <= 12'b111101011100;
   37290: result <= 12'b111101011100;
   37291: result <= 12'b111101011100;
   37292: result <= 12'b111101011100;
   37293: result <= 12'b111101011100;
   37294: result <= 12'b111101011101;
   37295: result <= 12'b111101011101;
   37296: result <= 12'b111101011101;
   37297: result <= 12'b111101011101;
   37298: result <= 12'b111101011101;
   37299: result <= 12'b111101011101;
   37300: result <= 12'b111101011110;
   37301: result <= 12'b111101011110;
   37302: result <= 12'b111101011110;
   37303: result <= 12'b111101011110;
   37304: result <= 12'b111101011110;
   37305: result <= 12'b111101011111;
   37306: result <= 12'b111101011111;
   37307: result <= 12'b111101011111;
   37308: result <= 12'b111101011111;
   37309: result <= 12'b111101011111;
   37310: result <= 12'b111101011111;
   37311: result <= 12'b111101100000;
   37312: result <= 12'b111101100000;
   37313: result <= 12'b111101100000;
   37314: result <= 12'b111101100000;
   37315: result <= 12'b111101100000;
   37316: result <= 12'b111101100000;
   37317: result <= 12'b111101100001;
   37318: result <= 12'b111101100001;
   37319: result <= 12'b111101100001;
   37320: result <= 12'b111101100001;
   37321: result <= 12'b111101100001;
   37322: result <= 12'b111101100010;
   37323: result <= 12'b111101100010;
   37324: result <= 12'b111101100010;
   37325: result <= 12'b111101100010;
   37326: result <= 12'b111101100010;
   37327: result <= 12'b111101100010;
   37328: result <= 12'b111101100011;
   37329: result <= 12'b111101100011;
   37330: result <= 12'b111101100011;
   37331: result <= 12'b111101100011;
   37332: result <= 12'b111101100011;
   37333: result <= 12'b111101100011;
   37334: result <= 12'b111101100100;
   37335: result <= 12'b111101100100;
   37336: result <= 12'b111101100100;
   37337: result <= 12'b111101100100;
   37338: result <= 12'b111101100100;
   37339: result <= 12'b111101100101;
   37340: result <= 12'b111101100101;
   37341: result <= 12'b111101100101;
   37342: result <= 12'b111101100101;
   37343: result <= 12'b111101100101;
   37344: result <= 12'b111101100101;
   37345: result <= 12'b111101100110;
   37346: result <= 12'b111101100110;
   37347: result <= 12'b111101100110;
   37348: result <= 12'b111101100110;
   37349: result <= 12'b111101100110;
   37350: result <= 12'b111101100111;
   37351: result <= 12'b111101100111;
   37352: result <= 12'b111101100111;
   37353: result <= 12'b111101100111;
   37354: result <= 12'b111101100111;
   37355: result <= 12'b111101100111;
   37356: result <= 12'b111101101000;
   37357: result <= 12'b111101101000;
   37358: result <= 12'b111101101000;
   37359: result <= 12'b111101101000;
   37360: result <= 12'b111101101000;
   37361: result <= 12'b111101101000;
   37362: result <= 12'b111101101001;
   37363: result <= 12'b111101101001;
   37364: result <= 12'b111101101001;
   37365: result <= 12'b111101101001;
   37366: result <= 12'b111101101001;
   37367: result <= 12'b111101101010;
   37368: result <= 12'b111101101010;
   37369: result <= 12'b111101101010;
   37370: result <= 12'b111101101010;
   37371: result <= 12'b111101101010;
   37372: result <= 12'b111101101010;
   37373: result <= 12'b111101101011;
   37374: result <= 12'b111101101011;
   37375: result <= 12'b111101101011;
   37376: result <= 12'b111101101011;
   37377: result <= 12'b111101101011;
   37378: result <= 12'b111101101011;
   37379: result <= 12'b111101101100;
   37380: result <= 12'b111101101100;
   37381: result <= 12'b111101101100;
   37382: result <= 12'b111101101100;
   37383: result <= 12'b111101101100;
   37384: result <= 12'b111101101101;
   37385: result <= 12'b111101101101;
   37386: result <= 12'b111101101101;
   37387: result <= 12'b111101101101;
   37388: result <= 12'b111101101101;
   37389: result <= 12'b111101101101;
   37390: result <= 12'b111101101110;
   37391: result <= 12'b111101101110;
   37392: result <= 12'b111101101110;
   37393: result <= 12'b111101101110;
   37394: result <= 12'b111101101110;
   37395: result <= 12'b111101101111;
   37396: result <= 12'b111101101111;
   37397: result <= 12'b111101101111;
   37398: result <= 12'b111101101111;
   37399: result <= 12'b111101101111;
   37400: result <= 12'b111101101111;
   37401: result <= 12'b111101110000;
   37402: result <= 12'b111101110000;
   37403: result <= 12'b111101110000;
   37404: result <= 12'b111101110000;
   37405: result <= 12'b111101110000;
   37406: result <= 12'b111101110000;
   37407: result <= 12'b111101110001;
   37408: result <= 12'b111101110001;
   37409: result <= 12'b111101110001;
   37410: result <= 12'b111101110001;
   37411: result <= 12'b111101110001;
   37412: result <= 12'b111101110010;
   37413: result <= 12'b111101110010;
   37414: result <= 12'b111101110010;
   37415: result <= 12'b111101110010;
   37416: result <= 12'b111101110010;
   37417: result <= 12'b111101110010;
   37418: result <= 12'b111101110011;
   37419: result <= 12'b111101110011;
   37420: result <= 12'b111101110011;
   37421: result <= 12'b111101110011;
   37422: result <= 12'b111101110011;
   37423: result <= 12'b111101110011;
   37424: result <= 12'b111101110100;
   37425: result <= 12'b111101110100;
   37426: result <= 12'b111101110100;
   37427: result <= 12'b111101110100;
   37428: result <= 12'b111101110100;
   37429: result <= 12'b111101110101;
   37430: result <= 12'b111101110101;
   37431: result <= 12'b111101110101;
   37432: result <= 12'b111101110101;
   37433: result <= 12'b111101110101;
   37434: result <= 12'b111101110101;
   37435: result <= 12'b111101110110;
   37436: result <= 12'b111101110110;
   37437: result <= 12'b111101110110;
   37438: result <= 12'b111101110110;
   37439: result <= 12'b111101110110;
   37440: result <= 12'b111101110110;
   37441: result <= 12'b111101110111;
   37442: result <= 12'b111101110111;
   37443: result <= 12'b111101110111;
   37444: result <= 12'b111101110111;
   37445: result <= 12'b111101110111;
   37446: result <= 12'b111101111000;
   37447: result <= 12'b111101111000;
   37448: result <= 12'b111101111000;
   37449: result <= 12'b111101111000;
   37450: result <= 12'b111101111000;
   37451: result <= 12'b111101111000;
   37452: result <= 12'b111101111001;
   37453: result <= 12'b111101111001;
   37454: result <= 12'b111101111001;
   37455: result <= 12'b111101111001;
   37456: result <= 12'b111101111001;
   37457: result <= 12'b111101111001;
   37458: result <= 12'b111101111010;
   37459: result <= 12'b111101111010;
   37460: result <= 12'b111101111010;
   37461: result <= 12'b111101111010;
   37462: result <= 12'b111101111010;
   37463: result <= 12'b111101111011;
   37464: result <= 12'b111101111011;
   37465: result <= 12'b111101111011;
   37466: result <= 12'b111101111011;
   37467: result <= 12'b111101111011;
   37468: result <= 12'b111101111011;
   37469: result <= 12'b111101111100;
   37470: result <= 12'b111101111100;
   37471: result <= 12'b111101111100;
   37472: result <= 12'b111101111100;
   37473: result <= 12'b111101111100;
   37474: result <= 12'b111101111100;
   37475: result <= 12'b111101111101;
   37476: result <= 12'b111101111101;
   37477: result <= 12'b111101111101;
   37478: result <= 12'b111101111101;
   37479: result <= 12'b111101111101;
   37480: result <= 12'b111101111110;
   37481: result <= 12'b111101111110;
   37482: result <= 12'b111101111110;
   37483: result <= 12'b111101111110;
   37484: result <= 12'b111101111110;
   37485: result <= 12'b111101111110;
   37486: result <= 12'b111101111111;
   37487: result <= 12'b111101111111;
   37488: result <= 12'b111101111111;
   37489: result <= 12'b111101111111;
   37490: result <= 12'b111101111111;
   37491: result <= 12'b111101111111;
   37492: result <= 12'b111110000000;
   37493: result <= 12'b111110000000;
   37494: result <= 12'b111110000000;
   37495: result <= 12'b111110000000;
   37496: result <= 12'b111110000000;
   37497: result <= 12'b111110000001;
   37498: result <= 12'b111110000001;
   37499: result <= 12'b111110000001;
   37500: result <= 12'b111110000001;
   37501: result <= 12'b111110000001;
   37502: result <= 12'b111110000001;
   37503: result <= 12'b111110000010;
   37504: result <= 12'b111110000010;
   37505: result <= 12'b111110000010;
   37506: result <= 12'b111110000010;
   37507: result <= 12'b111110000010;
   37508: result <= 12'b111110000010;
   37509: result <= 12'b111110000011;
   37510: result <= 12'b111110000011;
   37511: result <= 12'b111110000011;
   37512: result <= 12'b111110000011;
   37513: result <= 12'b111110000011;
   37514: result <= 12'b111110000100;
   37515: result <= 12'b111110000100;
   37516: result <= 12'b111110000100;
   37517: result <= 12'b111110000100;
   37518: result <= 12'b111110000100;
   37519: result <= 12'b111110000100;
   37520: result <= 12'b111110000101;
   37521: result <= 12'b111110000101;
   37522: result <= 12'b111110000101;
   37523: result <= 12'b111110000101;
   37524: result <= 12'b111110000101;
   37525: result <= 12'b111110000101;
   37526: result <= 12'b111110000110;
   37527: result <= 12'b111110000110;
   37528: result <= 12'b111110000110;
   37529: result <= 12'b111110000110;
   37530: result <= 12'b111110000110;
   37531: result <= 12'b111110000111;
   37532: result <= 12'b111110000111;
   37533: result <= 12'b111110000111;
   37534: result <= 12'b111110000111;
   37535: result <= 12'b111110000111;
   37536: result <= 12'b111110000111;
   37537: result <= 12'b111110001000;
   37538: result <= 12'b111110001000;
   37539: result <= 12'b111110001000;
   37540: result <= 12'b111110001000;
   37541: result <= 12'b111110001000;
   37542: result <= 12'b111110001000;
   37543: result <= 12'b111110001001;
   37544: result <= 12'b111110001001;
   37545: result <= 12'b111110001001;
   37546: result <= 12'b111110001001;
   37547: result <= 12'b111110001001;
   37548: result <= 12'b111110001010;
   37549: result <= 12'b111110001010;
   37550: result <= 12'b111110001010;
   37551: result <= 12'b111110001010;
   37552: result <= 12'b111110001010;
   37553: result <= 12'b111110001010;
   37554: result <= 12'b111110001011;
   37555: result <= 12'b111110001011;
   37556: result <= 12'b111110001011;
   37557: result <= 12'b111110001011;
   37558: result <= 12'b111110001011;
   37559: result <= 12'b111110001011;
   37560: result <= 12'b111110001100;
   37561: result <= 12'b111110001100;
   37562: result <= 12'b111110001100;
   37563: result <= 12'b111110001100;
   37564: result <= 12'b111110001100;
   37565: result <= 12'b111110001101;
   37566: result <= 12'b111110001101;
   37567: result <= 12'b111110001101;
   37568: result <= 12'b111110001101;
   37569: result <= 12'b111110001101;
   37570: result <= 12'b111110001101;
   37571: result <= 12'b111110001110;
   37572: result <= 12'b111110001110;
   37573: result <= 12'b111110001110;
   37574: result <= 12'b111110001110;
   37575: result <= 12'b111110001110;
   37576: result <= 12'b111110001110;
   37577: result <= 12'b111110001111;
   37578: result <= 12'b111110001111;
   37579: result <= 12'b111110001111;
   37580: result <= 12'b111110001111;
   37581: result <= 12'b111110001111;
   37582: result <= 12'b111110010000;
   37583: result <= 12'b111110010000;
   37584: result <= 12'b111110010000;
   37585: result <= 12'b111110010000;
   37586: result <= 12'b111110010000;
   37587: result <= 12'b111110010000;
   37588: result <= 12'b111110010001;
   37589: result <= 12'b111110010001;
   37590: result <= 12'b111110010001;
   37591: result <= 12'b111110010001;
   37592: result <= 12'b111110010001;
   37593: result <= 12'b111110010001;
   37594: result <= 12'b111110010010;
   37595: result <= 12'b111110010010;
   37596: result <= 12'b111110010010;
   37597: result <= 12'b111110010010;
   37598: result <= 12'b111110010010;
   37599: result <= 12'b111110010011;
   37600: result <= 12'b111110010011;
   37601: result <= 12'b111110010011;
   37602: result <= 12'b111110010011;
   37603: result <= 12'b111110010011;
   37604: result <= 12'b111110010011;
   37605: result <= 12'b111110010100;
   37606: result <= 12'b111110010100;
   37607: result <= 12'b111110010100;
   37608: result <= 12'b111110010100;
   37609: result <= 12'b111110010100;
   37610: result <= 12'b111110010100;
   37611: result <= 12'b111110010101;
   37612: result <= 12'b111110010101;
   37613: result <= 12'b111110010101;
   37614: result <= 12'b111110010101;
   37615: result <= 12'b111110010101;
   37616: result <= 12'b111110010101;
   37617: result <= 12'b111110010110;
   37618: result <= 12'b111110010110;
   37619: result <= 12'b111110010110;
   37620: result <= 12'b111110010110;
   37621: result <= 12'b111110010110;
   37622: result <= 12'b111110010111;
   37623: result <= 12'b111110010111;
   37624: result <= 12'b111110010111;
   37625: result <= 12'b111110010111;
   37626: result <= 12'b111110010111;
   37627: result <= 12'b111110010111;
   37628: result <= 12'b111110011000;
   37629: result <= 12'b111110011000;
   37630: result <= 12'b111110011000;
   37631: result <= 12'b111110011000;
   37632: result <= 12'b111110011000;
   37633: result <= 12'b111110011000;
   37634: result <= 12'b111110011001;
   37635: result <= 12'b111110011001;
   37636: result <= 12'b111110011001;
   37637: result <= 12'b111110011001;
   37638: result <= 12'b111110011001;
   37639: result <= 12'b111110011010;
   37640: result <= 12'b111110011010;
   37641: result <= 12'b111110011010;
   37642: result <= 12'b111110011010;
   37643: result <= 12'b111110011010;
   37644: result <= 12'b111110011010;
   37645: result <= 12'b111110011011;
   37646: result <= 12'b111110011011;
   37647: result <= 12'b111110011011;
   37648: result <= 12'b111110011011;
   37649: result <= 12'b111110011011;
   37650: result <= 12'b111110011011;
   37651: result <= 12'b111110011100;
   37652: result <= 12'b111110011100;
   37653: result <= 12'b111110011100;
   37654: result <= 12'b111110011100;
   37655: result <= 12'b111110011100;
   37656: result <= 12'b111110011101;
   37657: result <= 12'b111110011101;
   37658: result <= 12'b111110011101;
   37659: result <= 12'b111110011101;
   37660: result <= 12'b111110011101;
   37661: result <= 12'b111110011101;
   37662: result <= 12'b111110011110;
   37663: result <= 12'b111110011110;
   37664: result <= 12'b111110011110;
   37665: result <= 12'b111110011110;
   37666: result <= 12'b111110011110;
   37667: result <= 12'b111110011110;
   37668: result <= 12'b111110011111;
   37669: result <= 12'b111110011111;
   37670: result <= 12'b111110011111;
   37671: result <= 12'b111110011111;
   37672: result <= 12'b111110011111;
   37673: result <= 12'b111110011111;
   37674: result <= 12'b111110100000;
   37675: result <= 12'b111110100000;
   37676: result <= 12'b111110100000;
   37677: result <= 12'b111110100000;
   37678: result <= 12'b111110100000;
   37679: result <= 12'b111110100001;
   37680: result <= 12'b111110100001;
   37681: result <= 12'b111110100001;
   37682: result <= 12'b111110100001;
   37683: result <= 12'b111110100001;
   37684: result <= 12'b111110100001;
   37685: result <= 12'b111110100010;
   37686: result <= 12'b111110100010;
   37687: result <= 12'b111110100010;
   37688: result <= 12'b111110100010;
   37689: result <= 12'b111110100010;
   37690: result <= 12'b111110100010;
   37691: result <= 12'b111110100011;
   37692: result <= 12'b111110100011;
   37693: result <= 12'b111110100011;
   37694: result <= 12'b111110100011;
   37695: result <= 12'b111110100011;
   37696: result <= 12'b111110100100;
   37697: result <= 12'b111110100100;
   37698: result <= 12'b111110100100;
   37699: result <= 12'b111110100100;
   37700: result <= 12'b111110100100;
   37701: result <= 12'b111110100100;
   37702: result <= 12'b111110100101;
   37703: result <= 12'b111110100101;
   37704: result <= 12'b111110100101;
   37705: result <= 12'b111110100101;
   37706: result <= 12'b111110100101;
   37707: result <= 12'b111110100101;
   37708: result <= 12'b111110100110;
   37709: result <= 12'b111110100110;
   37710: result <= 12'b111110100110;
   37711: result <= 12'b111110100110;
   37712: result <= 12'b111110100110;
   37713: result <= 12'b111110100110;
   37714: result <= 12'b111110100111;
   37715: result <= 12'b111110100111;
   37716: result <= 12'b111110100111;
   37717: result <= 12'b111110100111;
   37718: result <= 12'b111110100111;
   37719: result <= 12'b111110101000;
   37720: result <= 12'b111110101000;
   37721: result <= 12'b111110101000;
   37722: result <= 12'b111110101000;
   37723: result <= 12'b111110101000;
   37724: result <= 12'b111110101000;
   37725: result <= 12'b111110101001;
   37726: result <= 12'b111110101001;
   37727: result <= 12'b111110101001;
   37728: result <= 12'b111110101001;
   37729: result <= 12'b111110101001;
   37730: result <= 12'b111110101001;
   37731: result <= 12'b111110101010;
   37732: result <= 12'b111110101010;
   37733: result <= 12'b111110101010;
   37734: result <= 12'b111110101010;
   37735: result <= 12'b111110101010;
   37736: result <= 12'b111110101010;
   37737: result <= 12'b111110101011;
   37738: result <= 12'b111110101011;
   37739: result <= 12'b111110101011;
   37740: result <= 12'b111110101011;
   37741: result <= 12'b111110101011;
   37742: result <= 12'b111110101100;
   37743: result <= 12'b111110101100;
   37744: result <= 12'b111110101100;
   37745: result <= 12'b111110101100;
   37746: result <= 12'b111110101100;
   37747: result <= 12'b111110101100;
   37748: result <= 12'b111110101101;
   37749: result <= 12'b111110101101;
   37750: result <= 12'b111110101101;
   37751: result <= 12'b111110101101;
   37752: result <= 12'b111110101101;
   37753: result <= 12'b111110101101;
   37754: result <= 12'b111110101110;
   37755: result <= 12'b111110101110;
   37756: result <= 12'b111110101110;
   37757: result <= 12'b111110101110;
   37758: result <= 12'b111110101110;
   37759: result <= 12'b111110101111;
   37760: result <= 12'b111110101111;
   37761: result <= 12'b111110101111;
   37762: result <= 12'b111110101111;
   37763: result <= 12'b111110101111;
   37764: result <= 12'b111110101111;
   37765: result <= 12'b111110110000;
   37766: result <= 12'b111110110000;
   37767: result <= 12'b111110110000;
   37768: result <= 12'b111110110000;
   37769: result <= 12'b111110110000;
   37770: result <= 12'b111110110000;
   37771: result <= 12'b111110110001;
   37772: result <= 12'b111110110001;
   37773: result <= 12'b111110110001;
   37774: result <= 12'b111110110001;
   37775: result <= 12'b111110110001;
   37776: result <= 12'b111110110001;
   37777: result <= 12'b111110110010;
   37778: result <= 12'b111110110010;
   37779: result <= 12'b111110110010;
   37780: result <= 12'b111110110010;
   37781: result <= 12'b111110110010;
   37782: result <= 12'b111110110011;
   37783: result <= 12'b111110110011;
   37784: result <= 12'b111110110011;
   37785: result <= 12'b111110110011;
   37786: result <= 12'b111110110011;
   37787: result <= 12'b111110110011;
   37788: result <= 12'b111110110100;
   37789: result <= 12'b111110110100;
   37790: result <= 12'b111110110100;
   37791: result <= 12'b111110110100;
   37792: result <= 12'b111110110100;
   37793: result <= 12'b111110110100;
   37794: result <= 12'b111110110101;
   37795: result <= 12'b111110110101;
   37796: result <= 12'b111110110101;
   37797: result <= 12'b111110110101;
   37798: result <= 12'b111110110101;
   37799: result <= 12'b111110110101;
   37800: result <= 12'b111110110110;
   37801: result <= 12'b111110110110;
   37802: result <= 12'b111110110110;
   37803: result <= 12'b111110110110;
   37804: result <= 12'b111110110110;
   37805: result <= 12'b111110110111;
   37806: result <= 12'b111110110111;
   37807: result <= 12'b111110110111;
   37808: result <= 12'b111110110111;
   37809: result <= 12'b111110110111;
   37810: result <= 12'b111110110111;
   37811: result <= 12'b111110111000;
   37812: result <= 12'b111110111000;
   37813: result <= 12'b111110111000;
   37814: result <= 12'b111110111000;
   37815: result <= 12'b111110111000;
   37816: result <= 12'b111110111000;
   37817: result <= 12'b111110111001;
   37818: result <= 12'b111110111001;
   37819: result <= 12'b111110111001;
   37820: result <= 12'b111110111001;
   37821: result <= 12'b111110111001;
   37822: result <= 12'b111110111001;
   37823: result <= 12'b111110111010;
   37824: result <= 12'b111110111010;
   37825: result <= 12'b111110111010;
   37826: result <= 12'b111110111010;
   37827: result <= 12'b111110111010;
   37828: result <= 12'b111110111011;
   37829: result <= 12'b111110111011;
   37830: result <= 12'b111110111011;
   37831: result <= 12'b111110111011;
   37832: result <= 12'b111110111011;
   37833: result <= 12'b111110111011;
   37834: result <= 12'b111110111100;
   37835: result <= 12'b111110111100;
   37836: result <= 12'b111110111100;
   37837: result <= 12'b111110111100;
   37838: result <= 12'b111110111100;
   37839: result <= 12'b111110111100;
   37840: result <= 12'b111110111101;
   37841: result <= 12'b111110111101;
   37842: result <= 12'b111110111101;
   37843: result <= 12'b111110111101;
   37844: result <= 12'b111110111101;
   37845: result <= 12'b111110111101;
   37846: result <= 12'b111110111110;
   37847: result <= 12'b111110111110;
   37848: result <= 12'b111110111110;
   37849: result <= 12'b111110111110;
   37850: result <= 12'b111110111110;
   37851: result <= 12'b111110111111;
   37852: result <= 12'b111110111111;
   37853: result <= 12'b111110111111;
   37854: result <= 12'b111110111111;
   37855: result <= 12'b111110111111;
   37856: result <= 12'b111110111111;
   37857: result <= 12'b111111000000;
   37858: result <= 12'b111111000000;
   37859: result <= 12'b111111000000;
   37860: result <= 12'b111111000000;
   37861: result <= 12'b111111000000;
   37862: result <= 12'b111111000000;
   37863: result <= 12'b111111000001;
   37864: result <= 12'b111111000001;
   37865: result <= 12'b111111000001;
   37866: result <= 12'b111111000001;
   37867: result <= 12'b111111000001;
   37868: result <= 12'b111111000001;
   37869: result <= 12'b111111000010;
   37870: result <= 12'b111111000010;
   37871: result <= 12'b111111000010;
   37872: result <= 12'b111111000010;
   37873: result <= 12'b111111000010;
   37874: result <= 12'b111111000010;
   37875: result <= 12'b111111000011;
   37876: result <= 12'b111111000011;
   37877: result <= 12'b111111000011;
   37878: result <= 12'b111111000011;
   37879: result <= 12'b111111000011;
   37880: result <= 12'b111111000100;
   37881: result <= 12'b111111000100;
   37882: result <= 12'b111111000100;
   37883: result <= 12'b111111000100;
   37884: result <= 12'b111111000100;
   37885: result <= 12'b111111000100;
   37886: result <= 12'b111111000101;
   37887: result <= 12'b111111000101;
   37888: result <= 12'b111111000101;
   37889: result <= 12'b111111000101;
   37890: result <= 12'b111111000101;
   37891: result <= 12'b111111000101;
   37892: result <= 12'b111111000110;
   37893: result <= 12'b111111000110;
   37894: result <= 12'b111111000110;
   37895: result <= 12'b111111000110;
   37896: result <= 12'b111111000110;
   37897: result <= 12'b111111000110;
   37898: result <= 12'b111111000111;
   37899: result <= 12'b111111000111;
   37900: result <= 12'b111111000111;
   37901: result <= 12'b111111000111;
   37902: result <= 12'b111111000111;
   37903: result <= 12'b111111001000;
   37904: result <= 12'b111111001000;
   37905: result <= 12'b111111001000;
   37906: result <= 12'b111111001000;
   37907: result <= 12'b111111001000;
   37908: result <= 12'b111111001000;
   37909: result <= 12'b111111001001;
   37910: result <= 12'b111111001001;
   37911: result <= 12'b111111001001;
   37912: result <= 12'b111111001001;
   37913: result <= 12'b111111001001;
   37914: result <= 12'b111111001001;
   37915: result <= 12'b111111001010;
   37916: result <= 12'b111111001010;
   37917: result <= 12'b111111001010;
   37918: result <= 12'b111111001010;
   37919: result <= 12'b111111001010;
   37920: result <= 12'b111111001010;
   37921: result <= 12'b111111001011;
   37922: result <= 12'b111111001011;
   37923: result <= 12'b111111001011;
   37924: result <= 12'b111111001011;
   37925: result <= 12'b111111001011;
   37926: result <= 12'b111111001011;
   37927: result <= 12'b111111001100;
   37928: result <= 12'b111111001100;
   37929: result <= 12'b111111001100;
   37930: result <= 12'b111111001100;
   37931: result <= 12'b111111001100;
   37932: result <= 12'b111111001101;
   37933: result <= 12'b111111001101;
   37934: result <= 12'b111111001101;
   37935: result <= 12'b111111001101;
   37936: result <= 12'b111111001101;
   37937: result <= 12'b111111001101;
   37938: result <= 12'b111111001110;
   37939: result <= 12'b111111001110;
   37940: result <= 12'b111111001110;
   37941: result <= 12'b111111001110;
   37942: result <= 12'b111111001110;
   37943: result <= 12'b111111001110;
   37944: result <= 12'b111111001111;
   37945: result <= 12'b111111001111;
   37946: result <= 12'b111111001111;
   37947: result <= 12'b111111001111;
   37948: result <= 12'b111111001111;
   37949: result <= 12'b111111001111;
   37950: result <= 12'b111111010000;
   37951: result <= 12'b111111010000;
   37952: result <= 12'b111111010000;
   37953: result <= 12'b111111010000;
   37954: result <= 12'b111111010000;
   37955: result <= 12'b111111010001;
   37956: result <= 12'b111111010001;
   37957: result <= 12'b111111010001;
   37958: result <= 12'b111111010001;
   37959: result <= 12'b111111010001;
   37960: result <= 12'b111111010001;
   37961: result <= 12'b111111010010;
   37962: result <= 12'b111111010010;
   37963: result <= 12'b111111010010;
   37964: result <= 12'b111111010010;
   37965: result <= 12'b111111010010;
   37966: result <= 12'b111111010010;
   37967: result <= 12'b111111010011;
   37968: result <= 12'b111111010011;
   37969: result <= 12'b111111010011;
   37970: result <= 12'b111111010011;
   37971: result <= 12'b111111010011;
   37972: result <= 12'b111111010011;
   37973: result <= 12'b111111010100;
   37974: result <= 12'b111111010100;
   37975: result <= 12'b111111010100;
   37976: result <= 12'b111111010100;
   37977: result <= 12'b111111010100;
   37978: result <= 12'b111111010100;
   37979: result <= 12'b111111010101;
   37980: result <= 12'b111111010101;
   37981: result <= 12'b111111010101;
   37982: result <= 12'b111111010101;
   37983: result <= 12'b111111010101;
   37984: result <= 12'b111111010110;
   37985: result <= 12'b111111010110;
   37986: result <= 12'b111111010110;
   37987: result <= 12'b111111010110;
   37988: result <= 12'b111111010110;
   37989: result <= 12'b111111010110;
   37990: result <= 12'b111111010111;
   37991: result <= 12'b111111010111;
   37992: result <= 12'b111111010111;
   37993: result <= 12'b111111010111;
   37994: result <= 12'b111111010111;
   37995: result <= 12'b111111010111;
   37996: result <= 12'b111111011000;
   37997: result <= 12'b111111011000;
   37998: result <= 12'b111111011000;
   37999: result <= 12'b111111011000;
   38000: result <= 12'b111111011000;
   38001: result <= 12'b111111011000;
   38002: result <= 12'b111111011001;
   38003: result <= 12'b111111011001;
   38004: result <= 12'b111111011001;
   38005: result <= 12'b111111011001;
   38006: result <= 12'b111111011001;
   38007: result <= 12'b111111011001;
   38008: result <= 12'b111111011010;
   38009: result <= 12'b111111011010;
   38010: result <= 12'b111111011010;
   38011: result <= 12'b111111011010;
   38012: result <= 12'b111111011010;
   38013: result <= 12'b111111011010;
   38014: result <= 12'b111111011011;
   38015: result <= 12'b111111011011;
   38016: result <= 12'b111111011011;
   38017: result <= 12'b111111011011;
   38018: result <= 12'b111111011011;
   38019: result <= 12'b111111011100;
   38020: result <= 12'b111111011100;
   38021: result <= 12'b111111011100;
   38022: result <= 12'b111111011100;
   38023: result <= 12'b111111011100;
   38024: result <= 12'b111111011100;
   38025: result <= 12'b111111011101;
   38026: result <= 12'b111111011101;
   38027: result <= 12'b111111011101;
   38028: result <= 12'b111111011101;
   38029: result <= 12'b111111011101;
   38030: result <= 12'b111111011101;
   38031: result <= 12'b111111011110;
   38032: result <= 12'b111111011110;
   38033: result <= 12'b111111011110;
   38034: result <= 12'b111111011110;
   38035: result <= 12'b111111011110;
   38036: result <= 12'b111111011110;
   38037: result <= 12'b111111011111;
   38038: result <= 12'b111111011111;
   38039: result <= 12'b111111011111;
   38040: result <= 12'b111111011111;
   38041: result <= 12'b111111011111;
   38042: result <= 12'b111111011111;
   38043: result <= 12'b111111100000;
   38044: result <= 12'b111111100000;
   38045: result <= 12'b111111100000;
   38046: result <= 12'b111111100000;
   38047: result <= 12'b111111100000;
   38048: result <= 12'b111111100001;
   38049: result <= 12'b111111100001;
   38050: result <= 12'b111111100001;
   38051: result <= 12'b111111100001;
   38052: result <= 12'b111111100001;
   38053: result <= 12'b111111100001;
   38054: result <= 12'b111111100010;
   38055: result <= 12'b111111100010;
   38056: result <= 12'b111111100010;
   38057: result <= 12'b111111100010;
   38058: result <= 12'b111111100010;
   38059: result <= 12'b111111100010;
   38060: result <= 12'b111111100011;
   38061: result <= 12'b111111100011;
   38062: result <= 12'b111111100011;
   38063: result <= 12'b111111100011;
   38064: result <= 12'b111111100011;
   38065: result <= 12'b111111100011;
   38066: result <= 12'b111111100100;
   38067: result <= 12'b111111100100;
   38068: result <= 12'b111111100100;
   38069: result <= 12'b111111100100;
   38070: result <= 12'b111111100100;
   38071: result <= 12'b111111100100;
   38072: result <= 12'b111111100101;
   38073: result <= 12'b111111100101;
   38074: result <= 12'b111111100101;
   38075: result <= 12'b111111100101;
   38076: result <= 12'b111111100101;
   38077: result <= 12'b111111100101;
   38078: result <= 12'b111111100110;
   38079: result <= 12'b111111100110;
   38080: result <= 12'b111111100110;
   38081: result <= 12'b111111100110;
   38082: result <= 12'b111111100110;
   38083: result <= 12'b111111100111;
   38084: result <= 12'b111111100111;
   38085: result <= 12'b111111100111;
   38086: result <= 12'b111111100111;
   38087: result <= 12'b111111100111;
   38088: result <= 12'b111111100111;
   38089: result <= 12'b111111101000;
   38090: result <= 12'b111111101000;
   38091: result <= 12'b111111101000;
   38092: result <= 12'b111111101000;
   38093: result <= 12'b111111101000;
   38094: result <= 12'b111111101000;
   38095: result <= 12'b111111101001;
   38096: result <= 12'b111111101001;
   38097: result <= 12'b111111101001;
   38098: result <= 12'b111111101001;
   38099: result <= 12'b111111101001;
   38100: result <= 12'b111111101001;
   38101: result <= 12'b111111101010;
   38102: result <= 12'b111111101010;
   38103: result <= 12'b111111101010;
   38104: result <= 12'b111111101010;
   38105: result <= 12'b111111101010;
   38106: result <= 12'b111111101010;
   38107: result <= 12'b111111101011;
   38108: result <= 12'b111111101011;
   38109: result <= 12'b111111101011;
   38110: result <= 12'b111111101011;
   38111: result <= 12'b111111101011;
   38112: result <= 12'b111111101011;
   38113: result <= 12'b111111101100;
   38114: result <= 12'b111111101100;
   38115: result <= 12'b111111101100;
   38116: result <= 12'b111111101100;
   38117: result <= 12'b111111101100;
   38118: result <= 12'b111111101101;
   38119: result <= 12'b111111101101;
   38120: result <= 12'b111111101101;
   38121: result <= 12'b111111101101;
   38122: result <= 12'b111111101101;
   38123: result <= 12'b111111101101;
   38124: result <= 12'b111111101110;
   38125: result <= 12'b111111101110;
   38126: result <= 12'b111111101110;
   38127: result <= 12'b111111101110;
   38128: result <= 12'b111111101110;
   38129: result <= 12'b111111101110;
   38130: result <= 12'b111111101111;
   38131: result <= 12'b111111101111;
   38132: result <= 12'b111111101111;
   38133: result <= 12'b111111101111;
   38134: result <= 12'b111111101111;
   38135: result <= 12'b111111101111;
   38136: result <= 12'b111111110000;
   38137: result <= 12'b111111110000;
   38138: result <= 12'b111111110000;
   38139: result <= 12'b111111110000;
   38140: result <= 12'b111111110000;
   38141: result <= 12'b111111110000;
   38142: result <= 12'b111111110001;
   38143: result <= 12'b111111110001;
   38144: result <= 12'b111111110001;
   38145: result <= 12'b111111110001;
   38146: result <= 12'b111111110001;
   38147: result <= 12'b111111110001;
   38148: result <= 12'b111111110010;
   38149: result <= 12'b111111110010;
   38150: result <= 12'b111111110010;
   38151: result <= 12'b111111110010;
   38152: result <= 12'b111111110010;
   38153: result <= 12'b111111110010;
   38154: result <= 12'b111111110011;
   38155: result <= 12'b111111110011;
   38156: result <= 12'b111111110011;
   38157: result <= 12'b111111110011;
   38158: result <= 12'b111111110011;
   38159: result <= 12'b111111110100;
   38160: result <= 12'b111111110100;
   38161: result <= 12'b111111110100;
   38162: result <= 12'b111111110100;
   38163: result <= 12'b111111110100;
   38164: result <= 12'b111111110100;
   38165: result <= 12'b111111110101;
   38166: result <= 12'b111111110101;
   38167: result <= 12'b111111110101;
   38168: result <= 12'b111111110101;
   38169: result <= 12'b111111110101;
   38170: result <= 12'b111111110101;
   38171: result <= 12'b111111110110;
   38172: result <= 12'b111111110110;
   38173: result <= 12'b111111110110;
   38174: result <= 12'b111111110110;
   38175: result <= 12'b111111110110;
   38176: result <= 12'b111111110110;
   38177: result <= 12'b111111110111;
   38178: result <= 12'b111111110111;
   38179: result <= 12'b111111110111;
   38180: result <= 12'b111111110111;
   38181: result <= 12'b111111110111;
   38182: result <= 12'b111111110111;
   38183: result <= 12'b111111111000;
   38184: result <= 12'b111111111000;
   38185: result <= 12'b111111111000;
   38186: result <= 12'b111111111000;
   38187: result <= 12'b111111111000;
   38188: result <= 12'b111111111000;
   38189: result <= 12'b111111111001;
   38190: result <= 12'b111111111001;
   38191: result <= 12'b111111111001;
   38192: result <= 12'b111111111001;
   38193: result <= 12'b111111111001;
   38194: result <= 12'b111111111001;
   38195: result <= 12'b111111111010;
   38196: result <= 12'b111111111010;
   38197: result <= 12'b111111111010;
   38198: result <= 12'b111111111010;
   38199: result <= 12'b111111111010;
   38200: result <= 12'b111111111011;
   38201: result <= 12'b111111111011;
   38202: result <= 12'b111111111011;
   38203: result <= 12'b111111111011;
   38204: result <= 12'b111111111011;
   38205: result <= 12'b111111111011;
   38206: result <= 12'b111111111100;
   38207: result <= 12'b111111111100;
   38208: result <= 12'b111111111100;
   38209: result <= 12'b111111111100;
   38210: result <= 12'b111111111100;
   38211: result <= 12'b111111111100;
   38212: result <= 12'b111111111101;
   38213: result <= 12'b111111111101;
   38214: result <= 12'b111111111101;
   38215: result <= 12'b111111111101;
   38216: result <= 12'b111111111101;
   38217: result <= 12'b111111111101;
   38218: result <= 12'b111111111110;
   38219: result <= 12'b111111111110;
   38220: result <= 12'b111111111110;
   38221: result <= 12'b111111111110;
   38222: result <= 12'b111111111110;
   38223: result <= 12'b111111111110;
   38224: result <= 12'b111111111111;
   38225: result <= 12'b111111111111;
   38226: result <= 12'b111111111111;
   38227: result <= 12'b111111111111;
   38228: result <= 12'b111111111111;
   38229: result <= 12'b111111111111;
   38230: result <= 12'b110000000000;
   38231: result <= 12'b110000000000;
   38232: result <= 12'b110000000000;
   38233: result <= 12'b110000000000;
   38234: result <= 12'b110000000000;
   38235: result <= 12'b110000000000;
   38236: result <= 12'b110000000001;
   38237: result <= 12'b110000000001;
   38238: result <= 12'b110000000001;
   38239: result <= 12'b110000000001;
   38240: result <= 12'b110000000001;
   38241: result <= 12'b110000000001;
   38242: result <= 12'b110000000010;
   38243: result <= 12'b110000000010;
   38244: result <= 12'b110000000010;
   38245: result <= 12'b110000000010;
   38246: result <= 12'b110000000010;
   38247: result <= 12'b110000000011;
   38248: result <= 12'b110000000011;
   38249: result <= 12'b110000000011;
   38250: result <= 12'b110000000011;
   38251: result <= 12'b110000000011;
   38252: result <= 12'b110000000011;
   38253: result <= 12'b110000000100;
   38254: result <= 12'b110000000100;
   38255: result <= 12'b110000000100;
   38256: result <= 12'b110000000100;
   38257: result <= 12'b110000000100;
   38258: result <= 12'b110000000100;
   38259: result <= 12'b110000000101;
   38260: result <= 12'b110000000101;
   38261: result <= 12'b110000000101;
   38262: result <= 12'b110000000101;
   38263: result <= 12'b110000000101;
   38264: result <= 12'b110000000101;
   38265: result <= 12'b110000000110;
   38266: result <= 12'b110000000110;
   38267: result <= 12'b110000000110;
   38268: result <= 12'b110000000110;
   38269: result <= 12'b110000000110;
   38270: result <= 12'b110000000110;
   38271: result <= 12'b110000000111;
   38272: result <= 12'b110000000111;
   38273: result <= 12'b110000000111;
   38274: result <= 12'b110000000111;
   38275: result <= 12'b110000000111;
   38276: result <= 12'b110000000111;
   38277: result <= 12'b110000001000;
   38278: result <= 12'b110000001000;
   38279: result <= 12'b110000001000;
   38280: result <= 12'b110000001000;
   38281: result <= 12'b110000001000;
   38282: result <= 12'b110000001000;
   38283: result <= 12'b110000001001;
   38284: result <= 12'b110000001001;
   38285: result <= 12'b110000001001;
   38286: result <= 12'b110000001001;
   38287: result <= 12'b110000001001;
   38288: result <= 12'b110000001001;
   38289: result <= 12'b110000001010;
   38290: result <= 12'b110000001010;
   38291: result <= 12'b110000001010;
   38292: result <= 12'b110000001010;
   38293: result <= 12'b110000001010;
   38294: result <= 12'b110000001010;
   38295: result <= 12'b110000001011;
   38296: result <= 12'b110000001011;
   38297: result <= 12'b110000001011;
   38298: result <= 12'b110000001011;
   38299: result <= 12'b110000001011;
   38300: result <= 12'b110000001011;
   38301: result <= 12'b110000001100;
   38302: result <= 12'b110000001100;
   38303: result <= 12'b110000001100;
   38304: result <= 12'b110000001100;
   38305: result <= 12'b110000001100;
   38306: result <= 12'b110000001101;
   38307: result <= 12'b110000001101;
   38308: result <= 12'b110000001101;
   38309: result <= 12'b110000001101;
   38310: result <= 12'b110000001101;
   38311: result <= 12'b110000001101;
   38312: result <= 12'b110000001110;
   38313: result <= 12'b110000001110;
   38314: result <= 12'b110000001110;
   38315: result <= 12'b110000001110;
   38316: result <= 12'b110000001110;
   38317: result <= 12'b110000001110;
   38318: result <= 12'b110000001111;
   38319: result <= 12'b110000001111;
   38320: result <= 12'b110000001111;
   38321: result <= 12'b110000001111;
   38322: result <= 12'b110000001111;
   38323: result <= 12'b110000001111;
   38324: result <= 12'b110000010000;
   38325: result <= 12'b110000010000;
   38326: result <= 12'b110000010000;
   38327: result <= 12'b110000010000;
   38328: result <= 12'b110000010000;
   38329: result <= 12'b110000010000;
   38330: result <= 12'b110000010001;
   38331: result <= 12'b110000010001;
   38332: result <= 12'b110000010001;
   38333: result <= 12'b110000010001;
   38334: result <= 12'b110000010001;
   38335: result <= 12'b110000010001;
   38336: result <= 12'b110000010010;
   38337: result <= 12'b110000010010;
   38338: result <= 12'b110000010010;
   38339: result <= 12'b110000010010;
   38340: result <= 12'b110000010010;
   38341: result <= 12'b110000010010;
   38342: result <= 12'b110000010011;
   38343: result <= 12'b110000010011;
   38344: result <= 12'b110000010011;
   38345: result <= 12'b110000010011;
   38346: result <= 12'b110000010011;
   38347: result <= 12'b110000010011;
   38348: result <= 12'b110000010100;
   38349: result <= 12'b110000010100;
   38350: result <= 12'b110000010100;
   38351: result <= 12'b110000010100;
   38352: result <= 12'b110000010100;
   38353: result <= 12'b110000010100;
   38354: result <= 12'b110000010101;
   38355: result <= 12'b110000010101;
   38356: result <= 12'b110000010101;
   38357: result <= 12'b110000010101;
   38358: result <= 12'b110000010101;
   38359: result <= 12'b110000010101;
   38360: result <= 12'b110000010110;
   38361: result <= 12'b110000010110;
   38362: result <= 12'b110000010110;
   38363: result <= 12'b110000010110;
   38364: result <= 12'b110000010110;
   38365: result <= 12'b110000010110;
   38366: result <= 12'b110000010111;
   38367: result <= 12'b110000010111;
   38368: result <= 12'b110000010111;
   38369: result <= 12'b110000010111;
   38370: result <= 12'b110000010111;
   38371: result <= 12'b110000010111;
   38372: result <= 12'b110000011000;
   38373: result <= 12'b110000011000;
   38374: result <= 12'b110000011000;
   38375: result <= 12'b110000011000;
   38376: result <= 12'b110000011000;
   38377: result <= 12'b110000011001;
   38378: result <= 12'b110000011001;
   38379: result <= 12'b110000011001;
   38380: result <= 12'b110000011001;
   38381: result <= 12'b110000011001;
   38382: result <= 12'b110000011001;
   38383: result <= 12'b110000011010;
   38384: result <= 12'b110000011010;
   38385: result <= 12'b110000011010;
   38386: result <= 12'b110000011010;
   38387: result <= 12'b110000011010;
   38388: result <= 12'b110000011010;
   38389: result <= 12'b110000011011;
   38390: result <= 12'b110000011011;
   38391: result <= 12'b110000011011;
   38392: result <= 12'b110000011011;
   38393: result <= 12'b110000011011;
   38394: result <= 12'b110000011011;
   38395: result <= 12'b110000011100;
   38396: result <= 12'b110000011100;
   38397: result <= 12'b110000011100;
   38398: result <= 12'b110000011100;
   38399: result <= 12'b110000011100;
   38400: result <= 12'b110000011100;
   38401: result <= 12'b110000011101;
   38402: result <= 12'b110000011101;
   38403: result <= 12'b110000011101;
   38404: result <= 12'b110000011101;
   38405: result <= 12'b110000011101;
   38406: result <= 12'b110000011101;
   38407: result <= 12'b110000011110;
   38408: result <= 12'b110000011110;
   38409: result <= 12'b110000011110;
   38410: result <= 12'b110000011110;
   38411: result <= 12'b110000011110;
   38412: result <= 12'b110000011110;
   38413: result <= 12'b110000011111;
   38414: result <= 12'b110000011111;
   38415: result <= 12'b110000011111;
   38416: result <= 12'b110000011111;
   38417: result <= 12'b110000011111;
   38418: result <= 12'b110000011111;
   38419: result <= 12'b110000100000;
   38420: result <= 12'b110000100000;
   38421: result <= 12'b110000100000;
   38422: result <= 12'b110000100000;
   38423: result <= 12'b110000100000;
   38424: result <= 12'b110000100000;
   38425: result <= 12'b110000100001;
   38426: result <= 12'b110000100001;
   38427: result <= 12'b110000100001;
   38428: result <= 12'b110000100001;
   38429: result <= 12'b110000100001;
   38430: result <= 12'b110000100001;
   38431: result <= 12'b110000100010;
   38432: result <= 12'b110000100010;
   38433: result <= 12'b110000100010;
   38434: result <= 12'b110000100010;
   38435: result <= 12'b110000100010;
   38436: result <= 12'b110000100010;
   38437: result <= 12'b110000100011;
   38438: result <= 12'b110000100011;
   38439: result <= 12'b110000100011;
   38440: result <= 12'b110000100011;
   38441: result <= 12'b110000100011;
   38442: result <= 12'b110000100011;
   38443: result <= 12'b110000100100;
   38444: result <= 12'b110000100100;
   38445: result <= 12'b110000100100;
   38446: result <= 12'b110000100100;
   38447: result <= 12'b110000100100;
   38448: result <= 12'b110000100100;
   38449: result <= 12'b110000100101;
   38450: result <= 12'b110000100101;
   38451: result <= 12'b110000100101;
   38452: result <= 12'b110000100101;
   38453: result <= 12'b110000100101;
   38454: result <= 12'b110000100101;
   38455: result <= 12'b110000100110;
   38456: result <= 12'b110000100110;
   38457: result <= 12'b110000100110;
   38458: result <= 12'b110000100110;
   38459: result <= 12'b110000100110;
   38460: result <= 12'b110000100110;
   38461: result <= 12'b110000100111;
   38462: result <= 12'b110000100111;
   38463: result <= 12'b110000100111;
   38464: result <= 12'b110000100111;
   38465: result <= 12'b110000100111;
   38466: result <= 12'b110000100111;
   38467: result <= 12'b110000101000;
   38468: result <= 12'b110000101000;
   38469: result <= 12'b110000101000;
   38470: result <= 12'b110000101000;
   38471: result <= 12'b110000101000;
   38472: result <= 12'b110000101000;
   38473: result <= 12'b110000101001;
   38474: result <= 12'b110000101001;
   38475: result <= 12'b110000101001;
   38476: result <= 12'b110000101001;
   38477: result <= 12'b110000101001;
   38478: result <= 12'b110000101001;
   38479: result <= 12'b110000101010;
   38480: result <= 12'b110000101010;
   38481: result <= 12'b110000101010;
   38482: result <= 12'b110000101010;
   38483: result <= 12'b110000101010;
   38484: result <= 12'b110000101010;
   38485: result <= 12'b110000101011;
   38486: result <= 12'b110000101011;
   38487: result <= 12'b110000101011;
   38488: result <= 12'b110000101011;
   38489: result <= 12'b110000101011;
   38490: result <= 12'b110000101100;
   38491: result <= 12'b110000101100;
   38492: result <= 12'b110000101100;
   38493: result <= 12'b110000101100;
   38494: result <= 12'b110000101100;
   38495: result <= 12'b110000101100;
   38496: result <= 12'b110000101101;
   38497: result <= 12'b110000101101;
   38498: result <= 12'b110000101101;
   38499: result <= 12'b110000101101;
   38500: result <= 12'b110000101101;
   38501: result <= 12'b110000101101;
   38502: result <= 12'b110000101110;
   38503: result <= 12'b110000101110;
   38504: result <= 12'b110000101110;
   38505: result <= 12'b110000101110;
   38506: result <= 12'b110000101110;
   38507: result <= 12'b110000101110;
   38508: result <= 12'b110000101111;
   38509: result <= 12'b110000101111;
   38510: result <= 12'b110000101111;
   38511: result <= 12'b110000101111;
   38512: result <= 12'b110000101111;
   38513: result <= 12'b110000101111;
   38514: result <= 12'b110000110000;
   38515: result <= 12'b110000110000;
   38516: result <= 12'b110000110000;
   38517: result <= 12'b110000110000;
   38518: result <= 12'b110000110000;
   38519: result <= 12'b110000110000;
   38520: result <= 12'b110000110001;
   38521: result <= 12'b110000110001;
   38522: result <= 12'b110000110001;
   38523: result <= 12'b110000110001;
   38524: result <= 12'b110000110001;
   38525: result <= 12'b110000110001;
   38526: result <= 12'b110000110010;
   38527: result <= 12'b110000110010;
   38528: result <= 12'b110000110010;
   38529: result <= 12'b110000110010;
   38530: result <= 12'b110000110010;
   38531: result <= 12'b110000110010;
   38532: result <= 12'b110000110011;
   38533: result <= 12'b110000110011;
   38534: result <= 12'b110000110011;
   38535: result <= 12'b110000110011;
   38536: result <= 12'b110000110011;
   38537: result <= 12'b110000110011;
   38538: result <= 12'b110000110100;
   38539: result <= 12'b110000110100;
   38540: result <= 12'b110000110100;
   38541: result <= 12'b110000110100;
   38542: result <= 12'b110000110100;
   38543: result <= 12'b110000110100;
   38544: result <= 12'b110000110101;
   38545: result <= 12'b110000110101;
   38546: result <= 12'b110000110101;
   38547: result <= 12'b110000110101;
   38548: result <= 12'b110000110101;
   38549: result <= 12'b110000110101;
   38550: result <= 12'b110000110110;
   38551: result <= 12'b110000110110;
   38552: result <= 12'b110000110110;
   38553: result <= 12'b110000110110;
   38554: result <= 12'b110000110110;
   38555: result <= 12'b110000110110;
   38556: result <= 12'b110000110111;
   38557: result <= 12'b110000110111;
   38558: result <= 12'b110000110111;
   38559: result <= 12'b110000110111;
   38560: result <= 12'b110000110111;
   38561: result <= 12'b110000110111;
   38562: result <= 12'b110000111000;
   38563: result <= 12'b110000111000;
   38564: result <= 12'b110000111000;
   38565: result <= 12'b110000111000;
   38566: result <= 12'b110000111000;
   38567: result <= 12'b110000111000;
   38568: result <= 12'b110000111001;
   38569: result <= 12'b110000111001;
   38570: result <= 12'b110000111001;
   38571: result <= 12'b110000111001;
   38572: result <= 12'b110000111001;
   38573: result <= 12'b110000111001;
   38574: result <= 12'b110000111010;
   38575: result <= 12'b110000111010;
   38576: result <= 12'b110000111010;
   38577: result <= 12'b110000111010;
   38578: result <= 12'b110000111010;
   38579: result <= 12'b110000111010;
   38580: result <= 12'b110000111011;
   38581: result <= 12'b110000111011;
   38582: result <= 12'b110000111011;
   38583: result <= 12'b110000111011;
   38584: result <= 12'b110000111011;
   38585: result <= 12'b110000111011;
   38586: result <= 12'b110000111100;
   38587: result <= 12'b110000111100;
   38588: result <= 12'b110000111100;
   38589: result <= 12'b110000111100;
   38590: result <= 12'b110000111100;
   38591: result <= 12'b110000111100;
   38592: result <= 12'b110000111101;
   38593: result <= 12'b110000111101;
   38594: result <= 12'b110000111101;
   38595: result <= 12'b110000111101;
   38596: result <= 12'b110000111101;
   38597: result <= 12'b110000111101;
   38598: result <= 12'b110000111110;
   38599: result <= 12'b110000111110;
   38600: result <= 12'b110000111110;
   38601: result <= 12'b110000111110;
   38602: result <= 12'b110000111110;
   38603: result <= 12'b110000111110;
   38604: result <= 12'b110000111111;
   38605: result <= 12'b110000111111;
   38606: result <= 12'b110000111111;
   38607: result <= 12'b110000111111;
   38608: result <= 12'b110000111111;
   38609: result <= 12'b110000111111;
   38610: result <= 12'b110001000000;
   38611: result <= 12'b110001000000;
   38612: result <= 12'b110001000000;
   38613: result <= 12'b110001000000;
   38614: result <= 12'b110001000000;
   38615: result <= 12'b110001000000;
   38616: result <= 12'b110001000001;
   38617: result <= 12'b110001000001;
   38618: result <= 12'b110001000001;
   38619: result <= 12'b110001000001;
   38620: result <= 12'b110001000001;
   38621: result <= 12'b110001000001;
   38622: result <= 12'b110001000010;
   38623: result <= 12'b110001000010;
   38624: result <= 12'b110001000010;
   38625: result <= 12'b110001000010;
   38626: result <= 12'b110001000010;
   38627: result <= 12'b110001000010;
   38628: result <= 12'b110001000011;
   38629: result <= 12'b110001000011;
   38630: result <= 12'b110001000011;
   38631: result <= 12'b110001000011;
   38632: result <= 12'b110001000011;
   38633: result <= 12'b110001000011;
   38634: result <= 12'b110001000100;
   38635: result <= 12'b110001000100;
   38636: result <= 12'b110001000100;
   38637: result <= 12'b110001000100;
   38638: result <= 12'b110001000100;
   38639: result <= 12'b110001000100;
   38640: result <= 12'b110001000101;
   38641: result <= 12'b110001000101;
   38642: result <= 12'b110001000101;
   38643: result <= 12'b110001000101;
   38644: result <= 12'b110001000101;
   38645: result <= 12'b110001000101;
   38646: result <= 12'b110001000110;
   38647: result <= 12'b110001000110;
   38648: result <= 12'b110001000110;
   38649: result <= 12'b110001000110;
   38650: result <= 12'b110001000110;
   38651: result <= 12'b110001000110;
   38652: result <= 12'b110001000111;
   38653: result <= 12'b110001000111;
   38654: result <= 12'b110001000111;
   38655: result <= 12'b110001000111;
   38656: result <= 12'b110001000111;
   38657: result <= 12'b110001000111;
   38658: result <= 12'b110001001000;
   38659: result <= 12'b110001001000;
   38660: result <= 12'b110001001000;
   38661: result <= 12'b110001001000;
   38662: result <= 12'b110001001000;
   38663: result <= 12'b110001001000;
   38664: result <= 12'b110001001001;
   38665: result <= 12'b110001001001;
   38666: result <= 12'b110001001001;
   38667: result <= 12'b110001001001;
   38668: result <= 12'b110001001001;
   38669: result <= 12'b110001001001;
   38670: result <= 12'b110001001001;
   38671: result <= 12'b110001001010;
   38672: result <= 12'b110001001010;
   38673: result <= 12'b110001001010;
   38674: result <= 12'b110001001010;
   38675: result <= 12'b110001001010;
   38676: result <= 12'b110001001010;
   38677: result <= 12'b110001001011;
   38678: result <= 12'b110001001011;
   38679: result <= 12'b110001001011;
   38680: result <= 12'b110001001011;
   38681: result <= 12'b110001001011;
   38682: result <= 12'b110001001011;
   38683: result <= 12'b110001001100;
   38684: result <= 12'b110001001100;
   38685: result <= 12'b110001001100;
   38686: result <= 12'b110001001100;
   38687: result <= 12'b110001001100;
   38688: result <= 12'b110001001100;
   38689: result <= 12'b110001001101;
   38690: result <= 12'b110001001101;
   38691: result <= 12'b110001001101;
   38692: result <= 12'b110001001101;
   38693: result <= 12'b110001001101;
   38694: result <= 12'b110001001101;
   38695: result <= 12'b110001001110;
   38696: result <= 12'b110001001110;
   38697: result <= 12'b110001001110;
   38698: result <= 12'b110001001110;
   38699: result <= 12'b110001001110;
   38700: result <= 12'b110001001110;
   38701: result <= 12'b110001001111;
   38702: result <= 12'b110001001111;
   38703: result <= 12'b110001001111;
   38704: result <= 12'b110001001111;
   38705: result <= 12'b110001001111;
   38706: result <= 12'b110001001111;
   38707: result <= 12'b110001010000;
   38708: result <= 12'b110001010000;
   38709: result <= 12'b110001010000;
   38710: result <= 12'b110001010000;
   38711: result <= 12'b110001010000;
   38712: result <= 12'b110001010000;
   38713: result <= 12'b110001010001;
   38714: result <= 12'b110001010001;
   38715: result <= 12'b110001010001;
   38716: result <= 12'b110001010001;
   38717: result <= 12'b110001010001;
   38718: result <= 12'b110001010001;
   38719: result <= 12'b110001010010;
   38720: result <= 12'b110001010010;
   38721: result <= 12'b110001010010;
   38722: result <= 12'b110001010010;
   38723: result <= 12'b110001010010;
   38724: result <= 12'b110001010010;
   38725: result <= 12'b110001010011;
   38726: result <= 12'b110001010011;
   38727: result <= 12'b110001010011;
   38728: result <= 12'b110001010011;
   38729: result <= 12'b110001010011;
   38730: result <= 12'b110001010011;
   38731: result <= 12'b110001010100;
   38732: result <= 12'b110001010100;
   38733: result <= 12'b110001010100;
   38734: result <= 12'b110001010100;
   38735: result <= 12'b110001010100;
   38736: result <= 12'b110001010100;
   38737: result <= 12'b110001010101;
   38738: result <= 12'b110001010101;
   38739: result <= 12'b110001010101;
   38740: result <= 12'b110001010101;
   38741: result <= 12'b110001010101;
   38742: result <= 12'b110001010101;
   38743: result <= 12'b110001010110;
   38744: result <= 12'b110001010110;
   38745: result <= 12'b110001010110;
   38746: result <= 12'b110001010110;
   38747: result <= 12'b110001010110;
   38748: result <= 12'b110001010110;
   38749: result <= 12'b110001010111;
   38750: result <= 12'b110001010111;
   38751: result <= 12'b110001010111;
   38752: result <= 12'b110001010111;
   38753: result <= 12'b110001010111;
   38754: result <= 12'b110001010111;
   38755: result <= 12'b110001011000;
   38756: result <= 12'b110001011000;
   38757: result <= 12'b110001011000;
   38758: result <= 12'b110001011000;
   38759: result <= 12'b110001011000;
   38760: result <= 12'b110001011000;
   38761: result <= 12'b110001011001;
   38762: result <= 12'b110001011001;
   38763: result <= 12'b110001011001;
   38764: result <= 12'b110001011001;
   38765: result <= 12'b110001011001;
   38766: result <= 12'b110001011001;
   38767: result <= 12'b110001011010;
   38768: result <= 12'b110001011010;
   38769: result <= 12'b110001011010;
   38770: result <= 12'b110001011010;
   38771: result <= 12'b110001011010;
   38772: result <= 12'b110001011010;
   38773: result <= 12'b110001011011;
   38774: result <= 12'b110001011011;
   38775: result <= 12'b110001011011;
   38776: result <= 12'b110001011011;
   38777: result <= 12'b110001011011;
   38778: result <= 12'b110001011011;
   38779: result <= 12'b110001011100;
   38780: result <= 12'b110001011100;
   38781: result <= 12'b110001011100;
   38782: result <= 12'b110001011100;
   38783: result <= 12'b110001011100;
   38784: result <= 12'b110001011100;
   38785: result <= 12'b110001011100;
   38786: result <= 12'b110001011101;
   38787: result <= 12'b110001011101;
   38788: result <= 12'b110001011101;
   38789: result <= 12'b110001011101;
   38790: result <= 12'b110001011101;
   38791: result <= 12'b110001011101;
   38792: result <= 12'b110001011110;
   38793: result <= 12'b110001011110;
   38794: result <= 12'b110001011110;
   38795: result <= 12'b110001011110;
   38796: result <= 12'b110001011110;
   38797: result <= 12'b110001011110;
   38798: result <= 12'b110001011111;
   38799: result <= 12'b110001011111;
   38800: result <= 12'b110001011111;
   38801: result <= 12'b110001011111;
   38802: result <= 12'b110001011111;
   38803: result <= 12'b110001011111;
   38804: result <= 12'b110001100000;
   38805: result <= 12'b110001100000;
   38806: result <= 12'b110001100000;
   38807: result <= 12'b110001100000;
   38808: result <= 12'b110001100000;
   38809: result <= 12'b110001100000;
   38810: result <= 12'b110001100001;
   38811: result <= 12'b110001100001;
   38812: result <= 12'b110001100001;
   38813: result <= 12'b110001100001;
   38814: result <= 12'b110001100001;
   38815: result <= 12'b110001100001;
   38816: result <= 12'b110001100010;
   38817: result <= 12'b110001100010;
   38818: result <= 12'b110001100010;
   38819: result <= 12'b110001100010;
   38820: result <= 12'b110001100010;
   38821: result <= 12'b110001100010;
   38822: result <= 12'b110001100011;
   38823: result <= 12'b110001100011;
   38824: result <= 12'b110001100011;
   38825: result <= 12'b110001100011;
   38826: result <= 12'b110001100011;
   38827: result <= 12'b110001100011;
   38828: result <= 12'b110001100100;
   38829: result <= 12'b110001100100;
   38830: result <= 12'b110001100100;
   38831: result <= 12'b110001100100;
   38832: result <= 12'b110001100100;
   38833: result <= 12'b110001100100;
   38834: result <= 12'b110001100101;
   38835: result <= 12'b110001100101;
   38836: result <= 12'b110001100101;
   38837: result <= 12'b110001100101;
   38838: result <= 12'b110001100101;
   38839: result <= 12'b110001100101;
   38840: result <= 12'b110001100110;
   38841: result <= 12'b110001100110;
   38842: result <= 12'b110001100110;
   38843: result <= 12'b110001100110;
   38844: result <= 12'b110001100110;
   38845: result <= 12'b110001100110;
   38846: result <= 12'b110001100111;
   38847: result <= 12'b110001100111;
   38848: result <= 12'b110001100111;
   38849: result <= 12'b110001100111;
   38850: result <= 12'b110001100111;
   38851: result <= 12'b110001100111;
   38852: result <= 12'b110001100111;
   38853: result <= 12'b110001101000;
   38854: result <= 12'b110001101000;
   38855: result <= 12'b110001101000;
   38856: result <= 12'b110001101000;
   38857: result <= 12'b110001101000;
   38858: result <= 12'b110001101000;
   38859: result <= 12'b110001101001;
   38860: result <= 12'b110001101001;
   38861: result <= 12'b110001101001;
   38862: result <= 12'b110001101001;
   38863: result <= 12'b110001101001;
   38864: result <= 12'b110001101001;
   38865: result <= 12'b110001101010;
   38866: result <= 12'b110001101010;
   38867: result <= 12'b110001101010;
   38868: result <= 12'b110001101010;
   38869: result <= 12'b110001101010;
   38870: result <= 12'b110001101010;
   38871: result <= 12'b110001101011;
   38872: result <= 12'b110001101011;
   38873: result <= 12'b110001101011;
   38874: result <= 12'b110001101011;
   38875: result <= 12'b110001101011;
   38876: result <= 12'b110001101011;
   38877: result <= 12'b110001101100;
   38878: result <= 12'b110001101100;
   38879: result <= 12'b110001101100;
   38880: result <= 12'b110001101100;
   38881: result <= 12'b110001101100;
   38882: result <= 12'b110001101100;
   38883: result <= 12'b110001101101;
   38884: result <= 12'b110001101101;
   38885: result <= 12'b110001101101;
   38886: result <= 12'b110001101101;
   38887: result <= 12'b110001101101;
   38888: result <= 12'b110001101101;
   38889: result <= 12'b110001101110;
   38890: result <= 12'b110001101110;
   38891: result <= 12'b110001101110;
   38892: result <= 12'b110001101110;
   38893: result <= 12'b110001101110;
   38894: result <= 12'b110001101110;
   38895: result <= 12'b110001101111;
   38896: result <= 12'b110001101111;
   38897: result <= 12'b110001101111;
   38898: result <= 12'b110001101111;
   38899: result <= 12'b110001101111;
   38900: result <= 12'b110001101111;
   38901: result <= 12'b110001110000;
   38902: result <= 12'b110001110000;
   38903: result <= 12'b110001110000;
   38904: result <= 12'b110001110000;
   38905: result <= 12'b110001110000;
   38906: result <= 12'b110001110000;
   38907: result <= 12'b110001110000;
   38908: result <= 12'b110001110001;
   38909: result <= 12'b110001110001;
   38910: result <= 12'b110001110001;
   38911: result <= 12'b110001110001;
   38912: result <= 12'b110001110001;
   38913: result <= 12'b110001110001;
   38914: result <= 12'b110001110010;
   38915: result <= 12'b110001110010;
   38916: result <= 12'b110001110010;
   38917: result <= 12'b110001110010;
   38918: result <= 12'b110001110010;
   38919: result <= 12'b110001110010;
   38920: result <= 12'b110001110011;
   38921: result <= 12'b110001110011;
   38922: result <= 12'b110001110011;
   38923: result <= 12'b110001110011;
   38924: result <= 12'b110001110011;
   38925: result <= 12'b110001110011;
   38926: result <= 12'b110001110100;
   38927: result <= 12'b110001110100;
   38928: result <= 12'b110001110100;
   38929: result <= 12'b110001110100;
   38930: result <= 12'b110001110100;
   38931: result <= 12'b110001110100;
   38932: result <= 12'b110001110101;
   38933: result <= 12'b110001110101;
   38934: result <= 12'b110001110101;
   38935: result <= 12'b110001110101;
   38936: result <= 12'b110001110101;
   38937: result <= 12'b110001110101;
   38938: result <= 12'b110001110110;
   38939: result <= 12'b110001110110;
   38940: result <= 12'b110001110110;
   38941: result <= 12'b110001110110;
   38942: result <= 12'b110001110110;
   38943: result <= 12'b110001110110;
   38944: result <= 12'b110001110111;
   38945: result <= 12'b110001110111;
   38946: result <= 12'b110001110111;
   38947: result <= 12'b110001110111;
   38948: result <= 12'b110001110111;
   38949: result <= 12'b110001110111;
   38950: result <= 12'b110001111000;
   38951: result <= 12'b110001111000;
   38952: result <= 12'b110001111000;
   38953: result <= 12'b110001111000;
   38954: result <= 12'b110001111000;
   38955: result <= 12'b110001111000;
   38956: result <= 12'b110001111000;
   38957: result <= 12'b110001111001;
   38958: result <= 12'b110001111001;
   38959: result <= 12'b110001111001;
   38960: result <= 12'b110001111001;
   38961: result <= 12'b110001111001;
   38962: result <= 12'b110001111001;
   38963: result <= 12'b110001111010;
   38964: result <= 12'b110001111010;
   38965: result <= 12'b110001111010;
   38966: result <= 12'b110001111010;
   38967: result <= 12'b110001111010;
   38968: result <= 12'b110001111010;
   38969: result <= 12'b110001111011;
   38970: result <= 12'b110001111011;
   38971: result <= 12'b110001111011;
   38972: result <= 12'b110001111011;
   38973: result <= 12'b110001111011;
   38974: result <= 12'b110001111011;
   38975: result <= 12'b110001111100;
   38976: result <= 12'b110001111100;
   38977: result <= 12'b110001111100;
   38978: result <= 12'b110001111100;
   38979: result <= 12'b110001111100;
   38980: result <= 12'b110001111100;
   38981: result <= 12'b110001111101;
   38982: result <= 12'b110001111101;
   38983: result <= 12'b110001111101;
   38984: result <= 12'b110001111101;
   38985: result <= 12'b110001111101;
   38986: result <= 12'b110001111101;
   38987: result <= 12'b110001111110;
   38988: result <= 12'b110001111110;
   38989: result <= 12'b110001111110;
   38990: result <= 12'b110001111110;
   38991: result <= 12'b110001111110;
   38992: result <= 12'b110001111110;
   38993: result <= 12'b110001111110;
   38994: result <= 12'b110001111111;
   38995: result <= 12'b110001111111;
   38996: result <= 12'b110001111111;
   38997: result <= 12'b110001111111;
   38998: result <= 12'b110001111111;
   38999: result <= 12'b110001111111;
   39000: result <= 12'b110010000000;
   39001: result <= 12'b110010000000;
   39002: result <= 12'b110010000000;
   39003: result <= 12'b110010000000;
   39004: result <= 12'b110010000000;
   39005: result <= 12'b110010000000;
   39006: result <= 12'b110010000001;
   39007: result <= 12'b110010000001;
   39008: result <= 12'b110010000001;
   39009: result <= 12'b110010000001;
   39010: result <= 12'b110010000001;
   39011: result <= 12'b110010000001;
   39012: result <= 12'b110010000010;
   39013: result <= 12'b110010000010;
   39014: result <= 12'b110010000010;
   39015: result <= 12'b110010000010;
   39016: result <= 12'b110010000010;
   39017: result <= 12'b110010000010;
   39018: result <= 12'b110010000011;
   39019: result <= 12'b110010000011;
   39020: result <= 12'b110010000011;
   39021: result <= 12'b110010000011;
   39022: result <= 12'b110010000011;
   39023: result <= 12'b110010000011;
   39024: result <= 12'b110010000100;
   39025: result <= 12'b110010000100;
   39026: result <= 12'b110010000100;
   39027: result <= 12'b110010000100;
   39028: result <= 12'b110010000100;
   39029: result <= 12'b110010000100;
   39030: result <= 12'b110010000100;
   39031: result <= 12'b110010000101;
   39032: result <= 12'b110010000101;
   39033: result <= 12'b110010000101;
   39034: result <= 12'b110010000101;
   39035: result <= 12'b110010000101;
   39036: result <= 12'b110010000101;
   39037: result <= 12'b110010000110;
   39038: result <= 12'b110010000110;
   39039: result <= 12'b110010000110;
   39040: result <= 12'b110010000110;
   39041: result <= 12'b110010000110;
   39042: result <= 12'b110010000110;
   39043: result <= 12'b110010000111;
   39044: result <= 12'b110010000111;
   39045: result <= 12'b110010000111;
   39046: result <= 12'b110010000111;
   39047: result <= 12'b110010000111;
   39048: result <= 12'b110010000111;
   39049: result <= 12'b110010001000;
   39050: result <= 12'b110010001000;
   39051: result <= 12'b110010001000;
   39052: result <= 12'b110010001000;
   39053: result <= 12'b110010001000;
   39054: result <= 12'b110010001000;
   39055: result <= 12'b110010001001;
   39056: result <= 12'b110010001001;
   39057: result <= 12'b110010001001;
   39058: result <= 12'b110010001001;
   39059: result <= 12'b110010001001;
   39060: result <= 12'b110010001001;
   39061: result <= 12'b110010001010;
   39062: result <= 12'b110010001010;
   39063: result <= 12'b110010001010;
   39064: result <= 12'b110010001010;
   39065: result <= 12'b110010001010;
   39066: result <= 12'b110010001010;
   39067: result <= 12'b110010001010;
   39068: result <= 12'b110010001011;
   39069: result <= 12'b110010001011;
   39070: result <= 12'b110010001011;
   39071: result <= 12'b110010001011;
   39072: result <= 12'b110010001011;
   39073: result <= 12'b110010001011;
   39074: result <= 12'b110010001100;
   39075: result <= 12'b110010001100;
   39076: result <= 12'b110010001100;
   39077: result <= 12'b110010001100;
   39078: result <= 12'b110010001100;
   39079: result <= 12'b110010001100;
   39080: result <= 12'b110010001101;
   39081: result <= 12'b110010001101;
   39082: result <= 12'b110010001101;
   39083: result <= 12'b110010001101;
   39084: result <= 12'b110010001101;
   39085: result <= 12'b110010001101;
   39086: result <= 12'b110010001110;
   39087: result <= 12'b110010001110;
   39088: result <= 12'b110010001110;
   39089: result <= 12'b110010001110;
   39090: result <= 12'b110010001110;
   39091: result <= 12'b110010001110;
   39092: result <= 12'b110010001111;
   39093: result <= 12'b110010001111;
   39094: result <= 12'b110010001111;
   39095: result <= 12'b110010001111;
   39096: result <= 12'b110010001111;
   39097: result <= 12'b110010001111;
   39098: result <= 12'b110010001111;
   39099: result <= 12'b110010010000;
   39100: result <= 12'b110010010000;
   39101: result <= 12'b110010010000;
   39102: result <= 12'b110010010000;
   39103: result <= 12'b110010010000;
   39104: result <= 12'b110010010000;
   39105: result <= 12'b110010010001;
   39106: result <= 12'b110010010001;
   39107: result <= 12'b110010010001;
   39108: result <= 12'b110010010001;
   39109: result <= 12'b110010010001;
   39110: result <= 12'b110010010001;
   39111: result <= 12'b110010010010;
   39112: result <= 12'b110010010010;
   39113: result <= 12'b110010010010;
   39114: result <= 12'b110010010010;
   39115: result <= 12'b110010010010;
   39116: result <= 12'b110010010010;
   39117: result <= 12'b110010010011;
   39118: result <= 12'b110010010011;
   39119: result <= 12'b110010010011;
   39120: result <= 12'b110010010011;
   39121: result <= 12'b110010010011;
   39122: result <= 12'b110010010011;
   39123: result <= 12'b110010010100;
   39124: result <= 12'b110010010100;
   39125: result <= 12'b110010010100;
   39126: result <= 12'b110010010100;
   39127: result <= 12'b110010010100;
   39128: result <= 12'b110010010100;
   39129: result <= 12'b110010010100;
   39130: result <= 12'b110010010101;
   39131: result <= 12'b110010010101;
   39132: result <= 12'b110010010101;
   39133: result <= 12'b110010010101;
   39134: result <= 12'b110010010101;
   39135: result <= 12'b110010010101;
   39136: result <= 12'b110010010110;
   39137: result <= 12'b110010010110;
   39138: result <= 12'b110010010110;
   39139: result <= 12'b110010010110;
   39140: result <= 12'b110010010110;
   39141: result <= 12'b110010010110;
   39142: result <= 12'b110010010111;
   39143: result <= 12'b110010010111;
   39144: result <= 12'b110010010111;
   39145: result <= 12'b110010010111;
   39146: result <= 12'b110010010111;
   39147: result <= 12'b110010010111;
   39148: result <= 12'b110010011000;
   39149: result <= 12'b110010011000;
   39150: result <= 12'b110010011000;
   39151: result <= 12'b110010011000;
   39152: result <= 12'b110010011000;
   39153: result <= 12'b110010011000;
   39154: result <= 12'b110010011001;
   39155: result <= 12'b110010011001;
   39156: result <= 12'b110010011001;
   39157: result <= 12'b110010011001;
   39158: result <= 12'b110010011001;
   39159: result <= 12'b110010011001;
   39160: result <= 12'b110010011001;
   39161: result <= 12'b110010011010;
   39162: result <= 12'b110010011010;
   39163: result <= 12'b110010011010;
   39164: result <= 12'b110010011010;
   39165: result <= 12'b110010011010;
   39166: result <= 12'b110010011010;
   39167: result <= 12'b110010011011;
   39168: result <= 12'b110010011011;
   39169: result <= 12'b110010011011;
   39170: result <= 12'b110010011011;
   39171: result <= 12'b110010011011;
   39172: result <= 12'b110010011011;
   39173: result <= 12'b110010011100;
   39174: result <= 12'b110010011100;
   39175: result <= 12'b110010011100;
   39176: result <= 12'b110010011100;
   39177: result <= 12'b110010011100;
   39178: result <= 12'b110010011100;
   39179: result <= 12'b110010011101;
   39180: result <= 12'b110010011101;
   39181: result <= 12'b110010011101;
   39182: result <= 12'b110010011101;
   39183: result <= 12'b110010011101;
   39184: result <= 12'b110010011101;
   39185: result <= 12'b110010011101;
   39186: result <= 12'b110010011110;
   39187: result <= 12'b110010011110;
   39188: result <= 12'b110010011110;
   39189: result <= 12'b110010011110;
   39190: result <= 12'b110010011110;
   39191: result <= 12'b110010011110;
   39192: result <= 12'b110010011111;
   39193: result <= 12'b110010011111;
   39194: result <= 12'b110010011111;
   39195: result <= 12'b110010011111;
   39196: result <= 12'b110010011111;
   39197: result <= 12'b110010011111;
   39198: result <= 12'b110010100000;
   39199: result <= 12'b110010100000;
   39200: result <= 12'b110010100000;
   39201: result <= 12'b110010100000;
   39202: result <= 12'b110010100000;
   39203: result <= 12'b110010100000;
   39204: result <= 12'b110010100001;
   39205: result <= 12'b110010100001;
   39206: result <= 12'b110010100001;
   39207: result <= 12'b110010100001;
   39208: result <= 12'b110010100001;
   39209: result <= 12'b110010100001;
   39210: result <= 12'b110010100001;
   39211: result <= 12'b110010100010;
   39212: result <= 12'b110010100010;
   39213: result <= 12'b110010100010;
   39214: result <= 12'b110010100010;
   39215: result <= 12'b110010100010;
   39216: result <= 12'b110010100010;
   39217: result <= 12'b110010100011;
   39218: result <= 12'b110010100011;
   39219: result <= 12'b110010100011;
   39220: result <= 12'b110010100011;
   39221: result <= 12'b110010100011;
   39222: result <= 12'b110010100011;
   39223: result <= 12'b110010100100;
   39224: result <= 12'b110010100100;
   39225: result <= 12'b110010100100;
   39226: result <= 12'b110010100100;
   39227: result <= 12'b110010100100;
   39228: result <= 12'b110010100100;
   39229: result <= 12'b110010100101;
   39230: result <= 12'b110010100101;
   39231: result <= 12'b110010100101;
   39232: result <= 12'b110010100101;
   39233: result <= 12'b110010100101;
   39234: result <= 12'b110010100101;
   39235: result <= 12'b110010100101;
   39236: result <= 12'b110010100110;
   39237: result <= 12'b110010100110;
   39238: result <= 12'b110010100110;
   39239: result <= 12'b110010100110;
   39240: result <= 12'b110010100110;
   39241: result <= 12'b110010100110;
   39242: result <= 12'b110010100111;
   39243: result <= 12'b110010100111;
   39244: result <= 12'b110010100111;
   39245: result <= 12'b110010100111;
   39246: result <= 12'b110010100111;
   39247: result <= 12'b110010100111;
   39248: result <= 12'b110010101000;
   39249: result <= 12'b110010101000;
   39250: result <= 12'b110010101000;
   39251: result <= 12'b110010101000;
   39252: result <= 12'b110010101000;
   39253: result <= 12'b110010101000;
   39254: result <= 12'b110010101001;
   39255: result <= 12'b110010101001;
   39256: result <= 12'b110010101001;
   39257: result <= 12'b110010101001;
   39258: result <= 12'b110010101001;
   39259: result <= 12'b110010101001;
   39260: result <= 12'b110010101001;
   39261: result <= 12'b110010101010;
   39262: result <= 12'b110010101010;
   39263: result <= 12'b110010101010;
   39264: result <= 12'b110010101010;
   39265: result <= 12'b110010101010;
   39266: result <= 12'b110010101010;
   39267: result <= 12'b110010101011;
   39268: result <= 12'b110010101011;
   39269: result <= 12'b110010101011;
   39270: result <= 12'b110010101011;
   39271: result <= 12'b110010101011;
   39272: result <= 12'b110010101011;
   39273: result <= 12'b110010101100;
   39274: result <= 12'b110010101100;
   39275: result <= 12'b110010101100;
   39276: result <= 12'b110010101100;
   39277: result <= 12'b110010101100;
   39278: result <= 12'b110010101100;
   39279: result <= 12'b110010101101;
   39280: result <= 12'b110010101101;
   39281: result <= 12'b110010101101;
   39282: result <= 12'b110010101101;
   39283: result <= 12'b110010101101;
   39284: result <= 12'b110010101101;
   39285: result <= 12'b110010101101;
   39286: result <= 12'b110010101110;
   39287: result <= 12'b110010101110;
   39288: result <= 12'b110010101110;
   39289: result <= 12'b110010101110;
   39290: result <= 12'b110010101110;
   39291: result <= 12'b110010101110;
   39292: result <= 12'b110010101111;
   39293: result <= 12'b110010101111;
   39294: result <= 12'b110010101111;
   39295: result <= 12'b110010101111;
   39296: result <= 12'b110010101111;
   39297: result <= 12'b110010101111;
   39298: result <= 12'b110010110000;
   39299: result <= 12'b110010110000;
   39300: result <= 12'b110010110000;
   39301: result <= 12'b110010110000;
   39302: result <= 12'b110010110000;
   39303: result <= 12'b110010110000;
   39304: result <= 12'b110010110000;
   39305: result <= 12'b110010110001;
   39306: result <= 12'b110010110001;
   39307: result <= 12'b110010110001;
   39308: result <= 12'b110010110001;
   39309: result <= 12'b110010110001;
   39310: result <= 12'b110010110001;
   39311: result <= 12'b110010110010;
   39312: result <= 12'b110010110010;
   39313: result <= 12'b110010110010;
   39314: result <= 12'b110010110010;
   39315: result <= 12'b110010110010;
   39316: result <= 12'b110010110010;
   39317: result <= 12'b110010110011;
   39318: result <= 12'b110010110011;
   39319: result <= 12'b110010110011;
   39320: result <= 12'b110010110011;
   39321: result <= 12'b110010110011;
   39322: result <= 12'b110010110011;
   39323: result <= 12'b110010110100;
   39324: result <= 12'b110010110100;
   39325: result <= 12'b110010110100;
   39326: result <= 12'b110010110100;
   39327: result <= 12'b110010110100;
   39328: result <= 12'b110010110100;
   39329: result <= 12'b110010110100;
   39330: result <= 12'b110010110101;
   39331: result <= 12'b110010110101;
   39332: result <= 12'b110010110101;
   39333: result <= 12'b110010110101;
   39334: result <= 12'b110010110101;
   39335: result <= 12'b110010110101;
   39336: result <= 12'b110010110110;
   39337: result <= 12'b110010110110;
   39338: result <= 12'b110010110110;
   39339: result <= 12'b110010110110;
   39340: result <= 12'b110010110110;
   39341: result <= 12'b110010110110;
   39342: result <= 12'b110010110111;
   39343: result <= 12'b110010110111;
   39344: result <= 12'b110010110111;
   39345: result <= 12'b110010110111;
   39346: result <= 12'b110010110111;
   39347: result <= 12'b110010110111;
   39348: result <= 12'b110010110111;
   39349: result <= 12'b110010111000;
   39350: result <= 12'b110010111000;
   39351: result <= 12'b110010111000;
   39352: result <= 12'b110010111000;
   39353: result <= 12'b110010111000;
   39354: result <= 12'b110010111000;
   39355: result <= 12'b110010111001;
   39356: result <= 12'b110010111001;
   39357: result <= 12'b110010111001;
   39358: result <= 12'b110010111001;
   39359: result <= 12'b110010111001;
   39360: result <= 12'b110010111001;
   39361: result <= 12'b110010111010;
   39362: result <= 12'b110010111010;
   39363: result <= 12'b110010111010;
   39364: result <= 12'b110010111010;
   39365: result <= 12'b110010111010;
   39366: result <= 12'b110010111010;
   39367: result <= 12'b110010111010;
   39368: result <= 12'b110010111011;
   39369: result <= 12'b110010111011;
   39370: result <= 12'b110010111011;
   39371: result <= 12'b110010111011;
   39372: result <= 12'b110010111011;
   39373: result <= 12'b110010111011;
   39374: result <= 12'b110010111100;
   39375: result <= 12'b110010111100;
   39376: result <= 12'b110010111100;
   39377: result <= 12'b110010111100;
   39378: result <= 12'b110010111100;
   39379: result <= 12'b110010111100;
   39380: result <= 12'b110010111101;
   39381: result <= 12'b110010111101;
   39382: result <= 12'b110010111101;
   39383: result <= 12'b110010111101;
   39384: result <= 12'b110010111101;
   39385: result <= 12'b110010111101;
   39386: result <= 12'b110010111101;
   39387: result <= 12'b110010111110;
   39388: result <= 12'b110010111110;
   39389: result <= 12'b110010111110;
   39390: result <= 12'b110010111110;
   39391: result <= 12'b110010111110;
   39392: result <= 12'b110010111110;
   39393: result <= 12'b110010111111;
   39394: result <= 12'b110010111111;
   39395: result <= 12'b110010111111;
   39396: result <= 12'b110010111111;
   39397: result <= 12'b110010111111;
   39398: result <= 12'b110010111111;
   39399: result <= 12'b110011000000;
   39400: result <= 12'b110011000000;
   39401: result <= 12'b110011000000;
   39402: result <= 12'b110011000000;
   39403: result <= 12'b110011000000;
   39404: result <= 12'b110011000000;
   39405: result <= 12'b110011000000;
   39406: result <= 12'b110011000001;
   39407: result <= 12'b110011000001;
   39408: result <= 12'b110011000001;
   39409: result <= 12'b110011000001;
   39410: result <= 12'b110011000001;
   39411: result <= 12'b110011000001;
   39412: result <= 12'b110011000010;
   39413: result <= 12'b110011000010;
   39414: result <= 12'b110011000010;
   39415: result <= 12'b110011000010;
   39416: result <= 12'b110011000010;
   39417: result <= 12'b110011000010;
   39418: result <= 12'b110011000011;
   39419: result <= 12'b110011000011;
   39420: result <= 12'b110011000011;
   39421: result <= 12'b110011000011;
   39422: result <= 12'b110011000011;
   39423: result <= 12'b110011000011;
   39424: result <= 12'b110011000011;
   39425: result <= 12'b110011000100;
   39426: result <= 12'b110011000100;
   39427: result <= 12'b110011000100;
   39428: result <= 12'b110011000100;
   39429: result <= 12'b110011000100;
   39430: result <= 12'b110011000100;
   39431: result <= 12'b110011000101;
   39432: result <= 12'b110011000101;
   39433: result <= 12'b110011000101;
   39434: result <= 12'b110011000101;
   39435: result <= 12'b110011000101;
   39436: result <= 12'b110011000101;
   39437: result <= 12'b110011000110;
   39438: result <= 12'b110011000110;
   39439: result <= 12'b110011000110;
   39440: result <= 12'b110011000110;
   39441: result <= 12'b110011000110;
   39442: result <= 12'b110011000110;
   39443: result <= 12'b110011000110;
   39444: result <= 12'b110011000111;
   39445: result <= 12'b110011000111;
   39446: result <= 12'b110011000111;
   39447: result <= 12'b110011000111;
   39448: result <= 12'b110011000111;
   39449: result <= 12'b110011000111;
   39450: result <= 12'b110011001000;
   39451: result <= 12'b110011001000;
   39452: result <= 12'b110011001000;
   39453: result <= 12'b110011001000;
   39454: result <= 12'b110011001000;
   39455: result <= 12'b110011001000;
   39456: result <= 12'b110011001001;
   39457: result <= 12'b110011001001;
   39458: result <= 12'b110011001001;
   39459: result <= 12'b110011001001;
   39460: result <= 12'b110011001001;
   39461: result <= 12'b110011001001;
   39462: result <= 12'b110011001001;
   39463: result <= 12'b110011001010;
   39464: result <= 12'b110011001010;
   39465: result <= 12'b110011001010;
   39466: result <= 12'b110011001010;
   39467: result <= 12'b110011001010;
   39468: result <= 12'b110011001010;
   39469: result <= 12'b110011001011;
   39470: result <= 12'b110011001011;
   39471: result <= 12'b110011001011;
   39472: result <= 12'b110011001011;
   39473: result <= 12'b110011001011;
   39474: result <= 12'b110011001011;
   39475: result <= 12'b110011001100;
   39476: result <= 12'b110011001100;
   39477: result <= 12'b110011001100;
   39478: result <= 12'b110011001100;
   39479: result <= 12'b110011001100;
   39480: result <= 12'b110011001100;
   39481: result <= 12'b110011001100;
   39482: result <= 12'b110011001101;
   39483: result <= 12'b110011001101;
   39484: result <= 12'b110011001101;
   39485: result <= 12'b110011001101;
   39486: result <= 12'b110011001101;
   39487: result <= 12'b110011001101;
   39488: result <= 12'b110011001110;
   39489: result <= 12'b110011001110;
   39490: result <= 12'b110011001110;
   39491: result <= 12'b110011001110;
   39492: result <= 12'b110011001110;
   39493: result <= 12'b110011001110;
   39494: result <= 12'b110011001111;
   39495: result <= 12'b110011001111;
   39496: result <= 12'b110011001111;
   39497: result <= 12'b110011001111;
   39498: result <= 12'b110011001111;
   39499: result <= 12'b110011001111;
   39500: result <= 12'b110011001111;
   39501: result <= 12'b110011010000;
   39502: result <= 12'b110011010000;
   39503: result <= 12'b110011010000;
   39504: result <= 12'b110011010000;
   39505: result <= 12'b110011010000;
   39506: result <= 12'b110011010000;
   39507: result <= 12'b110011010001;
   39508: result <= 12'b110011010001;
   39509: result <= 12'b110011010001;
   39510: result <= 12'b110011010001;
   39511: result <= 12'b110011010001;
   39512: result <= 12'b110011010001;
   39513: result <= 12'b110011010001;
   39514: result <= 12'b110011010010;
   39515: result <= 12'b110011010010;
   39516: result <= 12'b110011010010;
   39517: result <= 12'b110011010010;
   39518: result <= 12'b110011010010;
   39519: result <= 12'b110011010010;
   39520: result <= 12'b110011010011;
   39521: result <= 12'b110011010011;
   39522: result <= 12'b110011010011;
   39523: result <= 12'b110011010011;
   39524: result <= 12'b110011010011;
   39525: result <= 12'b110011010011;
   39526: result <= 12'b110011010100;
   39527: result <= 12'b110011010100;
   39528: result <= 12'b110011010100;
   39529: result <= 12'b110011010100;
   39530: result <= 12'b110011010100;
   39531: result <= 12'b110011010100;
   39532: result <= 12'b110011010100;
   39533: result <= 12'b110011010101;
   39534: result <= 12'b110011010101;
   39535: result <= 12'b110011010101;
   39536: result <= 12'b110011010101;
   39537: result <= 12'b110011010101;
   39538: result <= 12'b110011010101;
   39539: result <= 12'b110011010110;
   39540: result <= 12'b110011010110;
   39541: result <= 12'b110011010110;
   39542: result <= 12'b110011010110;
   39543: result <= 12'b110011010110;
   39544: result <= 12'b110011010110;
   39545: result <= 12'b110011010110;
   39546: result <= 12'b110011010111;
   39547: result <= 12'b110011010111;
   39548: result <= 12'b110011010111;
   39549: result <= 12'b110011010111;
   39550: result <= 12'b110011010111;
   39551: result <= 12'b110011010111;
   39552: result <= 12'b110011011000;
   39553: result <= 12'b110011011000;
   39554: result <= 12'b110011011000;
   39555: result <= 12'b110011011000;
   39556: result <= 12'b110011011000;
   39557: result <= 12'b110011011000;
   39558: result <= 12'b110011011001;
   39559: result <= 12'b110011011001;
   39560: result <= 12'b110011011001;
   39561: result <= 12'b110011011001;
   39562: result <= 12'b110011011001;
   39563: result <= 12'b110011011001;
   39564: result <= 12'b110011011001;
   39565: result <= 12'b110011011010;
   39566: result <= 12'b110011011010;
   39567: result <= 12'b110011011010;
   39568: result <= 12'b110011011010;
   39569: result <= 12'b110011011010;
   39570: result <= 12'b110011011010;
   39571: result <= 12'b110011011011;
   39572: result <= 12'b110011011011;
   39573: result <= 12'b110011011011;
   39574: result <= 12'b110011011011;
   39575: result <= 12'b110011011011;
   39576: result <= 12'b110011011011;
   39577: result <= 12'b110011011011;
   39578: result <= 12'b110011011100;
   39579: result <= 12'b110011011100;
   39580: result <= 12'b110011011100;
   39581: result <= 12'b110011011100;
   39582: result <= 12'b110011011100;
   39583: result <= 12'b110011011100;
   39584: result <= 12'b110011011101;
   39585: result <= 12'b110011011101;
   39586: result <= 12'b110011011101;
   39587: result <= 12'b110011011101;
   39588: result <= 12'b110011011101;
   39589: result <= 12'b110011011101;
   39590: result <= 12'b110011011110;
   39591: result <= 12'b110011011110;
   39592: result <= 12'b110011011110;
   39593: result <= 12'b110011011110;
   39594: result <= 12'b110011011110;
   39595: result <= 12'b110011011110;
   39596: result <= 12'b110011011110;
   39597: result <= 12'b110011011111;
   39598: result <= 12'b110011011111;
   39599: result <= 12'b110011011111;
   39600: result <= 12'b110011011111;
   39601: result <= 12'b110011011111;
   39602: result <= 12'b110011011111;
   39603: result <= 12'b110011100000;
   39604: result <= 12'b110011100000;
   39605: result <= 12'b110011100000;
   39606: result <= 12'b110011100000;
   39607: result <= 12'b110011100000;
   39608: result <= 12'b110011100000;
   39609: result <= 12'b110011100000;
   39610: result <= 12'b110011100001;
   39611: result <= 12'b110011100001;
   39612: result <= 12'b110011100001;
   39613: result <= 12'b110011100001;
   39614: result <= 12'b110011100001;
   39615: result <= 12'b110011100001;
   39616: result <= 12'b110011100010;
   39617: result <= 12'b110011100010;
   39618: result <= 12'b110011100010;
   39619: result <= 12'b110011100010;
   39620: result <= 12'b110011100010;
   39621: result <= 12'b110011100010;
   39622: result <= 12'b110011100010;
   39623: result <= 12'b110011100011;
   39624: result <= 12'b110011100011;
   39625: result <= 12'b110011100011;
   39626: result <= 12'b110011100011;
   39627: result <= 12'b110011100011;
   39628: result <= 12'b110011100011;
   39629: result <= 12'b110011100100;
   39630: result <= 12'b110011100100;
   39631: result <= 12'b110011100100;
   39632: result <= 12'b110011100100;
   39633: result <= 12'b110011100100;
   39634: result <= 12'b110011100100;
   39635: result <= 12'b110011100101;
   39636: result <= 12'b110011100101;
   39637: result <= 12'b110011100101;
   39638: result <= 12'b110011100101;
   39639: result <= 12'b110011100101;
   39640: result <= 12'b110011100101;
   39641: result <= 12'b110011100101;
   39642: result <= 12'b110011100110;
   39643: result <= 12'b110011100110;
   39644: result <= 12'b110011100110;
   39645: result <= 12'b110011100110;
   39646: result <= 12'b110011100110;
   39647: result <= 12'b110011100110;
   39648: result <= 12'b110011100111;
   39649: result <= 12'b110011100111;
   39650: result <= 12'b110011100111;
   39651: result <= 12'b110011100111;
   39652: result <= 12'b110011100111;
   39653: result <= 12'b110011100111;
   39654: result <= 12'b110011100111;
   39655: result <= 12'b110011101000;
   39656: result <= 12'b110011101000;
   39657: result <= 12'b110011101000;
   39658: result <= 12'b110011101000;
   39659: result <= 12'b110011101000;
   39660: result <= 12'b110011101000;
   39661: result <= 12'b110011101001;
   39662: result <= 12'b110011101001;
   39663: result <= 12'b110011101001;
   39664: result <= 12'b110011101001;
   39665: result <= 12'b110011101001;
   39666: result <= 12'b110011101001;
   39667: result <= 12'b110011101001;
   39668: result <= 12'b110011101010;
   39669: result <= 12'b110011101010;
   39670: result <= 12'b110011101010;
   39671: result <= 12'b110011101010;
   39672: result <= 12'b110011101010;
   39673: result <= 12'b110011101010;
   39674: result <= 12'b110011101011;
   39675: result <= 12'b110011101011;
   39676: result <= 12'b110011101011;
   39677: result <= 12'b110011101011;
   39678: result <= 12'b110011101011;
   39679: result <= 12'b110011101011;
   39680: result <= 12'b110011101011;
   39681: result <= 12'b110011101100;
   39682: result <= 12'b110011101100;
   39683: result <= 12'b110011101100;
   39684: result <= 12'b110011101100;
   39685: result <= 12'b110011101100;
   39686: result <= 12'b110011101100;
   39687: result <= 12'b110011101101;
   39688: result <= 12'b110011101101;
   39689: result <= 12'b110011101101;
   39690: result <= 12'b110011101101;
   39691: result <= 12'b110011101101;
   39692: result <= 12'b110011101101;
   39693: result <= 12'b110011101110;
   39694: result <= 12'b110011101110;
   39695: result <= 12'b110011101110;
   39696: result <= 12'b110011101110;
   39697: result <= 12'b110011101110;
   39698: result <= 12'b110011101110;
   39699: result <= 12'b110011101110;
   39700: result <= 12'b110011101111;
   39701: result <= 12'b110011101111;
   39702: result <= 12'b110011101111;
   39703: result <= 12'b110011101111;
   39704: result <= 12'b110011101111;
   39705: result <= 12'b110011101111;
   39706: result <= 12'b110011110000;
   39707: result <= 12'b110011110000;
   39708: result <= 12'b110011110000;
   39709: result <= 12'b110011110000;
   39710: result <= 12'b110011110000;
   39711: result <= 12'b110011110000;
   39712: result <= 12'b110011110000;
   39713: result <= 12'b110011110001;
   39714: result <= 12'b110011110001;
   39715: result <= 12'b110011110001;
   39716: result <= 12'b110011110001;
   39717: result <= 12'b110011110001;
   39718: result <= 12'b110011110001;
   39719: result <= 12'b110011110010;
   39720: result <= 12'b110011110010;
   39721: result <= 12'b110011110010;
   39722: result <= 12'b110011110010;
   39723: result <= 12'b110011110010;
   39724: result <= 12'b110011110010;
   39725: result <= 12'b110011110010;
   39726: result <= 12'b110011110011;
   39727: result <= 12'b110011110011;
   39728: result <= 12'b110011110011;
   39729: result <= 12'b110011110011;
   39730: result <= 12'b110011110011;
   39731: result <= 12'b110011110011;
   39732: result <= 12'b110011110100;
   39733: result <= 12'b110011110100;
   39734: result <= 12'b110011110100;
   39735: result <= 12'b110011110100;
   39736: result <= 12'b110011110100;
   39737: result <= 12'b110011110100;
   39738: result <= 12'b110011110100;
   39739: result <= 12'b110011110101;
   39740: result <= 12'b110011110101;
   39741: result <= 12'b110011110101;
   39742: result <= 12'b110011110101;
   39743: result <= 12'b110011110101;
   39744: result <= 12'b110011110101;
   39745: result <= 12'b110011110110;
   39746: result <= 12'b110011110110;
   39747: result <= 12'b110011110110;
   39748: result <= 12'b110011110110;
   39749: result <= 12'b110011110110;
   39750: result <= 12'b110011110110;
   39751: result <= 12'b110011110110;
   39752: result <= 12'b110011110111;
   39753: result <= 12'b110011110111;
   39754: result <= 12'b110011110111;
   39755: result <= 12'b110011110111;
   39756: result <= 12'b110011110111;
   39757: result <= 12'b110011110111;
   39758: result <= 12'b110011111000;
   39759: result <= 12'b110011111000;
   39760: result <= 12'b110011111000;
   39761: result <= 12'b110011111000;
   39762: result <= 12'b110011111000;
   39763: result <= 12'b110011111000;
   39764: result <= 12'b110011111000;
   39765: result <= 12'b110011111001;
   39766: result <= 12'b110011111001;
   39767: result <= 12'b110011111001;
   39768: result <= 12'b110011111001;
   39769: result <= 12'b110011111001;
   39770: result <= 12'b110011111001;
   39771: result <= 12'b110011111010;
   39772: result <= 12'b110011111010;
   39773: result <= 12'b110011111010;
   39774: result <= 12'b110011111010;
   39775: result <= 12'b110011111010;
   39776: result <= 12'b110011111010;
   39777: result <= 12'b110011111010;
   39778: result <= 12'b110011111011;
   39779: result <= 12'b110011111011;
   39780: result <= 12'b110011111011;
   39781: result <= 12'b110011111011;
   39782: result <= 12'b110011111011;
   39783: result <= 12'b110011111011;
   39784: result <= 12'b110011111100;
   39785: result <= 12'b110011111100;
   39786: result <= 12'b110011111100;
   39787: result <= 12'b110011111100;
   39788: result <= 12'b110011111100;
   39789: result <= 12'b110011111100;
   39790: result <= 12'b110011111100;
   39791: result <= 12'b110011111101;
   39792: result <= 12'b110011111101;
   39793: result <= 12'b110011111101;
   39794: result <= 12'b110011111101;
   39795: result <= 12'b110011111101;
   39796: result <= 12'b110011111101;
   39797: result <= 12'b110011111110;
   39798: result <= 12'b110011111110;
   39799: result <= 12'b110011111110;
   39800: result <= 12'b110011111110;
   39801: result <= 12'b110011111110;
   39802: result <= 12'b110011111110;
   39803: result <= 12'b110011111110;
   39804: result <= 12'b110011111111;
   39805: result <= 12'b110011111111;
   39806: result <= 12'b110011111111;
   39807: result <= 12'b110011111111;
   39808: result <= 12'b110011111111;
   39809: result <= 12'b110011111111;
   39810: result <= 12'b110100000000;
   39811: result <= 12'b110100000000;
   39812: result <= 12'b110100000000;
   39813: result <= 12'b110100000000;
   39814: result <= 12'b110100000000;
   39815: result <= 12'b110100000000;
   39816: result <= 12'b110100000000;
   39817: result <= 12'b110100000001;
   39818: result <= 12'b110100000001;
   39819: result <= 12'b110100000001;
   39820: result <= 12'b110100000001;
   39821: result <= 12'b110100000001;
   39822: result <= 12'b110100000001;
   39823: result <= 12'b110100000010;
   39824: result <= 12'b110100000010;
   39825: result <= 12'b110100000010;
   39826: result <= 12'b110100000010;
   39827: result <= 12'b110100000010;
   39828: result <= 12'b110100000010;
   39829: result <= 12'b110100000010;
   39830: result <= 12'b110100000011;
   39831: result <= 12'b110100000011;
   39832: result <= 12'b110100000011;
   39833: result <= 12'b110100000011;
   39834: result <= 12'b110100000011;
   39835: result <= 12'b110100000011;
   39836: result <= 12'b110100000011;
   39837: result <= 12'b110100000100;
   39838: result <= 12'b110100000100;
   39839: result <= 12'b110100000100;
   39840: result <= 12'b110100000100;
   39841: result <= 12'b110100000100;
   39842: result <= 12'b110100000100;
   39843: result <= 12'b110100000101;
   39844: result <= 12'b110100000101;
   39845: result <= 12'b110100000101;
   39846: result <= 12'b110100000101;
   39847: result <= 12'b110100000101;
   39848: result <= 12'b110100000101;
   39849: result <= 12'b110100000101;
   39850: result <= 12'b110100000110;
   39851: result <= 12'b110100000110;
   39852: result <= 12'b110100000110;
   39853: result <= 12'b110100000110;
   39854: result <= 12'b110100000110;
   39855: result <= 12'b110100000110;
   39856: result <= 12'b110100000111;
   39857: result <= 12'b110100000111;
   39858: result <= 12'b110100000111;
   39859: result <= 12'b110100000111;
   39860: result <= 12'b110100000111;
   39861: result <= 12'b110100000111;
   39862: result <= 12'b110100000111;
   39863: result <= 12'b110100001000;
   39864: result <= 12'b110100001000;
   39865: result <= 12'b110100001000;
   39866: result <= 12'b110100001000;
   39867: result <= 12'b110100001000;
   39868: result <= 12'b110100001000;
   39869: result <= 12'b110100001001;
   39870: result <= 12'b110100001001;
   39871: result <= 12'b110100001001;
   39872: result <= 12'b110100001001;
   39873: result <= 12'b110100001001;
   39874: result <= 12'b110100001001;
   39875: result <= 12'b110100001001;
   39876: result <= 12'b110100001010;
   39877: result <= 12'b110100001010;
   39878: result <= 12'b110100001010;
   39879: result <= 12'b110100001010;
   39880: result <= 12'b110100001010;
   39881: result <= 12'b110100001010;
   39882: result <= 12'b110100001011;
   39883: result <= 12'b110100001011;
   39884: result <= 12'b110100001011;
   39885: result <= 12'b110100001011;
   39886: result <= 12'b110100001011;
   39887: result <= 12'b110100001011;
   39888: result <= 12'b110100001011;
   39889: result <= 12'b110100001100;
   39890: result <= 12'b110100001100;
   39891: result <= 12'b110100001100;
   39892: result <= 12'b110100001100;
   39893: result <= 12'b110100001100;
   39894: result <= 12'b110100001100;
   39895: result <= 12'b110100001101;
   39896: result <= 12'b110100001101;
   39897: result <= 12'b110100001101;
   39898: result <= 12'b110100001101;
   39899: result <= 12'b110100001101;
   39900: result <= 12'b110100001101;
   39901: result <= 12'b110100001101;
   39902: result <= 12'b110100001110;
   39903: result <= 12'b110100001110;
   39904: result <= 12'b110100001110;
   39905: result <= 12'b110100001110;
   39906: result <= 12'b110100001110;
   39907: result <= 12'b110100001110;
   39908: result <= 12'b110100001110;
   39909: result <= 12'b110100001111;
   39910: result <= 12'b110100001111;
   39911: result <= 12'b110100001111;
   39912: result <= 12'b110100001111;
   39913: result <= 12'b110100001111;
   39914: result <= 12'b110100001111;
   39915: result <= 12'b110100010000;
   39916: result <= 12'b110100010000;
   39917: result <= 12'b110100010000;
   39918: result <= 12'b110100010000;
   39919: result <= 12'b110100010000;
   39920: result <= 12'b110100010000;
   39921: result <= 12'b110100010000;
   39922: result <= 12'b110100010001;
   39923: result <= 12'b110100010001;
   39924: result <= 12'b110100010001;
   39925: result <= 12'b110100010001;
   39926: result <= 12'b110100010001;
   39927: result <= 12'b110100010001;
   39928: result <= 12'b110100010010;
   39929: result <= 12'b110100010010;
   39930: result <= 12'b110100010010;
   39931: result <= 12'b110100010010;
   39932: result <= 12'b110100010010;
   39933: result <= 12'b110100010010;
   39934: result <= 12'b110100010010;
   39935: result <= 12'b110100010011;
   39936: result <= 12'b110100010011;
   39937: result <= 12'b110100010011;
   39938: result <= 12'b110100010011;
   39939: result <= 12'b110100010011;
   39940: result <= 12'b110100010011;
   39941: result <= 12'b110100010011;
   39942: result <= 12'b110100010100;
   39943: result <= 12'b110100010100;
   39944: result <= 12'b110100010100;
   39945: result <= 12'b110100010100;
   39946: result <= 12'b110100010100;
   39947: result <= 12'b110100010100;
   39948: result <= 12'b110100010101;
   39949: result <= 12'b110100010101;
   39950: result <= 12'b110100010101;
   39951: result <= 12'b110100010101;
   39952: result <= 12'b110100010101;
   39953: result <= 12'b110100010101;
   39954: result <= 12'b110100010101;
   39955: result <= 12'b110100010110;
   39956: result <= 12'b110100010110;
   39957: result <= 12'b110100010110;
   39958: result <= 12'b110100010110;
   39959: result <= 12'b110100010110;
   39960: result <= 12'b110100010110;
   39961: result <= 12'b110100010111;
   39962: result <= 12'b110100010111;
   39963: result <= 12'b110100010111;
   39964: result <= 12'b110100010111;
   39965: result <= 12'b110100010111;
   39966: result <= 12'b110100010111;
   39967: result <= 12'b110100010111;
   39968: result <= 12'b110100011000;
   39969: result <= 12'b110100011000;
   39970: result <= 12'b110100011000;
   39971: result <= 12'b110100011000;
   39972: result <= 12'b110100011000;
   39973: result <= 12'b110100011000;
   39974: result <= 12'b110100011000;
   39975: result <= 12'b110100011001;
   39976: result <= 12'b110100011001;
   39977: result <= 12'b110100011001;
   39978: result <= 12'b110100011001;
   39979: result <= 12'b110100011001;
   39980: result <= 12'b110100011001;
   39981: result <= 12'b110100011010;
   39982: result <= 12'b110100011010;
   39983: result <= 12'b110100011010;
   39984: result <= 12'b110100011010;
   39985: result <= 12'b110100011010;
   39986: result <= 12'b110100011010;
   39987: result <= 12'b110100011010;
   39988: result <= 12'b110100011011;
   39989: result <= 12'b110100011011;
   39990: result <= 12'b110100011011;
   39991: result <= 12'b110100011011;
   39992: result <= 12'b110100011011;
   39993: result <= 12'b110100011011;
   39994: result <= 12'b110100011100;
   39995: result <= 12'b110100011100;
   39996: result <= 12'b110100011100;
   39997: result <= 12'b110100011100;
   39998: result <= 12'b110100011100;
   39999: result <= 12'b110100011100;
   40000: result <= 12'b110100011100;
   40001: result <= 12'b110100011101;
   40002: result <= 12'b110100011101;
   40003: result <= 12'b110100011101;
   40004: result <= 12'b110100011101;
   40005: result <= 12'b110100011101;
   40006: result <= 12'b110100011101;
   40007: result <= 12'b110100011101;
   40008: result <= 12'b110100011110;
   40009: result <= 12'b110100011110;
   40010: result <= 12'b110100011110;
   40011: result <= 12'b110100011110;
   40012: result <= 12'b110100011110;
   40013: result <= 12'b110100011110;
   40014: result <= 12'b110100011111;
   40015: result <= 12'b110100011111;
   40016: result <= 12'b110100011111;
   40017: result <= 12'b110100011111;
   40018: result <= 12'b110100011111;
   40019: result <= 12'b110100011111;
   40020: result <= 12'b110100011111;
   40021: result <= 12'b110100100000;
   40022: result <= 12'b110100100000;
   40023: result <= 12'b110100100000;
   40024: result <= 12'b110100100000;
   40025: result <= 12'b110100100000;
   40026: result <= 12'b110100100000;
   40027: result <= 12'b110100100000;
   40028: result <= 12'b110100100001;
   40029: result <= 12'b110100100001;
   40030: result <= 12'b110100100001;
   40031: result <= 12'b110100100001;
   40032: result <= 12'b110100100001;
   40033: result <= 12'b110100100001;
   40034: result <= 12'b110100100010;
   40035: result <= 12'b110100100010;
   40036: result <= 12'b110100100010;
   40037: result <= 12'b110100100010;
   40038: result <= 12'b110100100010;
   40039: result <= 12'b110100100010;
   40040: result <= 12'b110100100010;
   40041: result <= 12'b110100100011;
   40042: result <= 12'b110100100011;
   40043: result <= 12'b110100100011;
   40044: result <= 12'b110100100011;
   40045: result <= 12'b110100100011;
   40046: result <= 12'b110100100011;
   40047: result <= 12'b110100100100;
   40048: result <= 12'b110100100100;
   40049: result <= 12'b110100100100;
   40050: result <= 12'b110100100100;
   40051: result <= 12'b110100100100;
   40052: result <= 12'b110100100100;
   40053: result <= 12'b110100100100;
   40054: result <= 12'b110100100101;
   40055: result <= 12'b110100100101;
   40056: result <= 12'b110100100101;
   40057: result <= 12'b110100100101;
   40058: result <= 12'b110100100101;
   40059: result <= 12'b110100100101;
   40060: result <= 12'b110100100101;
   40061: result <= 12'b110100100110;
   40062: result <= 12'b110100100110;
   40063: result <= 12'b110100100110;
   40064: result <= 12'b110100100110;
   40065: result <= 12'b110100100110;
   40066: result <= 12'b110100100110;
   40067: result <= 12'b110100100111;
   40068: result <= 12'b110100100111;
   40069: result <= 12'b110100100111;
   40070: result <= 12'b110100100111;
   40071: result <= 12'b110100100111;
   40072: result <= 12'b110100100111;
   40073: result <= 12'b110100100111;
   40074: result <= 12'b110100101000;
   40075: result <= 12'b110100101000;
   40076: result <= 12'b110100101000;
   40077: result <= 12'b110100101000;
   40078: result <= 12'b110100101000;
   40079: result <= 12'b110100101000;
   40080: result <= 12'b110100101000;
   40081: result <= 12'b110100101001;
   40082: result <= 12'b110100101001;
   40083: result <= 12'b110100101001;
   40084: result <= 12'b110100101001;
   40085: result <= 12'b110100101001;
   40086: result <= 12'b110100101001;
   40087: result <= 12'b110100101010;
   40088: result <= 12'b110100101010;
   40089: result <= 12'b110100101010;
   40090: result <= 12'b110100101010;
   40091: result <= 12'b110100101010;
   40092: result <= 12'b110100101010;
   40093: result <= 12'b110100101010;
   40094: result <= 12'b110100101011;
   40095: result <= 12'b110100101011;
   40096: result <= 12'b110100101011;
   40097: result <= 12'b110100101011;
   40098: result <= 12'b110100101011;
   40099: result <= 12'b110100101011;
   40100: result <= 12'b110100101011;
   40101: result <= 12'b110100101100;
   40102: result <= 12'b110100101100;
   40103: result <= 12'b110100101100;
   40104: result <= 12'b110100101100;
   40105: result <= 12'b110100101100;
   40106: result <= 12'b110100101100;
   40107: result <= 12'b110100101101;
   40108: result <= 12'b110100101101;
   40109: result <= 12'b110100101101;
   40110: result <= 12'b110100101101;
   40111: result <= 12'b110100101101;
   40112: result <= 12'b110100101101;
   40113: result <= 12'b110100101101;
   40114: result <= 12'b110100101110;
   40115: result <= 12'b110100101110;
   40116: result <= 12'b110100101110;
   40117: result <= 12'b110100101110;
   40118: result <= 12'b110100101110;
   40119: result <= 12'b110100101110;
   40120: result <= 12'b110100101110;
   40121: result <= 12'b110100101111;
   40122: result <= 12'b110100101111;
   40123: result <= 12'b110100101111;
   40124: result <= 12'b110100101111;
   40125: result <= 12'b110100101111;
   40126: result <= 12'b110100101111;
   40127: result <= 12'b110100110000;
   40128: result <= 12'b110100110000;
   40129: result <= 12'b110100110000;
   40130: result <= 12'b110100110000;
   40131: result <= 12'b110100110000;
   40132: result <= 12'b110100110000;
   40133: result <= 12'b110100110000;
   40134: result <= 12'b110100110001;
   40135: result <= 12'b110100110001;
   40136: result <= 12'b110100110001;
   40137: result <= 12'b110100110001;
   40138: result <= 12'b110100110001;
   40139: result <= 12'b110100110001;
   40140: result <= 12'b110100110001;
   40141: result <= 12'b110100110010;
   40142: result <= 12'b110100110010;
   40143: result <= 12'b110100110010;
   40144: result <= 12'b110100110010;
   40145: result <= 12'b110100110010;
   40146: result <= 12'b110100110010;
   40147: result <= 12'b110100110010;
   40148: result <= 12'b110100110011;
   40149: result <= 12'b110100110011;
   40150: result <= 12'b110100110011;
   40151: result <= 12'b110100110011;
   40152: result <= 12'b110100110011;
   40153: result <= 12'b110100110011;
   40154: result <= 12'b110100110100;
   40155: result <= 12'b110100110100;
   40156: result <= 12'b110100110100;
   40157: result <= 12'b110100110100;
   40158: result <= 12'b110100110100;
   40159: result <= 12'b110100110100;
   40160: result <= 12'b110100110100;
   40161: result <= 12'b110100110101;
   40162: result <= 12'b110100110101;
   40163: result <= 12'b110100110101;
   40164: result <= 12'b110100110101;
   40165: result <= 12'b110100110101;
   40166: result <= 12'b110100110101;
   40167: result <= 12'b110100110101;
   40168: result <= 12'b110100110110;
   40169: result <= 12'b110100110110;
   40170: result <= 12'b110100110110;
   40171: result <= 12'b110100110110;
   40172: result <= 12'b110100110110;
   40173: result <= 12'b110100110110;
   40174: result <= 12'b110100110111;
   40175: result <= 12'b110100110111;
   40176: result <= 12'b110100110111;
   40177: result <= 12'b110100110111;
   40178: result <= 12'b110100110111;
   40179: result <= 12'b110100110111;
   40180: result <= 12'b110100110111;
   40181: result <= 12'b110100111000;
   40182: result <= 12'b110100111000;
   40183: result <= 12'b110100111000;
   40184: result <= 12'b110100111000;
   40185: result <= 12'b110100111000;
   40186: result <= 12'b110100111000;
   40187: result <= 12'b110100111000;
   40188: result <= 12'b110100111001;
   40189: result <= 12'b110100111001;
   40190: result <= 12'b110100111001;
   40191: result <= 12'b110100111001;
   40192: result <= 12'b110100111001;
   40193: result <= 12'b110100111001;
   40194: result <= 12'b110100111001;
   40195: result <= 12'b110100111010;
   40196: result <= 12'b110100111010;
   40197: result <= 12'b110100111010;
   40198: result <= 12'b110100111010;
   40199: result <= 12'b110100111010;
   40200: result <= 12'b110100111010;
   40201: result <= 12'b110100111011;
   40202: result <= 12'b110100111011;
   40203: result <= 12'b110100111011;
   40204: result <= 12'b110100111011;
   40205: result <= 12'b110100111011;
   40206: result <= 12'b110100111011;
   40207: result <= 12'b110100111011;
   40208: result <= 12'b110100111100;
   40209: result <= 12'b110100111100;
   40210: result <= 12'b110100111100;
   40211: result <= 12'b110100111100;
   40212: result <= 12'b110100111100;
   40213: result <= 12'b110100111100;
   40214: result <= 12'b110100111100;
   40215: result <= 12'b110100111101;
   40216: result <= 12'b110100111101;
   40217: result <= 12'b110100111101;
   40218: result <= 12'b110100111101;
   40219: result <= 12'b110100111101;
   40220: result <= 12'b110100111101;
   40221: result <= 12'b110100111110;
   40222: result <= 12'b110100111110;
   40223: result <= 12'b110100111110;
   40224: result <= 12'b110100111110;
   40225: result <= 12'b110100111110;
   40226: result <= 12'b110100111110;
   40227: result <= 12'b110100111110;
   40228: result <= 12'b110100111111;
   40229: result <= 12'b110100111111;
   40230: result <= 12'b110100111111;
   40231: result <= 12'b110100111111;
   40232: result <= 12'b110100111111;
   40233: result <= 12'b110100111111;
   40234: result <= 12'b110100111111;
   40235: result <= 12'b110101000000;
   40236: result <= 12'b110101000000;
   40237: result <= 12'b110101000000;
   40238: result <= 12'b110101000000;
   40239: result <= 12'b110101000000;
   40240: result <= 12'b110101000000;
   40241: result <= 12'b110101000000;
   40242: result <= 12'b110101000001;
   40243: result <= 12'b110101000001;
   40244: result <= 12'b110101000001;
   40245: result <= 12'b110101000001;
   40246: result <= 12'b110101000001;
   40247: result <= 12'b110101000001;
   40248: result <= 12'b110101000010;
   40249: result <= 12'b110101000010;
   40250: result <= 12'b110101000010;
   40251: result <= 12'b110101000010;
   40252: result <= 12'b110101000010;
   40253: result <= 12'b110101000010;
   40254: result <= 12'b110101000010;
   40255: result <= 12'b110101000011;
   40256: result <= 12'b110101000011;
   40257: result <= 12'b110101000011;
   40258: result <= 12'b110101000011;
   40259: result <= 12'b110101000011;
   40260: result <= 12'b110101000011;
   40261: result <= 12'b110101000011;
   40262: result <= 12'b110101000100;
   40263: result <= 12'b110101000100;
   40264: result <= 12'b110101000100;
   40265: result <= 12'b110101000100;
   40266: result <= 12'b110101000100;
   40267: result <= 12'b110101000100;
   40268: result <= 12'b110101000100;
   40269: result <= 12'b110101000101;
   40270: result <= 12'b110101000101;
   40271: result <= 12'b110101000101;
   40272: result <= 12'b110101000101;
   40273: result <= 12'b110101000101;
   40274: result <= 12'b110101000101;
   40275: result <= 12'b110101000101;
   40276: result <= 12'b110101000110;
   40277: result <= 12'b110101000110;
   40278: result <= 12'b110101000110;
   40279: result <= 12'b110101000110;
   40280: result <= 12'b110101000110;
   40281: result <= 12'b110101000110;
   40282: result <= 12'b110101000111;
   40283: result <= 12'b110101000111;
   40284: result <= 12'b110101000111;
   40285: result <= 12'b110101000111;
   40286: result <= 12'b110101000111;
   40287: result <= 12'b110101000111;
   40288: result <= 12'b110101000111;
   40289: result <= 12'b110101001000;
   40290: result <= 12'b110101001000;
   40291: result <= 12'b110101001000;
   40292: result <= 12'b110101001000;
   40293: result <= 12'b110101001000;
   40294: result <= 12'b110101001000;
   40295: result <= 12'b110101001000;
   40296: result <= 12'b110101001001;
   40297: result <= 12'b110101001001;
   40298: result <= 12'b110101001001;
   40299: result <= 12'b110101001001;
   40300: result <= 12'b110101001001;
   40301: result <= 12'b110101001001;
   40302: result <= 12'b110101001001;
   40303: result <= 12'b110101001010;
   40304: result <= 12'b110101001010;
   40305: result <= 12'b110101001010;
   40306: result <= 12'b110101001010;
   40307: result <= 12'b110101001010;
   40308: result <= 12'b110101001010;
   40309: result <= 12'b110101001011;
   40310: result <= 12'b110101001011;
   40311: result <= 12'b110101001011;
   40312: result <= 12'b110101001011;
   40313: result <= 12'b110101001011;
   40314: result <= 12'b110101001011;
   40315: result <= 12'b110101001011;
   40316: result <= 12'b110101001100;
   40317: result <= 12'b110101001100;
   40318: result <= 12'b110101001100;
   40319: result <= 12'b110101001100;
   40320: result <= 12'b110101001100;
   40321: result <= 12'b110101001100;
   40322: result <= 12'b110101001100;
   40323: result <= 12'b110101001101;
   40324: result <= 12'b110101001101;
   40325: result <= 12'b110101001101;
   40326: result <= 12'b110101001101;
   40327: result <= 12'b110101001101;
   40328: result <= 12'b110101001101;
   40329: result <= 12'b110101001101;
   40330: result <= 12'b110101001110;
   40331: result <= 12'b110101001110;
   40332: result <= 12'b110101001110;
   40333: result <= 12'b110101001110;
   40334: result <= 12'b110101001110;
   40335: result <= 12'b110101001110;
   40336: result <= 12'b110101001110;
   40337: result <= 12'b110101001111;
   40338: result <= 12'b110101001111;
   40339: result <= 12'b110101001111;
   40340: result <= 12'b110101001111;
   40341: result <= 12'b110101001111;
   40342: result <= 12'b110101001111;
   40343: result <= 12'b110101010000;
   40344: result <= 12'b110101010000;
   40345: result <= 12'b110101010000;
   40346: result <= 12'b110101010000;
   40347: result <= 12'b110101010000;
   40348: result <= 12'b110101010000;
   40349: result <= 12'b110101010000;
   40350: result <= 12'b110101010001;
   40351: result <= 12'b110101010001;
   40352: result <= 12'b110101010001;
   40353: result <= 12'b110101010001;
   40354: result <= 12'b110101010001;
   40355: result <= 12'b110101010001;
   40356: result <= 12'b110101010001;
   40357: result <= 12'b110101010010;
   40358: result <= 12'b110101010010;
   40359: result <= 12'b110101010010;
   40360: result <= 12'b110101010010;
   40361: result <= 12'b110101010010;
   40362: result <= 12'b110101010010;
   40363: result <= 12'b110101010010;
   40364: result <= 12'b110101010011;
   40365: result <= 12'b110101010011;
   40366: result <= 12'b110101010011;
   40367: result <= 12'b110101010011;
   40368: result <= 12'b110101010011;
   40369: result <= 12'b110101010011;
   40370: result <= 12'b110101010011;
   40371: result <= 12'b110101010100;
   40372: result <= 12'b110101010100;
   40373: result <= 12'b110101010100;
   40374: result <= 12'b110101010100;
   40375: result <= 12'b110101010100;
   40376: result <= 12'b110101010100;
   40377: result <= 12'b110101010100;
   40378: result <= 12'b110101010101;
   40379: result <= 12'b110101010101;
   40380: result <= 12'b110101010101;
   40381: result <= 12'b110101010101;
   40382: result <= 12'b110101010101;
   40383: result <= 12'b110101010101;
   40384: result <= 12'b110101010110;
   40385: result <= 12'b110101010110;
   40386: result <= 12'b110101010110;
   40387: result <= 12'b110101010110;
   40388: result <= 12'b110101010110;
   40389: result <= 12'b110101010110;
   40390: result <= 12'b110101010110;
   40391: result <= 12'b110101010111;
   40392: result <= 12'b110101010111;
   40393: result <= 12'b110101010111;
   40394: result <= 12'b110101010111;
   40395: result <= 12'b110101010111;
   40396: result <= 12'b110101010111;
   40397: result <= 12'b110101010111;
   40398: result <= 12'b110101011000;
   40399: result <= 12'b110101011000;
   40400: result <= 12'b110101011000;
   40401: result <= 12'b110101011000;
   40402: result <= 12'b110101011000;
   40403: result <= 12'b110101011000;
   40404: result <= 12'b110101011000;
   40405: result <= 12'b110101011001;
   40406: result <= 12'b110101011001;
   40407: result <= 12'b110101011001;
   40408: result <= 12'b110101011001;
   40409: result <= 12'b110101011001;
   40410: result <= 12'b110101011001;
   40411: result <= 12'b110101011001;
   40412: result <= 12'b110101011010;
   40413: result <= 12'b110101011010;
   40414: result <= 12'b110101011010;
   40415: result <= 12'b110101011010;
   40416: result <= 12'b110101011010;
   40417: result <= 12'b110101011010;
   40418: result <= 12'b110101011010;
   40419: result <= 12'b110101011011;
   40420: result <= 12'b110101011011;
   40421: result <= 12'b110101011011;
   40422: result <= 12'b110101011011;
   40423: result <= 12'b110101011011;
   40424: result <= 12'b110101011011;
   40425: result <= 12'b110101011100;
   40426: result <= 12'b110101011100;
   40427: result <= 12'b110101011100;
   40428: result <= 12'b110101011100;
   40429: result <= 12'b110101011100;
   40430: result <= 12'b110101011100;
   40431: result <= 12'b110101011100;
   40432: result <= 12'b110101011101;
   40433: result <= 12'b110101011101;
   40434: result <= 12'b110101011101;
   40435: result <= 12'b110101011101;
   40436: result <= 12'b110101011101;
   40437: result <= 12'b110101011101;
   40438: result <= 12'b110101011101;
   40439: result <= 12'b110101011110;
   40440: result <= 12'b110101011110;
   40441: result <= 12'b110101011110;
   40442: result <= 12'b110101011110;
   40443: result <= 12'b110101011110;
   40444: result <= 12'b110101011110;
   40445: result <= 12'b110101011110;
   40446: result <= 12'b110101011111;
   40447: result <= 12'b110101011111;
   40448: result <= 12'b110101011111;
   40449: result <= 12'b110101011111;
   40450: result <= 12'b110101011111;
   40451: result <= 12'b110101011111;
   40452: result <= 12'b110101011111;
   40453: result <= 12'b110101100000;
   40454: result <= 12'b110101100000;
   40455: result <= 12'b110101100000;
   40456: result <= 12'b110101100000;
   40457: result <= 12'b110101100000;
   40458: result <= 12'b110101100000;
   40459: result <= 12'b110101100000;
   40460: result <= 12'b110101100001;
   40461: result <= 12'b110101100001;
   40462: result <= 12'b110101100001;
   40463: result <= 12'b110101100001;
   40464: result <= 12'b110101100001;
   40465: result <= 12'b110101100001;
   40466: result <= 12'b110101100001;
   40467: result <= 12'b110101100010;
   40468: result <= 12'b110101100010;
   40469: result <= 12'b110101100010;
   40470: result <= 12'b110101100010;
   40471: result <= 12'b110101100010;
   40472: result <= 12'b110101100010;
   40473: result <= 12'b110101100010;
   40474: result <= 12'b110101100011;
   40475: result <= 12'b110101100011;
   40476: result <= 12'b110101100011;
   40477: result <= 12'b110101100011;
   40478: result <= 12'b110101100011;
   40479: result <= 12'b110101100011;
   40480: result <= 12'b110101100100;
   40481: result <= 12'b110101100100;
   40482: result <= 12'b110101100100;
   40483: result <= 12'b110101100100;
   40484: result <= 12'b110101100100;
   40485: result <= 12'b110101100100;
   40486: result <= 12'b110101100100;
   40487: result <= 12'b110101100101;
   40488: result <= 12'b110101100101;
   40489: result <= 12'b110101100101;
   40490: result <= 12'b110101100101;
   40491: result <= 12'b110101100101;
   40492: result <= 12'b110101100101;
   40493: result <= 12'b110101100101;
   40494: result <= 12'b110101100110;
   40495: result <= 12'b110101100110;
   40496: result <= 12'b110101100110;
   40497: result <= 12'b110101100110;
   40498: result <= 12'b110101100110;
   40499: result <= 12'b110101100110;
   40500: result <= 12'b110101100110;
   40501: result <= 12'b110101100111;
   40502: result <= 12'b110101100111;
   40503: result <= 12'b110101100111;
   40504: result <= 12'b110101100111;
   40505: result <= 12'b110101100111;
   40506: result <= 12'b110101100111;
   40507: result <= 12'b110101100111;
   40508: result <= 12'b110101101000;
   40509: result <= 12'b110101101000;
   40510: result <= 12'b110101101000;
   40511: result <= 12'b110101101000;
   40512: result <= 12'b110101101000;
   40513: result <= 12'b110101101000;
   40514: result <= 12'b110101101000;
   40515: result <= 12'b110101101001;
   40516: result <= 12'b110101101001;
   40517: result <= 12'b110101101001;
   40518: result <= 12'b110101101001;
   40519: result <= 12'b110101101001;
   40520: result <= 12'b110101101001;
   40521: result <= 12'b110101101001;
   40522: result <= 12'b110101101010;
   40523: result <= 12'b110101101010;
   40524: result <= 12'b110101101010;
   40525: result <= 12'b110101101010;
   40526: result <= 12'b110101101010;
   40527: result <= 12'b110101101010;
   40528: result <= 12'b110101101010;
   40529: result <= 12'b110101101011;
   40530: result <= 12'b110101101011;
   40531: result <= 12'b110101101011;
   40532: result <= 12'b110101101011;
   40533: result <= 12'b110101101011;
   40534: result <= 12'b110101101011;
   40535: result <= 12'b110101101011;
   40536: result <= 12'b110101101100;
   40537: result <= 12'b110101101100;
   40538: result <= 12'b110101101100;
   40539: result <= 12'b110101101100;
   40540: result <= 12'b110101101100;
   40541: result <= 12'b110101101100;
   40542: result <= 12'b110101101100;
   40543: result <= 12'b110101101101;
   40544: result <= 12'b110101101101;
   40545: result <= 12'b110101101101;
   40546: result <= 12'b110101101101;
   40547: result <= 12'b110101101101;
   40548: result <= 12'b110101101101;
   40549: result <= 12'b110101101101;
   40550: result <= 12'b110101101110;
   40551: result <= 12'b110101101110;
   40552: result <= 12'b110101101110;
   40553: result <= 12'b110101101110;
   40554: result <= 12'b110101101110;
   40555: result <= 12'b110101101110;
   40556: result <= 12'b110101101110;
   40557: result <= 12'b110101101111;
   40558: result <= 12'b110101101111;
   40559: result <= 12'b110101101111;
   40560: result <= 12'b110101101111;
   40561: result <= 12'b110101101111;
   40562: result <= 12'b110101101111;
   40563: result <= 12'b110101101111;
   40564: result <= 12'b110101110000;
   40565: result <= 12'b110101110000;
   40566: result <= 12'b110101110000;
   40567: result <= 12'b110101110000;
   40568: result <= 12'b110101110000;
   40569: result <= 12'b110101110000;
   40570: result <= 12'b110101110001;
   40571: result <= 12'b110101110001;
   40572: result <= 12'b110101110001;
   40573: result <= 12'b110101110001;
   40574: result <= 12'b110101110001;
   40575: result <= 12'b110101110001;
   40576: result <= 12'b110101110001;
   40577: result <= 12'b110101110010;
   40578: result <= 12'b110101110010;
   40579: result <= 12'b110101110010;
   40580: result <= 12'b110101110010;
   40581: result <= 12'b110101110010;
   40582: result <= 12'b110101110010;
   40583: result <= 12'b110101110010;
   40584: result <= 12'b110101110011;
   40585: result <= 12'b110101110011;
   40586: result <= 12'b110101110011;
   40587: result <= 12'b110101110011;
   40588: result <= 12'b110101110011;
   40589: result <= 12'b110101110011;
   40590: result <= 12'b110101110011;
   40591: result <= 12'b110101110100;
   40592: result <= 12'b110101110100;
   40593: result <= 12'b110101110100;
   40594: result <= 12'b110101110100;
   40595: result <= 12'b110101110100;
   40596: result <= 12'b110101110100;
   40597: result <= 12'b110101110100;
   40598: result <= 12'b110101110101;
   40599: result <= 12'b110101110101;
   40600: result <= 12'b110101110101;
   40601: result <= 12'b110101110101;
   40602: result <= 12'b110101110101;
   40603: result <= 12'b110101110101;
   40604: result <= 12'b110101110101;
   40605: result <= 12'b110101110110;
   40606: result <= 12'b110101110110;
   40607: result <= 12'b110101110110;
   40608: result <= 12'b110101110110;
   40609: result <= 12'b110101110110;
   40610: result <= 12'b110101110110;
   40611: result <= 12'b110101110110;
   40612: result <= 12'b110101110111;
   40613: result <= 12'b110101110111;
   40614: result <= 12'b110101110111;
   40615: result <= 12'b110101110111;
   40616: result <= 12'b110101110111;
   40617: result <= 12'b110101110111;
   40618: result <= 12'b110101110111;
   40619: result <= 12'b110101111000;
   40620: result <= 12'b110101111000;
   40621: result <= 12'b110101111000;
   40622: result <= 12'b110101111000;
   40623: result <= 12'b110101111000;
   40624: result <= 12'b110101111000;
   40625: result <= 12'b110101111000;
   40626: result <= 12'b110101111001;
   40627: result <= 12'b110101111001;
   40628: result <= 12'b110101111001;
   40629: result <= 12'b110101111001;
   40630: result <= 12'b110101111001;
   40631: result <= 12'b110101111001;
   40632: result <= 12'b110101111001;
   40633: result <= 12'b110101111010;
   40634: result <= 12'b110101111010;
   40635: result <= 12'b110101111010;
   40636: result <= 12'b110101111010;
   40637: result <= 12'b110101111010;
   40638: result <= 12'b110101111010;
   40639: result <= 12'b110101111010;
   40640: result <= 12'b110101111011;
   40641: result <= 12'b110101111011;
   40642: result <= 12'b110101111011;
   40643: result <= 12'b110101111011;
   40644: result <= 12'b110101111011;
   40645: result <= 12'b110101111011;
   40646: result <= 12'b110101111011;
   40647: result <= 12'b110101111100;
   40648: result <= 12'b110101111100;
   40649: result <= 12'b110101111100;
   40650: result <= 12'b110101111100;
   40651: result <= 12'b110101111100;
   40652: result <= 12'b110101111100;
   40653: result <= 12'b110101111100;
   40654: result <= 12'b110101111101;
   40655: result <= 12'b110101111101;
   40656: result <= 12'b110101111101;
   40657: result <= 12'b110101111101;
   40658: result <= 12'b110101111101;
   40659: result <= 12'b110101111101;
   40660: result <= 12'b110101111101;
   40661: result <= 12'b110101111110;
   40662: result <= 12'b110101111110;
   40663: result <= 12'b110101111110;
   40664: result <= 12'b110101111110;
   40665: result <= 12'b110101111110;
   40666: result <= 12'b110101111110;
   40667: result <= 12'b110101111110;
   40668: result <= 12'b110101111111;
   40669: result <= 12'b110101111111;
   40670: result <= 12'b110101111111;
   40671: result <= 12'b110101111111;
   40672: result <= 12'b110101111111;
   40673: result <= 12'b110101111111;
   40674: result <= 12'b110101111111;
   40675: result <= 12'b110110000000;
   40676: result <= 12'b110110000000;
   40677: result <= 12'b110110000000;
   40678: result <= 12'b110110000000;
   40679: result <= 12'b110110000000;
   40680: result <= 12'b110110000000;
   40681: result <= 12'b110110000000;
   40682: result <= 12'b110110000001;
   40683: result <= 12'b110110000001;
   40684: result <= 12'b110110000001;
   40685: result <= 12'b110110000001;
   40686: result <= 12'b110110000001;
   40687: result <= 12'b110110000001;
   40688: result <= 12'b110110000001;
   40689: result <= 12'b110110000010;
   40690: result <= 12'b110110000010;
   40691: result <= 12'b110110000010;
   40692: result <= 12'b110110000010;
   40693: result <= 12'b110110000010;
   40694: result <= 12'b110110000010;
   40695: result <= 12'b110110000010;
   40696: result <= 12'b110110000011;
   40697: result <= 12'b110110000011;
   40698: result <= 12'b110110000011;
   40699: result <= 12'b110110000011;
   40700: result <= 12'b110110000011;
   40701: result <= 12'b110110000011;
   40702: result <= 12'b110110000011;
   40703: result <= 12'b110110000100;
   40704: result <= 12'b110110000100;
   40705: result <= 12'b110110000100;
   40706: result <= 12'b110110000100;
   40707: result <= 12'b110110000100;
   40708: result <= 12'b110110000100;
   40709: result <= 12'b110110000100;
   40710: result <= 12'b110110000101;
   40711: result <= 12'b110110000101;
   40712: result <= 12'b110110000101;
   40713: result <= 12'b110110000101;
   40714: result <= 12'b110110000101;
   40715: result <= 12'b110110000101;
   40716: result <= 12'b110110000101;
   40717: result <= 12'b110110000110;
   40718: result <= 12'b110110000110;
   40719: result <= 12'b110110000110;
   40720: result <= 12'b110110000110;
   40721: result <= 12'b110110000110;
   40722: result <= 12'b110110000110;
   40723: result <= 12'b110110000110;
   40724: result <= 12'b110110000111;
   40725: result <= 12'b110110000111;
   40726: result <= 12'b110110000111;
   40727: result <= 12'b110110000111;
   40728: result <= 12'b110110000111;
   40729: result <= 12'b110110000111;
   40730: result <= 12'b110110000111;
   40731: result <= 12'b110110001000;
   40732: result <= 12'b110110001000;
   40733: result <= 12'b110110001000;
   40734: result <= 12'b110110001000;
   40735: result <= 12'b110110001000;
   40736: result <= 12'b110110001000;
   40737: result <= 12'b110110001000;
   40738: result <= 12'b110110001001;
   40739: result <= 12'b110110001001;
   40740: result <= 12'b110110001001;
   40741: result <= 12'b110110001001;
   40742: result <= 12'b110110001001;
   40743: result <= 12'b110110001001;
   40744: result <= 12'b110110001001;
   40745: result <= 12'b110110001001;
   40746: result <= 12'b110110001010;
   40747: result <= 12'b110110001010;
   40748: result <= 12'b110110001010;
   40749: result <= 12'b110110001010;
   40750: result <= 12'b110110001010;
   40751: result <= 12'b110110001010;
   40752: result <= 12'b110110001010;
   40753: result <= 12'b110110001011;
   40754: result <= 12'b110110001011;
   40755: result <= 12'b110110001011;
   40756: result <= 12'b110110001011;
   40757: result <= 12'b110110001011;
   40758: result <= 12'b110110001011;
   40759: result <= 12'b110110001011;
   40760: result <= 12'b110110001100;
   40761: result <= 12'b110110001100;
   40762: result <= 12'b110110001100;
   40763: result <= 12'b110110001100;
   40764: result <= 12'b110110001100;
   40765: result <= 12'b110110001100;
   40766: result <= 12'b110110001100;
   40767: result <= 12'b110110001101;
   40768: result <= 12'b110110001101;
   40769: result <= 12'b110110001101;
   40770: result <= 12'b110110001101;
   40771: result <= 12'b110110001101;
   40772: result <= 12'b110110001101;
   40773: result <= 12'b110110001101;
   40774: result <= 12'b110110001110;
   40775: result <= 12'b110110001110;
   40776: result <= 12'b110110001110;
   40777: result <= 12'b110110001110;
   40778: result <= 12'b110110001110;
   40779: result <= 12'b110110001110;
   40780: result <= 12'b110110001110;
   40781: result <= 12'b110110001111;
   40782: result <= 12'b110110001111;
   40783: result <= 12'b110110001111;
   40784: result <= 12'b110110001111;
   40785: result <= 12'b110110001111;
   40786: result <= 12'b110110001111;
   40787: result <= 12'b110110001111;
   40788: result <= 12'b110110010000;
   40789: result <= 12'b110110010000;
   40790: result <= 12'b110110010000;
   40791: result <= 12'b110110010000;
   40792: result <= 12'b110110010000;
   40793: result <= 12'b110110010000;
   40794: result <= 12'b110110010000;
   40795: result <= 12'b110110010001;
   40796: result <= 12'b110110010001;
   40797: result <= 12'b110110010001;
   40798: result <= 12'b110110010001;
   40799: result <= 12'b110110010001;
   40800: result <= 12'b110110010001;
   40801: result <= 12'b110110010001;
   40802: result <= 12'b110110010010;
   40803: result <= 12'b110110010010;
   40804: result <= 12'b110110010010;
   40805: result <= 12'b110110010010;
   40806: result <= 12'b110110010010;
   40807: result <= 12'b110110010010;
   40808: result <= 12'b110110010010;
   40809: result <= 12'b110110010011;
   40810: result <= 12'b110110010011;
   40811: result <= 12'b110110010011;
   40812: result <= 12'b110110010011;
   40813: result <= 12'b110110010011;
   40814: result <= 12'b110110010011;
   40815: result <= 12'b110110010011;
   40816: result <= 12'b110110010100;
   40817: result <= 12'b110110010100;
   40818: result <= 12'b110110010100;
   40819: result <= 12'b110110010100;
   40820: result <= 12'b110110010100;
   40821: result <= 12'b110110010100;
   40822: result <= 12'b110110010100;
   40823: result <= 12'b110110010101;
   40824: result <= 12'b110110010101;
   40825: result <= 12'b110110010101;
   40826: result <= 12'b110110010101;
   40827: result <= 12'b110110010101;
   40828: result <= 12'b110110010101;
   40829: result <= 12'b110110010101;
   40830: result <= 12'b110110010101;
   40831: result <= 12'b110110010110;
   40832: result <= 12'b110110010110;
   40833: result <= 12'b110110010110;
   40834: result <= 12'b110110010110;
   40835: result <= 12'b110110010110;
   40836: result <= 12'b110110010110;
   40837: result <= 12'b110110010110;
   40838: result <= 12'b110110010111;
   40839: result <= 12'b110110010111;
   40840: result <= 12'b110110010111;
   40841: result <= 12'b110110010111;
   40842: result <= 12'b110110010111;
   40843: result <= 12'b110110010111;
   40844: result <= 12'b110110010111;
   40845: result <= 12'b110110011000;
   40846: result <= 12'b110110011000;
   40847: result <= 12'b110110011000;
   40848: result <= 12'b110110011000;
   40849: result <= 12'b110110011000;
   40850: result <= 12'b110110011000;
   40851: result <= 12'b110110011000;
   40852: result <= 12'b110110011001;
   40853: result <= 12'b110110011001;
   40854: result <= 12'b110110011001;
   40855: result <= 12'b110110011001;
   40856: result <= 12'b110110011001;
   40857: result <= 12'b110110011001;
   40858: result <= 12'b110110011001;
   40859: result <= 12'b110110011010;
   40860: result <= 12'b110110011010;
   40861: result <= 12'b110110011010;
   40862: result <= 12'b110110011010;
   40863: result <= 12'b110110011010;
   40864: result <= 12'b110110011010;
   40865: result <= 12'b110110011010;
   40866: result <= 12'b110110011011;
   40867: result <= 12'b110110011011;
   40868: result <= 12'b110110011011;
   40869: result <= 12'b110110011011;
   40870: result <= 12'b110110011011;
   40871: result <= 12'b110110011011;
   40872: result <= 12'b110110011011;
   40873: result <= 12'b110110011100;
   40874: result <= 12'b110110011100;
   40875: result <= 12'b110110011100;
   40876: result <= 12'b110110011100;
   40877: result <= 12'b110110011100;
   40878: result <= 12'b110110011100;
   40879: result <= 12'b110110011100;
   40880: result <= 12'b110110011101;
   40881: result <= 12'b110110011101;
   40882: result <= 12'b110110011101;
   40883: result <= 12'b110110011101;
   40884: result <= 12'b110110011101;
   40885: result <= 12'b110110011101;
   40886: result <= 12'b110110011101;
   40887: result <= 12'b110110011101;
   40888: result <= 12'b110110011110;
   40889: result <= 12'b110110011110;
   40890: result <= 12'b110110011110;
   40891: result <= 12'b110110011110;
   40892: result <= 12'b110110011110;
   40893: result <= 12'b110110011110;
   40894: result <= 12'b110110011110;
   40895: result <= 12'b110110011111;
   40896: result <= 12'b110110011111;
   40897: result <= 12'b110110011111;
   40898: result <= 12'b110110011111;
   40899: result <= 12'b110110011111;
   40900: result <= 12'b110110011111;
   40901: result <= 12'b110110011111;
   40902: result <= 12'b110110100000;
   40903: result <= 12'b110110100000;
   40904: result <= 12'b110110100000;
   40905: result <= 12'b110110100000;
   40906: result <= 12'b110110100000;
   40907: result <= 12'b110110100000;
   40908: result <= 12'b110110100000;
   40909: result <= 12'b110110100001;
   40910: result <= 12'b110110100001;
   40911: result <= 12'b110110100001;
   40912: result <= 12'b110110100001;
   40913: result <= 12'b110110100001;
   40914: result <= 12'b110110100001;
   40915: result <= 12'b110110100001;
   40916: result <= 12'b110110100010;
   40917: result <= 12'b110110100010;
   40918: result <= 12'b110110100010;
   40919: result <= 12'b110110100010;
   40920: result <= 12'b110110100010;
   40921: result <= 12'b110110100010;
   40922: result <= 12'b110110100010;
   40923: result <= 12'b110110100011;
   40924: result <= 12'b110110100011;
   40925: result <= 12'b110110100011;
   40926: result <= 12'b110110100011;
   40927: result <= 12'b110110100011;
   40928: result <= 12'b110110100011;
   40929: result <= 12'b110110100011;
   40930: result <= 12'b110110100011;
   40931: result <= 12'b110110100100;
   40932: result <= 12'b110110100100;
   40933: result <= 12'b110110100100;
   40934: result <= 12'b110110100100;
   40935: result <= 12'b110110100100;
   40936: result <= 12'b110110100100;
   40937: result <= 12'b110110100100;
   40938: result <= 12'b110110100101;
   40939: result <= 12'b110110100101;
   40940: result <= 12'b110110100101;
   40941: result <= 12'b110110100101;
   40942: result <= 12'b110110100101;
   40943: result <= 12'b110110100101;
   40944: result <= 12'b110110100101;
   40945: result <= 12'b110110100110;
   40946: result <= 12'b110110100110;
   40947: result <= 12'b110110100110;
   40948: result <= 12'b110110100110;
   40949: result <= 12'b110110100110;
   40950: result <= 12'b110110100110;
   40951: result <= 12'b110110100110;
   40952: result <= 12'b110110100111;
   40953: result <= 12'b110110100111;
   40954: result <= 12'b110110100111;
   40955: result <= 12'b110110100111;
   40956: result <= 12'b110110100111;
   40957: result <= 12'b110110100111;
   40958: result <= 12'b110110100111;
   40959: result <= 12'b110110101000;
   40960: result <= 12'b110110101000;
   40961: result <= 12'b110110101000;
   40962: result <= 12'b110110101000;
   40963: result <= 12'b110110101000;
   40964: result <= 12'b110110101000;
   40965: result <= 12'b110110101000;
   40966: result <= 12'b110110101000;
   40967: result <= 12'b110110101001;
   40968: result <= 12'b110110101001;
   40969: result <= 12'b110110101001;
   40970: result <= 12'b110110101001;
   40971: result <= 12'b110110101001;
   40972: result <= 12'b110110101001;
   40973: result <= 12'b110110101001;
   40974: result <= 12'b110110101010;
   40975: result <= 12'b110110101010;
   40976: result <= 12'b110110101010;
   40977: result <= 12'b110110101010;
   40978: result <= 12'b110110101010;
   40979: result <= 12'b110110101010;
   40980: result <= 12'b110110101010;
   40981: result <= 12'b110110101011;
   40982: result <= 12'b110110101011;
   40983: result <= 12'b110110101011;
   40984: result <= 12'b110110101011;
   40985: result <= 12'b110110101011;
   40986: result <= 12'b110110101011;
   40987: result <= 12'b110110101011;
   40988: result <= 12'b110110101100;
   40989: result <= 12'b110110101100;
   40990: result <= 12'b110110101100;
   40991: result <= 12'b110110101100;
   40992: result <= 12'b110110101100;
   40993: result <= 12'b110110101100;
   40994: result <= 12'b110110101100;
   40995: result <= 12'b110110101101;
   40996: result <= 12'b110110101101;
   40997: result <= 12'b110110101101;
   40998: result <= 12'b110110101101;
   40999: result <= 12'b110110101101;
   41000: result <= 12'b110110101101;
   41001: result <= 12'b110110101101;
   41002: result <= 12'b110110101101;
   41003: result <= 12'b110110101110;
   41004: result <= 12'b110110101110;
   41005: result <= 12'b110110101110;
   41006: result <= 12'b110110101110;
   41007: result <= 12'b110110101110;
   41008: result <= 12'b110110101110;
   41009: result <= 12'b110110101110;
   41010: result <= 12'b110110101111;
   41011: result <= 12'b110110101111;
   41012: result <= 12'b110110101111;
   41013: result <= 12'b110110101111;
   41014: result <= 12'b110110101111;
   41015: result <= 12'b110110101111;
   41016: result <= 12'b110110101111;
   41017: result <= 12'b110110110000;
   41018: result <= 12'b110110110000;
   41019: result <= 12'b110110110000;
   41020: result <= 12'b110110110000;
   41021: result <= 12'b110110110000;
   41022: result <= 12'b110110110000;
   41023: result <= 12'b110110110000;
   41024: result <= 12'b110110110001;
   41025: result <= 12'b110110110001;
   41026: result <= 12'b110110110001;
   41027: result <= 12'b110110110001;
   41028: result <= 12'b110110110001;
   41029: result <= 12'b110110110001;
   41030: result <= 12'b110110110001;
   41031: result <= 12'b110110110001;
   41032: result <= 12'b110110110010;
   41033: result <= 12'b110110110010;
   41034: result <= 12'b110110110010;
   41035: result <= 12'b110110110010;
   41036: result <= 12'b110110110010;
   41037: result <= 12'b110110110010;
   41038: result <= 12'b110110110010;
   41039: result <= 12'b110110110011;
   41040: result <= 12'b110110110011;
   41041: result <= 12'b110110110011;
   41042: result <= 12'b110110110011;
   41043: result <= 12'b110110110011;
   41044: result <= 12'b110110110011;
   41045: result <= 12'b110110110011;
   41046: result <= 12'b110110110100;
   41047: result <= 12'b110110110100;
   41048: result <= 12'b110110110100;
   41049: result <= 12'b110110110100;
   41050: result <= 12'b110110110100;
   41051: result <= 12'b110110110100;
   41052: result <= 12'b110110110100;
   41053: result <= 12'b110110110101;
   41054: result <= 12'b110110110101;
   41055: result <= 12'b110110110101;
   41056: result <= 12'b110110110101;
   41057: result <= 12'b110110110101;
   41058: result <= 12'b110110110101;
   41059: result <= 12'b110110110101;
   41060: result <= 12'b110110110101;
   41061: result <= 12'b110110110110;
   41062: result <= 12'b110110110110;
   41063: result <= 12'b110110110110;
   41064: result <= 12'b110110110110;
   41065: result <= 12'b110110110110;
   41066: result <= 12'b110110110110;
   41067: result <= 12'b110110110110;
   41068: result <= 12'b110110110111;
   41069: result <= 12'b110110110111;
   41070: result <= 12'b110110110111;
   41071: result <= 12'b110110110111;
   41072: result <= 12'b110110110111;
   41073: result <= 12'b110110110111;
   41074: result <= 12'b110110110111;
   41075: result <= 12'b110110111000;
   41076: result <= 12'b110110111000;
   41077: result <= 12'b110110111000;
   41078: result <= 12'b110110111000;
   41079: result <= 12'b110110111000;
   41080: result <= 12'b110110111000;
   41081: result <= 12'b110110111000;
   41082: result <= 12'b110110111000;
   41083: result <= 12'b110110111001;
   41084: result <= 12'b110110111001;
   41085: result <= 12'b110110111001;
   41086: result <= 12'b110110111001;
   41087: result <= 12'b110110111001;
   41088: result <= 12'b110110111001;
   41089: result <= 12'b110110111001;
   41090: result <= 12'b110110111010;
   41091: result <= 12'b110110111010;
   41092: result <= 12'b110110111010;
   41093: result <= 12'b110110111010;
   41094: result <= 12'b110110111010;
   41095: result <= 12'b110110111010;
   41096: result <= 12'b110110111010;
   41097: result <= 12'b110110111011;
   41098: result <= 12'b110110111011;
   41099: result <= 12'b110110111011;
   41100: result <= 12'b110110111011;
   41101: result <= 12'b110110111011;
   41102: result <= 12'b110110111011;
   41103: result <= 12'b110110111011;
   41104: result <= 12'b110110111100;
   41105: result <= 12'b110110111100;
   41106: result <= 12'b110110111100;
   41107: result <= 12'b110110111100;
   41108: result <= 12'b110110111100;
   41109: result <= 12'b110110111100;
   41110: result <= 12'b110110111100;
   41111: result <= 12'b110110111100;
   41112: result <= 12'b110110111101;
   41113: result <= 12'b110110111101;
   41114: result <= 12'b110110111101;
   41115: result <= 12'b110110111101;
   41116: result <= 12'b110110111101;
   41117: result <= 12'b110110111101;
   41118: result <= 12'b110110111101;
   41119: result <= 12'b110110111110;
   41120: result <= 12'b110110111110;
   41121: result <= 12'b110110111110;
   41122: result <= 12'b110110111110;
   41123: result <= 12'b110110111110;
   41124: result <= 12'b110110111110;
   41125: result <= 12'b110110111110;
   41126: result <= 12'b110110111111;
   41127: result <= 12'b110110111111;
   41128: result <= 12'b110110111111;
   41129: result <= 12'b110110111111;
   41130: result <= 12'b110110111111;
   41131: result <= 12'b110110111111;
   41132: result <= 12'b110110111111;
   41133: result <= 12'b110110111111;
   41134: result <= 12'b110111000000;
   41135: result <= 12'b110111000000;
   41136: result <= 12'b110111000000;
   41137: result <= 12'b110111000000;
   41138: result <= 12'b110111000000;
   41139: result <= 12'b110111000000;
   41140: result <= 12'b110111000000;
   41141: result <= 12'b110111000001;
   41142: result <= 12'b110111000001;
   41143: result <= 12'b110111000001;
   41144: result <= 12'b110111000001;
   41145: result <= 12'b110111000001;
   41146: result <= 12'b110111000001;
   41147: result <= 12'b110111000001;
   41148: result <= 12'b110111000010;
   41149: result <= 12'b110111000010;
   41150: result <= 12'b110111000010;
   41151: result <= 12'b110111000010;
   41152: result <= 12'b110111000010;
   41153: result <= 12'b110111000010;
   41154: result <= 12'b110111000010;
   41155: result <= 12'b110111000010;
   41156: result <= 12'b110111000011;
   41157: result <= 12'b110111000011;
   41158: result <= 12'b110111000011;
   41159: result <= 12'b110111000011;
   41160: result <= 12'b110111000011;
   41161: result <= 12'b110111000011;
   41162: result <= 12'b110111000011;
   41163: result <= 12'b110111000100;
   41164: result <= 12'b110111000100;
   41165: result <= 12'b110111000100;
   41166: result <= 12'b110111000100;
   41167: result <= 12'b110111000100;
   41168: result <= 12'b110111000100;
   41169: result <= 12'b110111000100;
   41170: result <= 12'b110111000101;
   41171: result <= 12'b110111000101;
   41172: result <= 12'b110111000101;
   41173: result <= 12'b110111000101;
   41174: result <= 12'b110111000101;
   41175: result <= 12'b110111000101;
   41176: result <= 12'b110111000101;
   41177: result <= 12'b110111000101;
   41178: result <= 12'b110111000110;
   41179: result <= 12'b110111000110;
   41180: result <= 12'b110111000110;
   41181: result <= 12'b110111000110;
   41182: result <= 12'b110111000110;
   41183: result <= 12'b110111000110;
   41184: result <= 12'b110111000110;
   41185: result <= 12'b110111000111;
   41186: result <= 12'b110111000111;
   41187: result <= 12'b110111000111;
   41188: result <= 12'b110111000111;
   41189: result <= 12'b110111000111;
   41190: result <= 12'b110111000111;
   41191: result <= 12'b110111000111;
   41192: result <= 12'b110111001000;
   41193: result <= 12'b110111001000;
   41194: result <= 12'b110111001000;
   41195: result <= 12'b110111001000;
   41196: result <= 12'b110111001000;
   41197: result <= 12'b110111001000;
   41198: result <= 12'b110111001000;
   41199: result <= 12'b110111001000;
   41200: result <= 12'b110111001001;
   41201: result <= 12'b110111001001;
   41202: result <= 12'b110111001001;
   41203: result <= 12'b110111001001;
   41204: result <= 12'b110111001001;
   41205: result <= 12'b110111001001;
   41206: result <= 12'b110111001001;
   41207: result <= 12'b110111001010;
   41208: result <= 12'b110111001010;
   41209: result <= 12'b110111001010;
   41210: result <= 12'b110111001010;
   41211: result <= 12'b110111001010;
   41212: result <= 12'b110111001010;
   41213: result <= 12'b110111001010;
   41214: result <= 12'b110111001010;
   41215: result <= 12'b110111001011;
   41216: result <= 12'b110111001011;
   41217: result <= 12'b110111001011;
   41218: result <= 12'b110111001011;
   41219: result <= 12'b110111001011;
   41220: result <= 12'b110111001011;
   41221: result <= 12'b110111001011;
   41222: result <= 12'b110111001100;
   41223: result <= 12'b110111001100;
   41224: result <= 12'b110111001100;
   41225: result <= 12'b110111001100;
   41226: result <= 12'b110111001100;
   41227: result <= 12'b110111001100;
   41228: result <= 12'b110111001100;
   41229: result <= 12'b110111001101;
   41230: result <= 12'b110111001101;
   41231: result <= 12'b110111001101;
   41232: result <= 12'b110111001101;
   41233: result <= 12'b110111001101;
   41234: result <= 12'b110111001101;
   41235: result <= 12'b110111001101;
   41236: result <= 12'b110111001101;
   41237: result <= 12'b110111001110;
   41238: result <= 12'b110111001110;
   41239: result <= 12'b110111001110;
   41240: result <= 12'b110111001110;
   41241: result <= 12'b110111001110;
   41242: result <= 12'b110111001110;
   41243: result <= 12'b110111001110;
   41244: result <= 12'b110111001111;
   41245: result <= 12'b110111001111;
   41246: result <= 12'b110111001111;
   41247: result <= 12'b110111001111;
   41248: result <= 12'b110111001111;
   41249: result <= 12'b110111001111;
   41250: result <= 12'b110111001111;
   41251: result <= 12'b110111001111;
   41252: result <= 12'b110111010000;
   41253: result <= 12'b110111010000;
   41254: result <= 12'b110111010000;
   41255: result <= 12'b110111010000;
   41256: result <= 12'b110111010000;
   41257: result <= 12'b110111010000;
   41258: result <= 12'b110111010000;
   41259: result <= 12'b110111010001;
   41260: result <= 12'b110111010001;
   41261: result <= 12'b110111010001;
   41262: result <= 12'b110111010001;
   41263: result <= 12'b110111010001;
   41264: result <= 12'b110111010001;
   41265: result <= 12'b110111010001;
   41266: result <= 12'b110111010010;
   41267: result <= 12'b110111010010;
   41268: result <= 12'b110111010010;
   41269: result <= 12'b110111010010;
   41270: result <= 12'b110111010010;
   41271: result <= 12'b110111010010;
   41272: result <= 12'b110111010010;
   41273: result <= 12'b110111010010;
   41274: result <= 12'b110111010011;
   41275: result <= 12'b110111010011;
   41276: result <= 12'b110111010011;
   41277: result <= 12'b110111010011;
   41278: result <= 12'b110111010011;
   41279: result <= 12'b110111010011;
   41280: result <= 12'b110111010011;
   41281: result <= 12'b110111010100;
   41282: result <= 12'b110111010100;
   41283: result <= 12'b110111010100;
   41284: result <= 12'b110111010100;
   41285: result <= 12'b110111010100;
   41286: result <= 12'b110111010100;
   41287: result <= 12'b110111010100;
   41288: result <= 12'b110111010100;
   41289: result <= 12'b110111010101;
   41290: result <= 12'b110111010101;
   41291: result <= 12'b110111010101;
   41292: result <= 12'b110111010101;
   41293: result <= 12'b110111010101;
   41294: result <= 12'b110111010101;
   41295: result <= 12'b110111010101;
   41296: result <= 12'b110111010110;
   41297: result <= 12'b110111010110;
   41298: result <= 12'b110111010110;
   41299: result <= 12'b110111010110;
   41300: result <= 12'b110111010110;
   41301: result <= 12'b110111010110;
   41302: result <= 12'b110111010110;
   41303: result <= 12'b110111010110;
   41304: result <= 12'b110111010111;
   41305: result <= 12'b110111010111;
   41306: result <= 12'b110111010111;
   41307: result <= 12'b110111010111;
   41308: result <= 12'b110111010111;
   41309: result <= 12'b110111010111;
   41310: result <= 12'b110111010111;
   41311: result <= 12'b110111011000;
   41312: result <= 12'b110111011000;
   41313: result <= 12'b110111011000;
   41314: result <= 12'b110111011000;
   41315: result <= 12'b110111011000;
   41316: result <= 12'b110111011000;
   41317: result <= 12'b110111011000;
   41318: result <= 12'b110111011000;
   41319: result <= 12'b110111011001;
   41320: result <= 12'b110111011001;
   41321: result <= 12'b110111011001;
   41322: result <= 12'b110111011001;
   41323: result <= 12'b110111011001;
   41324: result <= 12'b110111011001;
   41325: result <= 12'b110111011001;
   41326: result <= 12'b110111011010;
   41327: result <= 12'b110111011010;
   41328: result <= 12'b110111011010;
   41329: result <= 12'b110111011010;
   41330: result <= 12'b110111011010;
   41331: result <= 12'b110111011010;
   41332: result <= 12'b110111011010;
   41333: result <= 12'b110111011011;
   41334: result <= 12'b110111011011;
   41335: result <= 12'b110111011011;
   41336: result <= 12'b110111011011;
   41337: result <= 12'b110111011011;
   41338: result <= 12'b110111011011;
   41339: result <= 12'b110111011011;
   41340: result <= 12'b110111011011;
   41341: result <= 12'b110111011100;
   41342: result <= 12'b110111011100;
   41343: result <= 12'b110111011100;
   41344: result <= 12'b110111011100;
   41345: result <= 12'b110111011100;
   41346: result <= 12'b110111011100;
   41347: result <= 12'b110111011100;
   41348: result <= 12'b110111011101;
   41349: result <= 12'b110111011101;
   41350: result <= 12'b110111011101;
   41351: result <= 12'b110111011101;
   41352: result <= 12'b110111011101;
   41353: result <= 12'b110111011101;
   41354: result <= 12'b110111011101;
   41355: result <= 12'b110111011101;
   41356: result <= 12'b110111011110;
   41357: result <= 12'b110111011110;
   41358: result <= 12'b110111011110;
   41359: result <= 12'b110111011110;
   41360: result <= 12'b110111011110;
   41361: result <= 12'b110111011110;
   41362: result <= 12'b110111011110;
   41363: result <= 12'b110111011111;
   41364: result <= 12'b110111011111;
   41365: result <= 12'b110111011111;
   41366: result <= 12'b110111011111;
   41367: result <= 12'b110111011111;
   41368: result <= 12'b110111011111;
   41369: result <= 12'b110111011111;
   41370: result <= 12'b110111011111;
   41371: result <= 12'b110111100000;
   41372: result <= 12'b110111100000;
   41373: result <= 12'b110111100000;
   41374: result <= 12'b110111100000;
   41375: result <= 12'b110111100000;
   41376: result <= 12'b110111100000;
   41377: result <= 12'b110111100000;
   41378: result <= 12'b110111100001;
   41379: result <= 12'b110111100001;
   41380: result <= 12'b110111100001;
   41381: result <= 12'b110111100001;
   41382: result <= 12'b110111100001;
   41383: result <= 12'b110111100001;
   41384: result <= 12'b110111100001;
   41385: result <= 12'b110111100001;
   41386: result <= 12'b110111100010;
   41387: result <= 12'b110111100010;
   41388: result <= 12'b110111100010;
   41389: result <= 12'b110111100010;
   41390: result <= 12'b110111100010;
   41391: result <= 12'b110111100010;
   41392: result <= 12'b110111100010;
   41393: result <= 12'b110111100011;
   41394: result <= 12'b110111100011;
   41395: result <= 12'b110111100011;
   41396: result <= 12'b110111100011;
   41397: result <= 12'b110111100011;
   41398: result <= 12'b110111100011;
   41399: result <= 12'b110111100011;
   41400: result <= 12'b110111100011;
   41401: result <= 12'b110111100100;
   41402: result <= 12'b110111100100;
   41403: result <= 12'b110111100100;
   41404: result <= 12'b110111100100;
   41405: result <= 12'b110111100100;
   41406: result <= 12'b110111100100;
   41407: result <= 12'b110111100100;
   41408: result <= 12'b110111100101;
   41409: result <= 12'b110111100101;
   41410: result <= 12'b110111100101;
   41411: result <= 12'b110111100101;
   41412: result <= 12'b110111100101;
   41413: result <= 12'b110111100101;
   41414: result <= 12'b110111100101;
   41415: result <= 12'b110111100101;
   41416: result <= 12'b110111100110;
   41417: result <= 12'b110111100110;
   41418: result <= 12'b110111100110;
   41419: result <= 12'b110111100110;
   41420: result <= 12'b110111100110;
   41421: result <= 12'b110111100110;
   41422: result <= 12'b110111100110;
   41423: result <= 12'b110111100110;
   41424: result <= 12'b110111100111;
   41425: result <= 12'b110111100111;
   41426: result <= 12'b110111100111;
   41427: result <= 12'b110111100111;
   41428: result <= 12'b110111100111;
   41429: result <= 12'b110111100111;
   41430: result <= 12'b110111100111;
   41431: result <= 12'b110111101000;
   41432: result <= 12'b110111101000;
   41433: result <= 12'b110111101000;
   41434: result <= 12'b110111101000;
   41435: result <= 12'b110111101000;
   41436: result <= 12'b110111101000;
   41437: result <= 12'b110111101000;
   41438: result <= 12'b110111101000;
   41439: result <= 12'b110111101001;
   41440: result <= 12'b110111101001;
   41441: result <= 12'b110111101001;
   41442: result <= 12'b110111101001;
   41443: result <= 12'b110111101001;
   41444: result <= 12'b110111101001;
   41445: result <= 12'b110111101001;
   41446: result <= 12'b110111101010;
   41447: result <= 12'b110111101010;
   41448: result <= 12'b110111101010;
   41449: result <= 12'b110111101010;
   41450: result <= 12'b110111101010;
   41451: result <= 12'b110111101010;
   41452: result <= 12'b110111101010;
   41453: result <= 12'b110111101010;
   41454: result <= 12'b110111101011;
   41455: result <= 12'b110111101011;
   41456: result <= 12'b110111101011;
   41457: result <= 12'b110111101011;
   41458: result <= 12'b110111101011;
   41459: result <= 12'b110111101011;
   41460: result <= 12'b110111101011;
   41461: result <= 12'b110111101100;
   41462: result <= 12'b110111101100;
   41463: result <= 12'b110111101100;
   41464: result <= 12'b110111101100;
   41465: result <= 12'b110111101100;
   41466: result <= 12'b110111101100;
   41467: result <= 12'b110111101100;
   41468: result <= 12'b110111101100;
   41469: result <= 12'b110111101101;
   41470: result <= 12'b110111101101;
   41471: result <= 12'b110111101101;
   41472: result <= 12'b110111101101;
   41473: result <= 12'b110111101101;
   41474: result <= 12'b110111101101;
   41475: result <= 12'b110111101101;
   41476: result <= 12'b110111101101;
   41477: result <= 12'b110111101110;
   41478: result <= 12'b110111101110;
   41479: result <= 12'b110111101110;
   41480: result <= 12'b110111101110;
   41481: result <= 12'b110111101110;
   41482: result <= 12'b110111101110;
   41483: result <= 12'b110111101110;
   41484: result <= 12'b110111101111;
   41485: result <= 12'b110111101111;
   41486: result <= 12'b110111101111;
   41487: result <= 12'b110111101111;
   41488: result <= 12'b110111101111;
   41489: result <= 12'b110111101111;
   41490: result <= 12'b110111101111;
   41491: result <= 12'b110111101111;
   41492: result <= 12'b110111110000;
   41493: result <= 12'b110111110000;
   41494: result <= 12'b110111110000;
   41495: result <= 12'b110111110000;
   41496: result <= 12'b110111110000;
   41497: result <= 12'b110111110000;
   41498: result <= 12'b110111110000;
   41499: result <= 12'b110111110001;
   41500: result <= 12'b110111110001;
   41501: result <= 12'b110111110001;
   41502: result <= 12'b110111110001;
   41503: result <= 12'b110111110001;
   41504: result <= 12'b110111110001;
   41505: result <= 12'b110111110001;
   41506: result <= 12'b110111110001;
   41507: result <= 12'b110111110010;
   41508: result <= 12'b110111110010;
   41509: result <= 12'b110111110010;
   41510: result <= 12'b110111110010;
   41511: result <= 12'b110111110010;
   41512: result <= 12'b110111110010;
   41513: result <= 12'b110111110010;
   41514: result <= 12'b110111110010;
   41515: result <= 12'b110111110011;
   41516: result <= 12'b110111110011;
   41517: result <= 12'b110111110011;
   41518: result <= 12'b110111110011;
   41519: result <= 12'b110111110011;
   41520: result <= 12'b110111110011;
   41521: result <= 12'b110111110011;
   41522: result <= 12'b110111110100;
   41523: result <= 12'b110111110100;
   41524: result <= 12'b110111110100;
   41525: result <= 12'b110111110100;
   41526: result <= 12'b110111110100;
   41527: result <= 12'b110111110100;
   41528: result <= 12'b110111110100;
   41529: result <= 12'b110111110100;
   41530: result <= 12'b110111110101;
   41531: result <= 12'b110111110101;
   41532: result <= 12'b110111110101;
   41533: result <= 12'b110111110101;
   41534: result <= 12'b110111110101;
   41535: result <= 12'b110111110101;
   41536: result <= 12'b110111110101;
   41537: result <= 12'b110111110110;
   41538: result <= 12'b110111110110;
   41539: result <= 12'b110111110110;
   41540: result <= 12'b110111110110;
   41541: result <= 12'b110111110110;
   41542: result <= 12'b110111110110;
   41543: result <= 12'b110111110110;
   41544: result <= 12'b110111110110;
   41545: result <= 12'b110111110111;
   41546: result <= 12'b110111110111;
   41547: result <= 12'b110111110111;
   41548: result <= 12'b110111110111;
   41549: result <= 12'b110111110111;
   41550: result <= 12'b110111110111;
   41551: result <= 12'b110111110111;
   41552: result <= 12'b110111110111;
   41553: result <= 12'b110111111000;
   41554: result <= 12'b110111111000;
   41555: result <= 12'b110111111000;
   41556: result <= 12'b110111111000;
   41557: result <= 12'b110111111000;
   41558: result <= 12'b110111111000;
   41559: result <= 12'b110111111000;
   41560: result <= 12'b110111111001;
   41561: result <= 12'b110111111001;
   41562: result <= 12'b110111111001;
   41563: result <= 12'b110111111001;
   41564: result <= 12'b110111111001;
   41565: result <= 12'b110111111001;
   41566: result <= 12'b110111111001;
   41567: result <= 12'b110111111001;
   41568: result <= 12'b110111111010;
   41569: result <= 12'b110111111010;
   41570: result <= 12'b110111111010;
   41571: result <= 12'b110111111010;
   41572: result <= 12'b110111111010;
   41573: result <= 12'b110111111010;
   41574: result <= 12'b110111111010;
   41575: result <= 12'b110111111010;
   41576: result <= 12'b110111111011;
   41577: result <= 12'b110111111011;
   41578: result <= 12'b110111111011;
   41579: result <= 12'b110111111011;
   41580: result <= 12'b110111111011;
   41581: result <= 12'b110111111011;
   41582: result <= 12'b110111111011;
   41583: result <= 12'b110111111100;
   41584: result <= 12'b110111111100;
   41585: result <= 12'b110111111100;
   41586: result <= 12'b110111111100;
   41587: result <= 12'b110111111100;
   41588: result <= 12'b110111111100;
   41589: result <= 12'b110111111100;
   41590: result <= 12'b110111111100;
   41591: result <= 12'b110111111101;
   41592: result <= 12'b110111111101;
   41593: result <= 12'b110111111101;
   41594: result <= 12'b110111111101;
   41595: result <= 12'b110111111101;
   41596: result <= 12'b110111111101;
   41597: result <= 12'b110111111101;
   41598: result <= 12'b110111111101;
   41599: result <= 12'b110111111110;
   41600: result <= 12'b110111111110;
   41601: result <= 12'b110111111110;
   41602: result <= 12'b110111111110;
   41603: result <= 12'b110111111110;
   41604: result <= 12'b110111111110;
   41605: result <= 12'b110111111110;
   41606: result <= 12'b110111111111;
   41607: result <= 12'b110111111111;
   41608: result <= 12'b110111111111;
   41609: result <= 12'b110111111111;
   41610: result <= 12'b110111111111;
   41611: result <= 12'b110111111111;
   41612: result <= 12'b110111111111;
   41613: result <= 12'b110111111111;
   41614: result <= 12'b111000000000;
   41615: result <= 12'b111000000000;
   41616: result <= 12'b111000000000;
   41617: result <= 12'b111000000000;
   41618: result <= 12'b111000000000;
   41619: result <= 12'b111000000000;
   41620: result <= 12'b111000000000;
   41621: result <= 12'b111000000000;
   41622: result <= 12'b111000000001;
   41623: result <= 12'b111000000001;
   41624: result <= 12'b111000000001;
   41625: result <= 12'b111000000001;
   41626: result <= 12'b111000000001;
   41627: result <= 12'b111000000001;
   41628: result <= 12'b111000000001;
   41629: result <= 12'b111000000001;
   41630: result <= 12'b111000000010;
   41631: result <= 12'b111000000010;
   41632: result <= 12'b111000000010;
   41633: result <= 12'b111000000010;
   41634: result <= 12'b111000000010;
   41635: result <= 12'b111000000010;
   41636: result <= 12'b111000000010;
   41637: result <= 12'b111000000011;
   41638: result <= 12'b111000000011;
   41639: result <= 12'b111000000011;
   41640: result <= 12'b111000000011;
   41641: result <= 12'b111000000011;
   41642: result <= 12'b111000000011;
   41643: result <= 12'b111000000011;
   41644: result <= 12'b111000000011;
   41645: result <= 12'b111000000100;
   41646: result <= 12'b111000000100;
   41647: result <= 12'b111000000100;
   41648: result <= 12'b111000000100;
   41649: result <= 12'b111000000100;
   41650: result <= 12'b111000000100;
   41651: result <= 12'b111000000100;
   41652: result <= 12'b111000000100;
   41653: result <= 12'b111000000101;
   41654: result <= 12'b111000000101;
   41655: result <= 12'b111000000101;
   41656: result <= 12'b111000000101;
   41657: result <= 12'b111000000101;
   41658: result <= 12'b111000000101;
   41659: result <= 12'b111000000101;
   41660: result <= 12'b111000000110;
   41661: result <= 12'b111000000110;
   41662: result <= 12'b111000000110;
   41663: result <= 12'b111000000110;
   41664: result <= 12'b111000000110;
   41665: result <= 12'b111000000110;
   41666: result <= 12'b111000000110;
   41667: result <= 12'b111000000110;
   41668: result <= 12'b111000000111;
   41669: result <= 12'b111000000111;
   41670: result <= 12'b111000000111;
   41671: result <= 12'b111000000111;
   41672: result <= 12'b111000000111;
   41673: result <= 12'b111000000111;
   41674: result <= 12'b111000000111;
   41675: result <= 12'b111000000111;
   41676: result <= 12'b111000001000;
   41677: result <= 12'b111000001000;
   41678: result <= 12'b111000001000;
   41679: result <= 12'b111000001000;
   41680: result <= 12'b111000001000;
   41681: result <= 12'b111000001000;
   41682: result <= 12'b111000001000;
   41683: result <= 12'b111000001000;
   41684: result <= 12'b111000001001;
   41685: result <= 12'b111000001001;
   41686: result <= 12'b111000001001;
   41687: result <= 12'b111000001001;
   41688: result <= 12'b111000001001;
   41689: result <= 12'b111000001001;
   41690: result <= 12'b111000001001;
   41691: result <= 12'b111000001010;
   41692: result <= 12'b111000001010;
   41693: result <= 12'b111000001010;
   41694: result <= 12'b111000001010;
   41695: result <= 12'b111000001010;
   41696: result <= 12'b111000001010;
   41697: result <= 12'b111000001010;
   41698: result <= 12'b111000001010;
   41699: result <= 12'b111000001011;
   41700: result <= 12'b111000001011;
   41701: result <= 12'b111000001011;
   41702: result <= 12'b111000001011;
   41703: result <= 12'b111000001011;
   41704: result <= 12'b111000001011;
   41705: result <= 12'b111000001011;
   41706: result <= 12'b111000001011;
   41707: result <= 12'b111000001100;
   41708: result <= 12'b111000001100;
   41709: result <= 12'b111000001100;
   41710: result <= 12'b111000001100;
   41711: result <= 12'b111000001100;
   41712: result <= 12'b111000001100;
   41713: result <= 12'b111000001100;
   41714: result <= 12'b111000001100;
   41715: result <= 12'b111000001101;
   41716: result <= 12'b111000001101;
   41717: result <= 12'b111000001101;
   41718: result <= 12'b111000001101;
   41719: result <= 12'b111000001101;
   41720: result <= 12'b111000001101;
   41721: result <= 12'b111000001101;
   41722: result <= 12'b111000001101;
   41723: result <= 12'b111000001110;
   41724: result <= 12'b111000001110;
   41725: result <= 12'b111000001110;
   41726: result <= 12'b111000001110;
   41727: result <= 12'b111000001110;
   41728: result <= 12'b111000001110;
   41729: result <= 12'b111000001110;
   41730: result <= 12'b111000001111;
   41731: result <= 12'b111000001111;
   41732: result <= 12'b111000001111;
   41733: result <= 12'b111000001111;
   41734: result <= 12'b111000001111;
   41735: result <= 12'b111000001111;
   41736: result <= 12'b111000001111;
   41737: result <= 12'b111000001111;
   41738: result <= 12'b111000010000;
   41739: result <= 12'b111000010000;
   41740: result <= 12'b111000010000;
   41741: result <= 12'b111000010000;
   41742: result <= 12'b111000010000;
   41743: result <= 12'b111000010000;
   41744: result <= 12'b111000010000;
   41745: result <= 12'b111000010000;
   41746: result <= 12'b111000010001;
   41747: result <= 12'b111000010001;
   41748: result <= 12'b111000010001;
   41749: result <= 12'b111000010001;
   41750: result <= 12'b111000010001;
   41751: result <= 12'b111000010001;
   41752: result <= 12'b111000010001;
   41753: result <= 12'b111000010001;
   41754: result <= 12'b111000010010;
   41755: result <= 12'b111000010010;
   41756: result <= 12'b111000010010;
   41757: result <= 12'b111000010010;
   41758: result <= 12'b111000010010;
   41759: result <= 12'b111000010010;
   41760: result <= 12'b111000010010;
   41761: result <= 12'b111000010010;
   41762: result <= 12'b111000010011;
   41763: result <= 12'b111000010011;
   41764: result <= 12'b111000010011;
   41765: result <= 12'b111000010011;
   41766: result <= 12'b111000010011;
   41767: result <= 12'b111000010011;
   41768: result <= 12'b111000010011;
   41769: result <= 12'b111000010100;
   41770: result <= 12'b111000010100;
   41771: result <= 12'b111000010100;
   41772: result <= 12'b111000010100;
   41773: result <= 12'b111000010100;
   41774: result <= 12'b111000010100;
   41775: result <= 12'b111000010100;
   41776: result <= 12'b111000010100;
   41777: result <= 12'b111000010101;
   41778: result <= 12'b111000010101;
   41779: result <= 12'b111000010101;
   41780: result <= 12'b111000010101;
   41781: result <= 12'b111000010101;
   41782: result <= 12'b111000010101;
   41783: result <= 12'b111000010101;
   41784: result <= 12'b111000010101;
   41785: result <= 12'b111000010110;
   41786: result <= 12'b111000010110;
   41787: result <= 12'b111000010110;
   41788: result <= 12'b111000010110;
   41789: result <= 12'b111000010110;
   41790: result <= 12'b111000010110;
   41791: result <= 12'b111000010110;
   41792: result <= 12'b111000010110;
   41793: result <= 12'b111000010111;
   41794: result <= 12'b111000010111;
   41795: result <= 12'b111000010111;
   41796: result <= 12'b111000010111;
   41797: result <= 12'b111000010111;
   41798: result <= 12'b111000010111;
   41799: result <= 12'b111000010111;
   41800: result <= 12'b111000010111;
   41801: result <= 12'b111000011000;
   41802: result <= 12'b111000011000;
   41803: result <= 12'b111000011000;
   41804: result <= 12'b111000011000;
   41805: result <= 12'b111000011000;
   41806: result <= 12'b111000011000;
   41807: result <= 12'b111000011000;
   41808: result <= 12'b111000011000;
   41809: result <= 12'b111000011001;
   41810: result <= 12'b111000011001;
   41811: result <= 12'b111000011001;
   41812: result <= 12'b111000011001;
   41813: result <= 12'b111000011001;
   41814: result <= 12'b111000011001;
   41815: result <= 12'b111000011001;
   41816: result <= 12'b111000011001;
   41817: result <= 12'b111000011010;
   41818: result <= 12'b111000011010;
   41819: result <= 12'b111000011010;
   41820: result <= 12'b111000011010;
   41821: result <= 12'b111000011010;
   41822: result <= 12'b111000011010;
   41823: result <= 12'b111000011010;
   41824: result <= 12'b111000011011;
   41825: result <= 12'b111000011011;
   41826: result <= 12'b111000011011;
   41827: result <= 12'b111000011011;
   41828: result <= 12'b111000011011;
   41829: result <= 12'b111000011011;
   41830: result <= 12'b111000011011;
   41831: result <= 12'b111000011011;
   41832: result <= 12'b111000011100;
   41833: result <= 12'b111000011100;
   41834: result <= 12'b111000011100;
   41835: result <= 12'b111000011100;
   41836: result <= 12'b111000011100;
   41837: result <= 12'b111000011100;
   41838: result <= 12'b111000011100;
   41839: result <= 12'b111000011100;
   41840: result <= 12'b111000011101;
   41841: result <= 12'b111000011101;
   41842: result <= 12'b111000011101;
   41843: result <= 12'b111000011101;
   41844: result <= 12'b111000011101;
   41845: result <= 12'b111000011101;
   41846: result <= 12'b111000011101;
   41847: result <= 12'b111000011101;
   41848: result <= 12'b111000011110;
   41849: result <= 12'b111000011110;
   41850: result <= 12'b111000011110;
   41851: result <= 12'b111000011110;
   41852: result <= 12'b111000011110;
   41853: result <= 12'b111000011110;
   41854: result <= 12'b111000011110;
   41855: result <= 12'b111000011110;
   41856: result <= 12'b111000011111;
   41857: result <= 12'b111000011111;
   41858: result <= 12'b111000011111;
   41859: result <= 12'b111000011111;
   41860: result <= 12'b111000011111;
   41861: result <= 12'b111000011111;
   41862: result <= 12'b111000011111;
   41863: result <= 12'b111000011111;
   41864: result <= 12'b111000100000;
   41865: result <= 12'b111000100000;
   41866: result <= 12'b111000100000;
   41867: result <= 12'b111000100000;
   41868: result <= 12'b111000100000;
   41869: result <= 12'b111000100000;
   41870: result <= 12'b111000100000;
   41871: result <= 12'b111000100000;
   41872: result <= 12'b111000100001;
   41873: result <= 12'b111000100001;
   41874: result <= 12'b111000100001;
   41875: result <= 12'b111000100001;
   41876: result <= 12'b111000100001;
   41877: result <= 12'b111000100001;
   41878: result <= 12'b111000100001;
   41879: result <= 12'b111000100001;
   41880: result <= 12'b111000100010;
   41881: result <= 12'b111000100010;
   41882: result <= 12'b111000100010;
   41883: result <= 12'b111000100010;
   41884: result <= 12'b111000100010;
   41885: result <= 12'b111000100010;
   41886: result <= 12'b111000100010;
   41887: result <= 12'b111000100010;
   41888: result <= 12'b111000100011;
   41889: result <= 12'b111000100011;
   41890: result <= 12'b111000100011;
   41891: result <= 12'b111000100011;
   41892: result <= 12'b111000100011;
   41893: result <= 12'b111000100011;
   41894: result <= 12'b111000100011;
   41895: result <= 12'b111000100011;
   41896: result <= 12'b111000100100;
   41897: result <= 12'b111000100100;
   41898: result <= 12'b111000100100;
   41899: result <= 12'b111000100100;
   41900: result <= 12'b111000100100;
   41901: result <= 12'b111000100100;
   41902: result <= 12'b111000100100;
   41903: result <= 12'b111000100100;
   41904: result <= 12'b111000100101;
   41905: result <= 12'b111000100101;
   41906: result <= 12'b111000100101;
   41907: result <= 12'b111000100101;
   41908: result <= 12'b111000100101;
   41909: result <= 12'b111000100101;
   41910: result <= 12'b111000100101;
   41911: result <= 12'b111000100101;
   41912: result <= 12'b111000100110;
   41913: result <= 12'b111000100110;
   41914: result <= 12'b111000100110;
   41915: result <= 12'b111000100110;
   41916: result <= 12'b111000100110;
   41917: result <= 12'b111000100110;
   41918: result <= 12'b111000100110;
   41919: result <= 12'b111000100110;
   41920: result <= 12'b111000100111;
   41921: result <= 12'b111000100111;
   41922: result <= 12'b111000100111;
   41923: result <= 12'b111000100111;
   41924: result <= 12'b111000100111;
   41925: result <= 12'b111000100111;
   41926: result <= 12'b111000100111;
   41927: result <= 12'b111000101000;
   41928: result <= 12'b111000101000;
   41929: result <= 12'b111000101000;
   41930: result <= 12'b111000101000;
   41931: result <= 12'b111000101000;
   41932: result <= 12'b111000101000;
   41933: result <= 12'b111000101000;
   41934: result <= 12'b111000101000;
   41935: result <= 12'b111000101001;
   41936: result <= 12'b111000101001;
   41937: result <= 12'b111000101001;
   41938: result <= 12'b111000101001;
   41939: result <= 12'b111000101001;
   41940: result <= 12'b111000101001;
   41941: result <= 12'b111000101001;
   41942: result <= 12'b111000101001;
   41943: result <= 12'b111000101010;
   41944: result <= 12'b111000101010;
   41945: result <= 12'b111000101010;
   41946: result <= 12'b111000101010;
   41947: result <= 12'b111000101010;
   41948: result <= 12'b111000101010;
   41949: result <= 12'b111000101010;
   41950: result <= 12'b111000101010;
   41951: result <= 12'b111000101011;
   41952: result <= 12'b111000101011;
   41953: result <= 12'b111000101011;
   41954: result <= 12'b111000101011;
   41955: result <= 12'b111000101011;
   41956: result <= 12'b111000101011;
   41957: result <= 12'b111000101011;
   41958: result <= 12'b111000101011;
   41959: result <= 12'b111000101100;
   41960: result <= 12'b111000101100;
   41961: result <= 12'b111000101100;
   41962: result <= 12'b111000101100;
   41963: result <= 12'b111000101100;
   41964: result <= 12'b111000101100;
   41965: result <= 12'b111000101100;
   41966: result <= 12'b111000101100;
   41967: result <= 12'b111000101101;
   41968: result <= 12'b111000101101;
   41969: result <= 12'b111000101101;
   41970: result <= 12'b111000101101;
   41971: result <= 12'b111000101101;
   41972: result <= 12'b111000101101;
   41973: result <= 12'b111000101101;
   41974: result <= 12'b111000101101;
   41975: result <= 12'b111000101110;
   41976: result <= 12'b111000101110;
   41977: result <= 12'b111000101110;
   41978: result <= 12'b111000101110;
   41979: result <= 12'b111000101110;
   41980: result <= 12'b111000101110;
   41981: result <= 12'b111000101110;
   41982: result <= 12'b111000101110;
   41983: result <= 12'b111000101111;
   41984: result <= 12'b111000101111;
   41985: result <= 12'b111000101111;
   41986: result <= 12'b111000101111;
   41987: result <= 12'b111000101111;
   41988: result <= 12'b111000101111;
   41989: result <= 12'b111000101111;
   41990: result <= 12'b111000101111;
   41991: result <= 12'b111000101111;
   41992: result <= 12'b111000110000;
   41993: result <= 12'b111000110000;
   41994: result <= 12'b111000110000;
   41995: result <= 12'b111000110000;
   41996: result <= 12'b111000110000;
   41997: result <= 12'b111000110000;
   41998: result <= 12'b111000110000;
   41999: result <= 12'b111000110000;
   42000: result <= 12'b111000110001;
   42001: result <= 12'b111000110001;
   42002: result <= 12'b111000110001;
   42003: result <= 12'b111000110001;
   42004: result <= 12'b111000110001;
   42005: result <= 12'b111000110001;
   42006: result <= 12'b111000110001;
   42007: result <= 12'b111000110001;
   42008: result <= 12'b111000110010;
   42009: result <= 12'b111000110010;
   42010: result <= 12'b111000110010;
   42011: result <= 12'b111000110010;
   42012: result <= 12'b111000110010;
   42013: result <= 12'b111000110010;
   42014: result <= 12'b111000110010;
   42015: result <= 12'b111000110010;
   42016: result <= 12'b111000110011;
   42017: result <= 12'b111000110011;
   42018: result <= 12'b111000110011;
   42019: result <= 12'b111000110011;
   42020: result <= 12'b111000110011;
   42021: result <= 12'b111000110011;
   42022: result <= 12'b111000110011;
   42023: result <= 12'b111000110011;
   42024: result <= 12'b111000110100;
   42025: result <= 12'b111000110100;
   42026: result <= 12'b111000110100;
   42027: result <= 12'b111000110100;
   42028: result <= 12'b111000110100;
   42029: result <= 12'b111000110100;
   42030: result <= 12'b111000110100;
   42031: result <= 12'b111000110100;
   42032: result <= 12'b111000110101;
   42033: result <= 12'b111000110101;
   42034: result <= 12'b111000110101;
   42035: result <= 12'b111000110101;
   42036: result <= 12'b111000110101;
   42037: result <= 12'b111000110101;
   42038: result <= 12'b111000110101;
   42039: result <= 12'b111000110101;
   42040: result <= 12'b111000110110;
   42041: result <= 12'b111000110110;
   42042: result <= 12'b111000110110;
   42043: result <= 12'b111000110110;
   42044: result <= 12'b111000110110;
   42045: result <= 12'b111000110110;
   42046: result <= 12'b111000110110;
   42047: result <= 12'b111000110110;
   42048: result <= 12'b111000110111;
   42049: result <= 12'b111000110111;
   42050: result <= 12'b111000110111;
   42051: result <= 12'b111000110111;
   42052: result <= 12'b111000110111;
   42053: result <= 12'b111000110111;
   42054: result <= 12'b111000110111;
   42055: result <= 12'b111000110111;
   42056: result <= 12'b111000111000;
   42057: result <= 12'b111000111000;
   42058: result <= 12'b111000111000;
   42059: result <= 12'b111000111000;
   42060: result <= 12'b111000111000;
   42061: result <= 12'b111000111000;
   42062: result <= 12'b111000111000;
   42063: result <= 12'b111000111000;
   42064: result <= 12'b111000111001;
   42065: result <= 12'b111000111001;
   42066: result <= 12'b111000111001;
   42067: result <= 12'b111000111001;
   42068: result <= 12'b111000111001;
   42069: result <= 12'b111000111001;
   42070: result <= 12'b111000111001;
   42071: result <= 12'b111000111001;
   42072: result <= 12'b111000111010;
   42073: result <= 12'b111000111010;
   42074: result <= 12'b111000111010;
   42075: result <= 12'b111000111010;
   42076: result <= 12'b111000111010;
   42077: result <= 12'b111000111010;
   42078: result <= 12'b111000111010;
   42079: result <= 12'b111000111010;
   42080: result <= 12'b111000111011;
   42081: result <= 12'b111000111011;
   42082: result <= 12'b111000111011;
   42083: result <= 12'b111000111011;
   42084: result <= 12'b111000111011;
   42085: result <= 12'b111000111011;
   42086: result <= 12'b111000111011;
   42087: result <= 12'b111000111011;
   42088: result <= 12'b111000111100;
   42089: result <= 12'b111000111100;
   42090: result <= 12'b111000111100;
   42091: result <= 12'b111000111100;
   42092: result <= 12'b111000111100;
   42093: result <= 12'b111000111100;
   42094: result <= 12'b111000111100;
   42095: result <= 12'b111000111100;
   42096: result <= 12'b111000111100;
   42097: result <= 12'b111000111101;
   42098: result <= 12'b111000111101;
   42099: result <= 12'b111000111101;
   42100: result <= 12'b111000111101;
   42101: result <= 12'b111000111101;
   42102: result <= 12'b111000111101;
   42103: result <= 12'b111000111101;
   42104: result <= 12'b111000111101;
   42105: result <= 12'b111000111110;
   42106: result <= 12'b111000111110;
   42107: result <= 12'b111000111110;
   42108: result <= 12'b111000111110;
   42109: result <= 12'b111000111110;
   42110: result <= 12'b111000111110;
   42111: result <= 12'b111000111110;
   42112: result <= 12'b111000111110;
   42113: result <= 12'b111000111111;
   42114: result <= 12'b111000111111;
   42115: result <= 12'b111000111111;
   42116: result <= 12'b111000111111;
   42117: result <= 12'b111000111111;
   42118: result <= 12'b111000111111;
   42119: result <= 12'b111000111111;
   42120: result <= 12'b111000111111;
   42121: result <= 12'b111001000000;
   42122: result <= 12'b111001000000;
   42123: result <= 12'b111001000000;
   42124: result <= 12'b111001000000;
   42125: result <= 12'b111001000000;
   42126: result <= 12'b111001000000;
   42127: result <= 12'b111001000000;
   42128: result <= 12'b111001000000;
   42129: result <= 12'b111001000001;
   42130: result <= 12'b111001000001;
   42131: result <= 12'b111001000001;
   42132: result <= 12'b111001000001;
   42133: result <= 12'b111001000001;
   42134: result <= 12'b111001000001;
   42135: result <= 12'b111001000001;
   42136: result <= 12'b111001000001;
   42137: result <= 12'b111001000010;
   42138: result <= 12'b111001000010;
   42139: result <= 12'b111001000010;
   42140: result <= 12'b111001000010;
   42141: result <= 12'b111001000010;
   42142: result <= 12'b111001000010;
   42143: result <= 12'b111001000010;
   42144: result <= 12'b111001000010;
   42145: result <= 12'b111001000010;
   42146: result <= 12'b111001000011;
   42147: result <= 12'b111001000011;
   42148: result <= 12'b111001000011;
   42149: result <= 12'b111001000011;
   42150: result <= 12'b111001000011;
   42151: result <= 12'b111001000011;
   42152: result <= 12'b111001000011;
   42153: result <= 12'b111001000011;
   42154: result <= 12'b111001000100;
   42155: result <= 12'b111001000100;
   42156: result <= 12'b111001000100;
   42157: result <= 12'b111001000100;
   42158: result <= 12'b111001000100;
   42159: result <= 12'b111001000100;
   42160: result <= 12'b111001000100;
   42161: result <= 12'b111001000100;
   42162: result <= 12'b111001000101;
   42163: result <= 12'b111001000101;
   42164: result <= 12'b111001000101;
   42165: result <= 12'b111001000101;
   42166: result <= 12'b111001000101;
   42167: result <= 12'b111001000101;
   42168: result <= 12'b111001000101;
   42169: result <= 12'b111001000101;
   42170: result <= 12'b111001000110;
   42171: result <= 12'b111001000110;
   42172: result <= 12'b111001000110;
   42173: result <= 12'b111001000110;
   42174: result <= 12'b111001000110;
   42175: result <= 12'b111001000110;
   42176: result <= 12'b111001000110;
   42177: result <= 12'b111001000110;
   42178: result <= 12'b111001000111;
   42179: result <= 12'b111001000111;
   42180: result <= 12'b111001000111;
   42181: result <= 12'b111001000111;
   42182: result <= 12'b111001000111;
   42183: result <= 12'b111001000111;
   42184: result <= 12'b111001000111;
   42185: result <= 12'b111001000111;
   42186: result <= 12'b111001000111;
   42187: result <= 12'b111001001000;
   42188: result <= 12'b111001001000;
   42189: result <= 12'b111001001000;
   42190: result <= 12'b111001001000;
   42191: result <= 12'b111001001000;
   42192: result <= 12'b111001001000;
   42193: result <= 12'b111001001000;
   42194: result <= 12'b111001001000;
   42195: result <= 12'b111001001001;
   42196: result <= 12'b111001001001;
   42197: result <= 12'b111001001001;
   42198: result <= 12'b111001001001;
   42199: result <= 12'b111001001001;
   42200: result <= 12'b111001001001;
   42201: result <= 12'b111001001001;
   42202: result <= 12'b111001001001;
   42203: result <= 12'b111001001010;
   42204: result <= 12'b111001001010;
   42205: result <= 12'b111001001010;
   42206: result <= 12'b111001001010;
   42207: result <= 12'b111001001010;
   42208: result <= 12'b111001001010;
   42209: result <= 12'b111001001010;
   42210: result <= 12'b111001001010;
   42211: result <= 12'b111001001011;
   42212: result <= 12'b111001001011;
   42213: result <= 12'b111001001011;
   42214: result <= 12'b111001001011;
   42215: result <= 12'b111001001011;
   42216: result <= 12'b111001001011;
   42217: result <= 12'b111001001011;
   42218: result <= 12'b111001001011;
   42219: result <= 12'b111001001011;
   42220: result <= 12'b111001001100;
   42221: result <= 12'b111001001100;
   42222: result <= 12'b111001001100;
   42223: result <= 12'b111001001100;
   42224: result <= 12'b111001001100;
   42225: result <= 12'b111001001100;
   42226: result <= 12'b111001001100;
   42227: result <= 12'b111001001100;
   42228: result <= 12'b111001001101;
   42229: result <= 12'b111001001101;
   42230: result <= 12'b111001001101;
   42231: result <= 12'b111001001101;
   42232: result <= 12'b111001001101;
   42233: result <= 12'b111001001101;
   42234: result <= 12'b111001001101;
   42235: result <= 12'b111001001101;
   42236: result <= 12'b111001001110;
   42237: result <= 12'b111001001110;
   42238: result <= 12'b111001001110;
   42239: result <= 12'b111001001110;
   42240: result <= 12'b111001001110;
   42241: result <= 12'b111001001110;
   42242: result <= 12'b111001001110;
   42243: result <= 12'b111001001110;
   42244: result <= 12'b111001001111;
   42245: result <= 12'b111001001111;
   42246: result <= 12'b111001001111;
   42247: result <= 12'b111001001111;
   42248: result <= 12'b111001001111;
   42249: result <= 12'b111001001111;
   42250: result <= 12'b111001001111;
   42251: result <= 12'b111001001111;
   42252: result <= 12'b111001001111;
   42253: result <= 12'b111001010000;
   42254: result <= 12'b111001010000;
   42255: result <= 12'b111001010000;
   42256: result <= 12'b111001010000;
   42257: result <= 12'b111001010000;
   42258: result <= 12'b111001010000;
   42259: result <= 12'b111001010000;
   42260: result <= 12'b111001010000;
   42261: result <= 12'b111001010001;
   42262: result <= 12'b111001010001;
   42263: result <= 12'b111001010001;
   42264: result <= 12'b111001010001;
   42265: result <= 12'b111001010001;
   42266: result <= 12'b111001010001;
   42267: result <= 12'b111001010001;
   42268: result <= 12'b111001010001;
   42269: result <= 12'b111001010010;
   42270: result <= 12'b111001010010;
   42271: result <= 12'b111001010010;
   42272: result <= 12'b111001010010;
   42273: result <= 12'b111001010010;
   42274: result <= 12'b111001010010;
   42275: result <= 12'b111001010010;
   42276: result <= 12'b111001010010;
   42277: result <= 12'b111001010010;
   42278: result <= 12'b111001010011;
   42279: result <= 12'b111001010011;
   42280: result <= 12'b111001010011;
   42281: result <= 12'b111001010011;
   42282: result <= 12'b111001010011;
   42283: result <= 12'b111001010011;
   42284: result <= 12'b111001010011;
   42285: result <= 12'b111001010011;
   42286: result <= 12'b111001010100;
   42287: result <= 12'b111001010100;
   42288: result <= 12'b111001010100;
   42289: result <= 12'b111001010100;
   42290: result <= 12'b111001010100;
   42291: result <= 12'b111001010100;
   42292: result <= 12'b111001010100;
   42293: result <= 12'b111001010100;
   42294: result <= 12'b111001010101;
   42295: result <= 12'b111001010101;
   42296: result <= 12'b111001010101;
   42297: result <= 12'b111001010101;
   42298: result <= 12'b111001010101;
   42299: result <= 12'b111001010101;
   42300: result <= 12'b111001010101;
   42301: result <= 12'b111001010101;
   42302: result <= 12'b111001010101;
   42303: result <= 12'b111001010110;
   42304: result <= 12'b111001010110;
   42305: result <= 12'b111001010110;
   42306: result <= 12'b111001010110;
   42307: result <= 12'b111001010110;
   42308: result <= 12'b111001010110;
   42309: result <= 12'b111001010110;
   42310: result <= 12'b111001010110;
   42311: result <= 12'b111001010111;
   42312: result <= 12'b111001010111;
   42313: result <= 12'b111001010111;
   42314: result <= 12'b111001010111;
   42315: result <= 12'b111001010111;
   42316: result <= 12'b111001010111;
   42317: result <= 12'b111001010111;
   42318: result <= 12'b111001010111;
   42319: result <= 12'b111001011000;
   42320: result <= 12'b111001011000;
   42321: result <= 12'b111001011000;
   42322: result <= 12'b111001011000;
   42323: result <= 12'b111001011000;
   42324: result <= 12'b111001011000;
   42325: result <= 12'b111001011000;
   42326: result <= 12'b111001011000;
   42327: result <= 12'b111001011000;
   42328: result <= 12'b111001011001;
   42329: result <= 12'b111001011001;
   42330: result <= 12'b111001011001;
   42331: result <= 12'b111001011001;
   42332: result <= 12'b111001011001;
   42333: result <= 12'b111001011001;
   42334: result <= 12'b111001011001;
   42335: result <= 12'b111001011001;
   42336: result <= 12'b111001011010;
   42337: result <= 12'b111001011010;
   42338: result <= 12'b111001011010;
   42339: result <= 12'b111001011010;
   42340: result <= 12'b111001011010;
   42341: result <= 12'b111001011010;
   42342: result <= 12'b111001011010;
   42343: result <= 12'b111001011010;
   42344: result <= 12'b111001011011;
   42345: result <= 12'b111001011011;
   42346: result <= 12'b111001011011;
   42347: result <= 12'b111001011011;
   42348: result <= 12'b111001011011;
   42349: result <= 12'b111001011011;
   42350: result <= 12'b111001011011;
   42351: result <= 12'b111001011011;
   42352: result <= 12'b111001011011;
   42353: result <= 12'b111001011100;
   42354: result <= 12'b111001011100;
   42355: result <= 12'b111001011100;
   42356: result <= 12'b111001011100;
   42357: result <= 12'b111001011100;
   42358: result <= 12'b111001011100;
   42359: result <= 12'b111001011100;
   42360: result <= 12'b111001011100;
   42361: result <= 12'b111001011101;
   42362: result <= 12'b111001011101;
   42363: result <= 12'b111001011101;
   42364: result <= 12'b111001011101;
   42365: result <= 12'b111001011101;
   42366: result <= 12'b111001011101;
   42367: result <= 12'b111001011101;
   42368: result <= 12'b111001011101;
   42369: result <= 12'b111001011101;
   42370: result <= 12'b111001011110;
   42371: result <= 12'b111001011110;
   42372: result <= 12'b111001011110;
   42373: result <= 12'b111001011110;
   42374: result <= 12'b111001011110;
   42375: result <= 12'b111001011110;
   42376: result <= 12'b111001011110;
   42377: result <= 12'b111001011110;
   42378: result <= 12'b111001011111;
   42379: result <= 12'b111001011111;
   42380: result <= 12'b111001011111;
   42381: result <= 12'b111001011111;
   42382: result <= 12'b111001011111;
   42383: result <= 12'b111001011111;
   42384: result <= 12'b111001011111;
   42385: result <= 12'b111001011111;
   42386: result <= 12'b111001100000;
   42387: result <= 12'b111001100000;
   42388: result <= 12'b111001100000;
   42389: result <= 12'b111001100000;
   42390: result <= 12'b111001100000;
   42391: result <= 12'b111001100000;
   42392: result <= 12'b111001100000;
   42393: result <= 12'b111001100000;
   42394: result <= 12'b111001100000;
   42395: result <= 12'b111001100001;
   42396: result <= 12'b111001100001;
   42397: result <= 12'b111001100001;
   42398: result <= 12'b111001100001;
   42399: result <= 12'b111001100001;
   42400: result <= 12'b111001100001;
   42401: result <= 12'b111001100001;
   42402: result <= 12'b111001100001;
   42403: result <= 12'b111001100010;
   42404: result <= 12'b111001100010;
   42405: result <= 12'b111001100010;
   42406: result <= 12'b111001100010;
   42407: result <= 12'b111001100010;
   42408: result <= 12'b111001100010;
   42409: result <= 12'b111001100010;
   42410: result <= 12'b111001100010;
   42411: result <= 12'b111001100010;
   42412: result <= 12'b111001100011;
   42413: result <= 12'b111001100011;
   42414: result <= 12'b111001100011;
   42415: result <= 12'b111001100011;
   42416: result <= 12'b111001100011;
   42417: result <= 12'b111001100011;
   42418: result <= 12'b111001100011;
   42419: result <= 12'b111001100011;
   42420: result <= 12'b111001100100;
   42421: result <= 12'b111001100100;
   42422: result <= 12'b111001100100;
   42423: result <= 12'b111001100100;
   42424: result <= 12'b111001100100;
   42425: result <= 12'b111001100100;
   42426: result <= 12'b111001100100;
   42427: result <= 12'b111001100100;
   42428: result <= 12'b111001100100;
   42429: result <= 12'b111001100101;
   42430: result <= 12'b111001100101;
   42431: result <= 12'b111001100101;
   42432: result <= 12'b111001100101;
   42433: result <= 12'b111001100101;
   42434: result <= 12'b111001100101;
   42435: result <= 12'b111001100101;
   42436: result <= 12'b111001100101;
   42437: result <= 12'b111001100110;
   42438: result <= 12'b111001100110;
   42439: result <= 12'b111001100110;
   42440: result <= 12'b111001100110;
   42441: result <= 12'b111001100110;
   42442: result <= 12'b111001100110;
   42443: result <= 12'b111001100110;
   42444: result <= 12'b111001100110;
   42445: result <= 12'b111001100110;
   42446: result <= 12'b111001100111;
   42447: result <= 12'b111001100111;
   42448: result <= 12'b111001100111;
   42449: result <= 12'b111001100111;
   42450: result <= 12'b111001100111;
   42451: result <= 12'b111001100111;
   42452: result <= 12'b111001100111;
   42453: result <= 12'b111001100111;
   42454: result <= 12'b111001101000;
   42455: result <= 12'b111001101000;
   42456: result <= 12'b111001101000;
   42457: result <= 12'b111001101000;
   42458: result <= 12'b111001101000;
   42459: result <= 12'b111001101000;
   42460: result <= 12'b111001101000;
   42461: result <= 12'b111001101000;
   42462: result <= 12'b111001101000;
   42463: result <= 12'b111001101001;
   42464: result <= 12'b111001101001;
   42465: result <= 12'b111001101001;
   42466: result <= 12'b111001101001;
   42467: result <= 12'b111001101001;
   42468: result <= 12'b111001101001;
   42469: result <= 12'b111001101001;
   42470: result <= 12'b111001101001;
   42471: result <= 12'b111001101010;
   42472: result <= 12'b111001101010;
   42473: result <= 12'b111001101010;
   42474: result <= 12'b111001101010;
   42475: result <= 12'b111001101010;
   42476: result <= 12'b111001101010;
   42477: result <= 12'b111001101010;
   42478: result <= 12'b111001101010;
   42479: result <= 12'b111001101010;
   42480: result <= 12'b111001101011;
   42481: result <= 12'b111001101011;
   42482: result <= 12'b111001101011;
   42483: result <= 12'b111001101011;
   42484: result <= 12'b111001101011;
   42485: result <= 12'b111001101011;
   42486: result <= 12'b111001101011;
   42487: result <= 12'b111001101011;
   42488: result <= 12'b111001101100;
   42489: result <= 12'b111001101100;
   42490: result <= 12'b111001101100;
   42491: result <= 12'b111001101100;
   42492: result <= 12'b111001101100;
   42493: result <= 12'b111001101100;
   42494: result <= 12'b111001101100;
   42495: result <= 12'b111001101100;
   42496: result <= 12'b111001101100;
   42497: result <= 12'b111001101101;
   42498: result <= 12'b111001101101;
   42499: result <= 12'b111001101101;
   42500: result <= 12'b111001101101;
   42501: result <= 12'b111001101101;
   42502: result <= 12'b111001101101;
   42503: result <= 12'b111001101101;
   42504: result <= 12'b111001101101;
   42505: result <= 12'b111001101110;
   42506: result <= 12'b111001101110;
   42507: result <= 12'b111001101110;
   42508: result <= 12'b111001101110;
   42509: result <= 12'b111001101110;
   42510: result <= 12'b111001101110;
   42511: result <= 12'b111001101110;
   42512: result <= 12'b111001101110;
   42513: result <= 12'b111001101110;
   42514: result <= 12'b111001101111;
   42515: result <= 12'b111001101111;
   42516: result <= 12'b111001101111;
   42517: result <= 12'b111001101111;
   42518: result <= 12'b111001101111;
   42519: result <= 12'b111001101111;
   42520: result <= 12'b111001101111;
   42521: result <= 12'b111001101111;
   42522: result <= 12'b111001110000;
   42523: result <= 12'b111001110000;
   42524: result <= 12'b111001110000;
   42525: result <= 12'b111001110000;
   42526: result <= 12'b111001110000;
   42527: result <= 12'b111001110000;
   42528: result <= 12'b111001110000;
   42529: result <= 12'b111001110000;
   42530: result <= 12'b111001110000;
   42531: result <= 12'b111001110001;
   42532: result <= 12'b111001110001;
   42533: result <= 12'b111001110001;
   42534: result <= 12'b111001110001;
   42535: result <= 12'b111001110001;
   42536: result <= 12'b111001110001;
   42537: result <= 12'b111001110001;
   42538: result <= 12'b111001110001;
   42539: result <= 12'b111001110001;
   42540: result <= 12'b111001110010;
   42541: result <= 12'b111001110010;
   42542: result <= 12'b111001110010;
   42543: result <= 12'b111001110010;
   42544: result <= 12'b111001110010;
   42545: result <= 12'b111001110010;
   42546: result <= 12'b111001110010;
   42547: result <= 12'b111001110010;
   42548: result <= 12'b111001110011;
   42549: result <= 12'b111001110011;
   42550: result <= 12'b111001110011;
   42551: result <= 12'b111001110011;
   42552: result <= 12'b111001110011;
   42553: result <= 12'b111001110011;
   42554: result <= 12'b111001110011;
   42555: result <= 12'b111001110011;
   42556: result <= 12'b111001110011;
   42557: result <= 12'b111001110100;
   42558: result <= 12'b111001110100;
   42559: result <= 12'b111001110100;
   42560: result <= 12'b111001110100;
   42561: result <= 12'b111001110100;
   42562: result <= 12'b111001110100;
   42563: result <= 12'b111001110100;
   42564: result <= 12'b111001110100;
   42565: result <= 12'b111001110101;
   42566: result <= 12'b111001110101;
   42567: result <= 12'b111001110101;
   42568: result <= 12'b111001110101;
   42569: result <= 12'b111001110101;
   42570: result <= 12'b111001110101;
   42571: result <= 12'b111001110101;
   42572: result <= 12'b111001110101;
   42573: result <= 12'b111001110101;
   42574: result <= 12'b111001110110;
   42575: result <= 12'b111001110110;
   42576: result <= 12'b111001110110;
   42577: result <= 12'b111001110110;
   42578: result <= 12'b111001110110;
   42579: result <= 12'b111001110110;
   42580: result <= 12'b111001110110;
   42581: result <= 12'b111001110110;
   42582: result <= 12'b111001110110;
   42583: result <= 12'b111001110111;
   42584: result <= 12'b111001110111;
   42585: result <= 12'b111001110111;
   42586: result <= 12'b111001110111;
   42587: result <= 12'b111001110111;
   42588: result <= 12'b111001110111;
   42589: result <= 12'b111001110111;
   42590: result <= 12'b111001110111;
   42591: result <= 12'b111001111000;
   42592: result <= 12'b111001111000;
   42593: result <= 12'b111001111000;
   42594: result <= 12'b111001111000;
   42595: result <= 12'b111001111000;
   42596: result <= 12'b111001111000;
   42597: result <= 12'b111001111000;
   42598: result <= 12'b111001111000;
   42599: result <= 12'b111001111000;
   42600: result <= 12'b111001111001;
   42601: result <= 12'b111001111001;
   42602: result <= 12'b111001111001;
   42603: result <= 12'b111001111001;
   42604: result <= 12'b111001111001;
   42605: result <= 12'b111001111001;
   42606: result <= 12'b111001111001;
   42607: result <= 12'b111001111001;
   42608: result <= 12'b111001111001;
   42609: result <= 12'b111001111010;
   42610: result <= 12'b111001111010;
   42611: result <= 12'b111001111010;
   42612: result <= 12'b111001111010;
   42613: result <= 12'b111001111010;
   42614: result <= 12'b111001111010;
   42615: result <= 12'b111001111010;
   42616: result <= 12'b111001111010;
   42617: result <= 12'b111001111011;
   42618: result <= 12'b111001111011;
   42619: result <= 12'b111001111011;
   42620: result <= 12'b111001111011;
   42621: result <= 12'b111001111011;
   42622: result <= 12'b111001111011;
   42623: result <= 12'b111001111011;
   42624: result <= 12'b111001111011;
   42625: result <= 12'b111001111011;
   42626: result <= 12'b111001111100;
   42627: result <= 12'b111001111100;
   42628: result <= 12'b111001111100;
   42629: result <= 12'b111001111100;
   42630: result <= 12'b111001111100;
   42631: result <= 12'b111001111100;
   42632: result <= 12'b111001111100;
   42633: result <= 12'b111001111100;
   42634: result <= 12'b111001111100;
   42635: result <= 12'b111001111101;
   42636: result <= 12'b111001111101;
   42637: result <= 12'b111001111101;
   42638: result <= 12'b111001111101;
   42639: result <= 12'b111001111101;
   42640: result <= 12'b111001111101;
   42641: result <= 12'b111001111101;
   42642: result <= 12'b111001111101;
   42643: result <= 12'b111001111101;
   42644: result <= 12'b111001111110;
   42645: result <= 12'b111001111110;
   42646: result <= 12'b111001111110;
   42647: result <= 12'b111001111110;
   42648: result <= 12'b111001111110;
   42649: result <= 12'b111001111110;
   42650: result <= 12'b111001111110;
   42651: result <= 12'b111001111110;
   42652: result <= 12'b111001111111;
   42653: result <= 12'b111001111111;
   42654: result <= 12'b111001111111;
   42655: result <= 12'b111001111111;
   42656: result <= 12'b111001111111;
   42657: result <= 12'b111001111111;
   42658: result <= 12'b111001111111;
   42659: result <= 12'b111001111111;
   42660: result <= 12'b111001111111;
   42661: result <= 12'b111010000000;
   42662: result <= 12'b111010000000;
   42663: result <= 12'b111010000000;
   42664: result <= 12'b111010000000;
   42665: result <= 12'b111010000000;
   42666: result <= 12'b111010000000;
   42667: result <= 12'b111010000000;
   42668: result <= 12'b111010000000;
   42669: result <= 12'b111010000000;
   42670: result <= 12'b111010000001;
   42671: result <= 12'b111010000001;
   42672: result <= 12'b111010000001;
   42673: result <= 12'b111010000001;
   42674: result <= 12'b111010000001;
   42675: result <= 12'b111010000001;
   42676: result <= 12'b111010000001;
   42677: result <= 12'b111010000001;
   42678: result <= 12'b111010000010;
   42679: result <= 12'b111010000010;
   42680: result <= 12'b111010000010;
   42681: result <= 12'b111010000010;
   42682: result <= 12'b111010000010;
   42683: result <= 12'b111010000010;
   42684: result <= 12'b111010000010;
   42685: result <= 12'b111010000010;
   42686: result <= 12'b111010000010;
   42687: result <= 12'b111010000011;
   42688: result <= 12'b111010000011;
   42689: result <= 12'b111010000011;
   42690: result <= 12'b111010000011;
   42691: result <= 12'b111010000011;
   42692: result <= 12'b111010000011;
   42693: result <= 12'b111010000011;
   42694: result <= 12'b111010000011;
   42695: result <= 12'b111010000011;
   42696: result <= 12'b111010000100;
   42697: result <= 12'b111010000100;
   42698: result <= 12'b111010000100;
   42699: result <= 12'b111010000100;
   42700: result <= 12'b111010000100;
   42701: result <= 12'b111010000100;
   42702: result <= 12'b111010000100;
   42703: result <= 12'b111010000100;
   42704: result <= 12'b111010000100;
   42705: result <= 12'b111010000101;
   42706: result <= 12'b111010000101;
   42707: result <= 12'b111010000101;
   42708: result <= 12'b111010000101;
   42709: result <= 12'b111010000101;
   42710: result <= 12'b111010000101;
   42711: result <= 12'b111010000101;
   42712: result <= 12'b111010000101;
   42713: result <= 12'b111010000101;
   42714: result <= 12'b111010000110;
   42715: result <= 12'b111010000110;
   42716: result <= 12'b111010000110;
   42717: result <= 12'b111010000110;
   42718: result <= 12'b111010000110;
   42719: result <= 12'b111010000110;
   42720: result <= 12'b111010000110;
   42721: result <= 12'b111010000110;
   42722: result <= 12'b111010000111;
   42723: result <= 12'b111010000111;
   42724: result <= 12'b111010000111;
   42725: result <= 12'b111010000111;
   42726: result <= 12'b111010000111;
   42727: result <= 12'b111010000111;
   42728: result <= 12'b111010000111;
   42729: result <= 12'b111010000111;
   42730: result <= 12'b111010000111;
   42731: result <= 12'b111010001000;
   42732: result <= 12'b111010001000;
   42733: result <= 12'b111010001000;
   42734: result <= 12'b111010001000;
   42735: result <= 12'b111010001000;
   42736: result <= 12'b111010001000;
   42737: result <= 12'b111010001000;
   42738: result <= 12'b111010001000;
   42739: result <= 12'b111010001000;
   42740: result <= 12'b111010001001;
   42741: result <= 12'b111010001001;
   42742: result <= 12'b111010001001;
   42743: result <= 12'b111010001001;
   42744: result <= 12'b111010001001;
   42745: result <= 12'b111010001001;
   42746: result <= 12'b111010001001;
   42747: result <= 12'b111010001001;
   42748: result <= 12'b111010001001;
   42749: result <= 12'b111010001010;
   42750: result <= 12'b111010001010;
   42751: result <= 12'b111010001010;
   42752: result <= 12'b111010001010;
   42753: result <= 12'b111010001010;
   42754: result <= 12'b111010001010;
   42755: result <= 12'b111010001010;
   42756: result <= 12'b111010001010;
   42757: result <= 12'b111010001010;
   42758: result <= 12'b111010001011;
   42759: result <= 12'b111010001011;
   42760: result <= 12'b111010001011;
   42761: result <= 12'b111010001011;
   42762: result <= 12'b111010001011;
   42763: result <= 12'b111010001011;
   42764: result <= 12'b111010001011;
   42765: result <= 12'b111010001011;
   42766: result <= 12'b111010001011;
   42767: result <= 12'b111010001100;
   42768: result <= 12'b111010001100;
   42769: result <= 12'b111010001100;
   42770: result <= 12'b111010001100;
   42771: result <= 12'b111010001100;
   42772: result <= 12'b111010001100;
   42773: result <= 12'b111010001100;
   42774: result <= 12'b111010001100;
   42775: result <= 12'b111010001101;
   42776: result <= 12'b111010001101;
   42777: result <= 12'b111010001101;
   42778: result <= 12'b111010001101;
   42779: result <= 12'b111010001101;
   42780: result <= 12'b111010001101;
   42781: result <= 12'b111010001101;
   42782: result <= 12'b111010001101;
   42783: result <= 12'b111010001101;
   42784: result <= 12'b111010001110;
   42785: result <= 12'b111010001110;
   42786: result <= 12'b111010001110;
   42787: result <= 12'b111010001110;
   42788: result <= 12'b111010001110;
   42789: result <= 12'b111010001110;
   42790: result <= 12'b111010001110;
   42791: result <= 12'b111010001110;
   42792: result <= 12'b111010001110;
   42793: result <= 12'b111010001111;
   42794: result <= 12'b111010001111;
   42795: result <= 12'b111010001111;
   42796: result <= 12'b111010001111;
   42797: result <= 12'b111010001111;
   42798: result <= 12'b111010001111;
   42799: result <= 12'b111010001111;
   42800: result <= 12'b111010001111;
   42801: result <= 12'b111010001111;
   42802: result <= 12'b111010010000;
   42803: result <= 12'b111010010000;
   42804: result <= 12'b111010010000;
   42805: result <= 12'b111010010000;
   42806: result <= 12'b111010010000;
   42807: result <= 12'b111010010000;
   42808: result <= 12'b111010010000;
   42809: result <= 12'b111010010000;
   42810: result <= 12'b111010010000;
   42811: result <= 12'b111010010001;
   42812: result <= 12'b111010010001;
   42813: result <= 12'b111010010001;
   42814: result <= 12'b111010010001;
   42815: result <= 12'b111010010001;
   42816: result <= 12'b111010010001;
   42817: result <= 12'b111010010001;
   42818: result <= 12'b111010010001;
   42819: result <= 12'b111010010001;
   42820: result <= 12'b111010010010;
   42821: result <= 12'b111010010010;
   42822: result <= 12'b111010010010;
   42823: result <= 12'b111010010010;
   42824: result <= 12'b111010010010;
   42825: result <= 12'b111010010010;
   42826: result <= 12'b111010010010;
   42827: result <= 12'b111010010010;
   42828: result <= 12'b111010010010;
   42829: result <= 12'b111010010011;
   42830: result <= 12'b111010010011;
   42831: result <= 12'b111010010011;
   42832: result <= 12'b111010010011;
   42833: result <= 12'b111010010011;
   42834: result <= 12'b111010010011;
   42835: result <= 12'b111010010011;
   42836: result <= 12'b111010010011;
   42837: result <= 12'b111010010011;
   42838: result <= 12'b111010010100;
   42839: result <= 12'b111010010100;
   42840: result <= 12'b111010010100;
   42841: result <= 12'b111010010100;
   42842: result <= 12'b111010010100;
   42843: result <= 12'b111010010100;
   42844: result <= 12'b111010010100;
   42845: result <= 12'b111010010100;
   42846: result <= 12'b111010010100;
   42847: result <= 12'b111010010101;
   42848: result <= 12'b111010010101;
   42849: result <= 12'b111010010101;
   42850: result <= 12'b111010010101;
   42851: result <= 12'b111010010101;
   42852: result <= 12'b111010010101;
   42853: result <= 12'b111010010101;
   42854: result <= 12'b111010010101;
   42855: result <= 12'b111010010101;
   42856: result <= 12'b111010010110;
   42857: result <= 12'b111010010110;
   42858: result <= 12'b111010010110;
   42859: result <= 12'b111010010110;
   42860: result <= 12'b111010010110;
   42861: result <= 12'b111010010110;
   42862: result <= 12'b111010010110;
   42863: result <= 12'b111010010110;
   42864: result <= 12'b111010010110;
   42865: result <= 12'b111010010111;
   42866: result <= 12'b111010010111;
   42867: result <= 12'b111010010111;
   42868: result <= 12'b111010010111;
   42869: result <= 12'b111010010111;
   42870: result <= 12'b111010010111;
   42871: result <= 12'b111010010111;
   42872: result <= 12'b111010010111;
   42873: result <= 12'b111010010111;
   42874: result <= 12'b111010011000;
   42875: result <= 12'b111010011000;
   42876: result <= 12'b111010011000;
   42877: result <= 12'b111010011000;
   42878: result <= 12'b111010011000;
   42879: result <= 12'b111010011000;
   42880: result <= 12'b111010011000;
   42881: result <= 12'b111010011000;
   42882: result <= 12'b111010011000;
   42883: result <= 12'b111010011001;
   42884: result <= 12'b111010011001;
   42885: result <= 12'b111010011001;
   42886: result <= 12'b111010011001;
   42887: result <= 12'b111010011001;
   42888: result <= 12'b111010011001;
   42889: result <= 12'b111010011001;
   42890: result <= 12'b111010011001;
   42891: result <= 12'b111010011001;
   42892: result <= 12'b111010011010;
   42893: result <= 12'b111010011010;
   42894: result <= 12'b111010011010;
   42895: result <= 12'b111010011010;
   42896: result <= 12'b111010011010;
   42897: result <= 12'b111010011010;
   42898: result <= 12'b111010011010;
   42899: result <= 12'b111010011010;
   42900: result <= 12'b111010011010;
   42901: result <= 12'b111010011011;
   42902: result <= 12'b111010011011;
   42903: result <= 12'b111010011011;
   42904: result <= 12'b111010011011;
   42905: result <= 12'b111010011011;
   42906: result <= 12'b111010011011;
   42907: result <= 12'b111010011011;
   42908: result <= 12'b111010011011;
   42909: result <= 12'b111010011011;
   42910: result <= 12'b111010011100;
   42911: result <= 12'b111010011100;
   42912: result <= 12'b111010011100;
   42913: result <= 12'b111010011100;
   42914: result <= 12'b111010011100;
   42915: result <= 12'b111010011100;
   42916: result <= 12'b111010011100;
   42917: result <= 12'b111010011100;
   42918: result <= 12'b111010011100;
   42919: result <= 12'b111010011101;
   42920: result <= 12'b111010011101;
   42921: result <= 12'b111010011101;
   42922: result <= 12'b111010011101;
   42923: result <= 12'b111010011101;
   42924: result <= 12'b111010011101;
   42925: result <= 12'b111010011101;
   42926: result <= 12'b111010011101;
   42927: result <= 12'b111010011101;
   42928: result <= 12'b111010011110;
   42929: result <= 12'b111010011110;
   42930: result <= 12'b111010011110;
   42931: result <= 12'b111010011110;
   42932: result <= 12'b111010011110;
   42933: result <= 12'b111010011110;
   42934: result <= 12'b111010011110;
   42935: result <= 12'b111010011110;
   42936: result <= 12'b111010011110;
   42937: result <= 12'b111010011111;
   42938: result <= 12'b111010011111;
   42939: result <= 12'b111010011111;
   42940: result <= 12'b111010011111;
   42941: result <= 12'b111010011111;
   42942: result <= 12'b111010011111;
   42943: result <= 12'b111010011111;
   42944: result <= 12'b111010011111;
   42945: result <= 12'b111010011111;
   42946: result <= 12'b111010100000;
   42947: result <= 12'b111010100000;
   42948: result <= 12'b111010100000;
   42949: result <= 12'b111010100000;
   42950: result <= 12'b111010100000;
   42951: result <= 12'b111010100000;
   42952: result <= 12'b111010100000;
   42953: result <= 12'b111010100000;
   42954: result <= 12'b111010100000;
   42955: result <= 12'b111010100001;
   42956: result <= 12'b111010100001;
   42957: result <= 12'b111010100001;
   42958: result <= 12'b111010100001;
   42959: result <= 12'b111010100001;
   42960: result <= 12'b111010100001;
   42961: result <= 12'b111010100001;
   42962: result <= 12'b111010100001;
   42963: result <= 12'b111010100001;
   42964: result <= 12'b111010100010;
   42965: result <= 12'b111010100010;
   42966: result <= 12'b111010100010;
   42967: result <= 12'b111010100010;
   42968: result <= 12'b111010100010;
   42969: result <= 12'b111010100010;
   42970: result <= 12'b111010100010;
   42971: result <= 12'b111010100010;
   42972: result <= 12'b111010100010;
   42973: result <= 12'b111010100011;
   42974: result <= 12'b111010100011;
   42975: result <= 12'b111010100011;
   42976: result <= 12'b111010100011;
   42977: result <= 12'b111010100011;
   42978: result <= 12'b111010100011;
   42979: result <= 12'b111010100011;
   42980: result <= 12'b111010100011;
   42981: result <= 12'b111010100011;
   42982: result <= 12'b111010100100;
   42983: result <= 12'b111010100100;
   42984: result <= 12'b111010100100;
   42985: result <= 12'b111010100100;
   42986: result <= 12'b111010100100;
   42987: result <= 12'b111010100100;
   42988: result <= 12'b111010100100;
   42989: result <= 12'b111010100100;
   42990: result <= 12'b111010100100;
   42991: result <= 12'b111010100100;
   42992: result <= 12'b111010100101;
   42993: result <= 12'b111010100101;
   42994: result <= 12'b111010100101;
   42995: result <= 12'b111010100101;
   42996: result <= 12'b111010100101;
   42997: result <= 12'b111010100101;
   42998: result <= 12'b111010100101;
   42999: result <= 12'b111010100101;
   43000: result <= 12'b111010100101;
   43001: result <= 12'b111010100110;
   43002: result <= 12'b111010100110;
   43003: result <= 12'b111010100110;
   43004: result <= 12'b111010100110;
   43005: result <= 12'b111010100110;
   43006: result <= 12'b111010100110;
   43007: result <= 12'b111010100110;
   43008: result <= 12'b111010100110;
   43009: result <= 12'b111010100110;
   43010: result <= 12'b111010100111;
   43011: result <= 12'b111010100111;
   43012: result <= 12'b111010100111;
   43013: result <= 12'b111010100111;
   43014: result <= 12'b111010100111;
   43015: result <= 12'b111010100111;
   43016: result <= 12'b111010100111;
   43017: result <= 12'b111010100111;
   43018: result <= 12'b111010100111;
   43019: result <= 12'b111010101000;
   43020: result <= 12'b111010101000;
   43021: result <= 12'b111010101000;
   43022: result <= 12'b111010101000;
   43023: result <= 12'b111010101000;
   43024: result <= 12'b111010101000;
   43025: result <= 12'b111010101000;
   43026: result <= 12'b111010101000;
   43027: result <= 12'b111010101000;
   43028: result <= 12'b111010101001;
   43029: result <= 12'b111010101001;
   43030: result <= 12'b111010101001;
   43031: result <= 12'b111010101001;
   43032: result <= 12'b111010101001;
   43033: result <= 12'b111010101001;
   43034: result <= 12'b111010101001;
   43035: result <= 12'b111010101001;
   43036: result <= 12'b111010101001;
   43037: result <= 12'b111010101010;
   43038: result <= 12'b111010101010;
   43039: result <= 12'b111010101010;
   43040: result <= 12'b111010101010;
   43041: result <= 12'b111010101010;
   43042: result <= 12'b111010101010;
   43043: result <= 12'b111010101010;
   43044: result <= 12'b111010101010;
   43045: result <= 12'b111010101010;
   43046: result <= 12'b111010101010;
   43047: result <= 12'b111010101011;
   43048: result <= 12'b111010101011;
   43049: result <= 12'b111010101011;
   43050: result <= 12'b111010101011;
   43051: result <= 12'b111010101011;
   43052: result <= 12'b111010101011;
   43053: result <= 12'b111010101011;
   43054: result <= 12'b111010101011;
   43055: result <= 12'b111010101011;
   43056: result <= 12'b111010101100;
   43057: result <= 12'b111010101100;
   43058: result <= 12'b111010101100;
   43059: result <= 12'b111010101100;
   43060: result <= 12'b111010101100;
   43061: result <= 12'b111010101100;
   43062: result <= 12'b111010101100;
   43063: result <= 12'b111010101100;
   43064: result <= 12'b111010101100;
   43065: result <= 12'b111010101101;
   43066: result <= 12'b111010101101;
   43067: result <= 12'b111010101101;
   43068: result <= 12'b111010101101;
   43069: result <= 12'b111010101101;
   43070: result <= 12'b111010101101;
   43071: result <= 12'b111010101101;
   43072: result <= 12'b111010101101;
   43073: result <= 12'b111010101101;
   43074: result <= 12'b111010101110;
   43075: result <= 12'b111010101110;
   43076: result <= 12'b111010101110;
   43077: result <= 12'b111010101110;
   43078: result <= 12'b111010101110;
   43079: result <= 12'b111010101110;
   43080: result <= 12'b111010101110;
   43081: result <= 12'b111010101110;
   43082: result <= 12'b111010101110;
   43083: result <= 12'b111010101110;
   43084: result <= 12'b111010101111;
   43085: result <= 12'b111010101111;
   43086: result <= 12'b111010101111;
   43087: result <= 12'b111010101111;
   43088: result <= 12'b111010101111;
   43089: result <= 12'b111010101111;
   43090: result <= 12'b111010101111;
   43091: result <= 12'b111010101111;
   43092: result <= 12'b111010101111;
   43093: result <= 12'b111010110000;
   43094: result <= 12'b111010110000;
   43095: result <= 12'b111010110000;
   43096: result <= 12'b111010110000;
   43097: result <= 12'b111010110000;
   43098: result <= 12'b111010110000;
   43099: result <= 12'b111010110000;
   43100: result <= 12'b111010110000;
   43101: result <= 12'b111010110000;
   43102: result <= 12'b111010110001;
   43103: result <= 12'b111010110001;
   43104: result <= 12'b111010110001;
   43105: result <= 12'b111010110001;
   43106: result <= 12'b111010110001;
   43107: result <= 12'b111010110001;
   43108: result <= 12'b111010110001;
   43109: result <= 12'b111010110001;
   43110: result <= 12'b111010110001;
   43111: result <= 12'b111010110010;
   43112: result <= 12'b111010110010;
   43113: result <= 12'b111010110010;
   43114: result <= 12'b111010110010;
   43115: result <= 12'b111010110010;
   43116: result <= 12'b111010110010;
   43117: result <= 12'b111010110010;
   43118: result <= 12'b111010110010;
   43119: result <= 12'b111010110010;
   43120: result <= 12'b111010110010;
   43121: result <= 12'b111010110011;
   43122: result <= 12'b111010110011;
   43123: result <= 12'b111010110011;
   43124: result <= 12'b111010110011;
   43125: result <= 12'b111010110011;
   43126: result <= 12'b111010110011;
   43127: result <= 12'b111010110011;
   43128: result <= 12'b111010110011;
   43129: result <= 12'b111010110011;
   43130: result <= 12'b111010110100;
   43131: result <= 12'b111010110100;
   43132: result <= 12'b111010110100;
   43133: result <= 12'b111010110100;
   43134: result <= 12'b111010110100;
   43135: result <= 12'b111010110100;
   43136: result <= 12'b111010110100;
   43137: result <= 12'b111010110100;
   43138: result <= 12'b111010110100;
   43139: result <= 12'b111010110101;
   43140: result <= 12'b111010110101;
   43141: result <= 12'b111010110101;
   43142: result <= 12'b111010110101;
   43143: result <= 12'b111010110101;
   43144: result <= 12'b111010110101;
   43145: result <= 12'b111010110101;
   43146: result <= 12'b111010110101;
   43147: result <= 12'b111010110101;
   43148: result <= 12'b111010110101;
   43149: result <= 12'b111010110110;
   43150: result <= 12'b111010110110;
   43151: result <= 12'b111010110110;
   43152: result <= 12'b111010110110;
   43153: result <= 12'b111010110110;
   43154: result <= 12'b111010110110;
   43155: result <= 12'b111010110110;
   43156: result <= 12'b111010110110;
   43157: result <= 12'b111010110110;
   43158: result <= 12'b111010110111;
   43159: result <= 12'b111010110111;
   43160: result <= 12'b111010110111;
   43161: result <= 12'b111010110111;
   43162: result <= 12'b111010110111;
   43163: result <= 12'b111010110111;
   43164: result <= 12'b111010110111;
   43165: result <= 12'b111010110111;
   43166: result <= 12'b111010110111;
   43167: result <= 12'b111010110111;
   43168: result <= 12'b111010111000;
   43169: result <= 12'b111010111000;
   43170: result <= 12'b111010111000;
   43171: result <= 12'b111010111000;
   43172: result <= 12'b111010111000;
   43173: result <= 12'b111010111000;
   43174: result <= 12'b111010111000;
   43175: result <= 12'b111010111000;
   43176: result <= 12'b111010111000;
   43177: result <= 12'b111010111001;
   43178: result <= 12'b111010111001;
   43179: result <= 12'b111010111001;
   43180: result <= 12'b111010111001;
   43181: result <= 12'b111010111001;
   43182: result <= 12'b111010111001;
   43183: result <= 12'b111010111001;
   43184: result <= 12'b111010111001;
   43185: result <= 12'b111010111001;
   43186: result <= 12'b111010111010;
   43187: result <= 12'b111010111010;
   43188: result <= 12'b111010111010;
   43189: result <= 12'b111010111010;
   43190: result <= 12'b111010111010;
   43191: result <= 12'b111010111010;
   43192: result <= 12'b111010111010;
   43193: result <= 12'b111010111010;
   43194: result <= 12'b111010111010;
   43195: result <= 12'b111010111010;
   43196: result <= 12'b111010111011;
   43197: result <= 12'b111010111011;
   43198: result <= 12'b111010111011;
   43199: result <= 12'b111010111011;
   43200: result <= 12'b111010111011;
   43201: result <= 12'b111010111011;
   43202: result <= 12'b111010111011;
   43203: result <= 12'b111010111011;
   43204: result <= 12'b111010111011;
   43205: result <= 12'b111010111100;
   43206: result <= 12'b111010111100;
   43207: result <= 12'b111010111100;
   43208: result <= 12'b111010111100;
   43209: result <= 12'b111010111100;
   43210: result <= 12'b111010111100;
   43211: result <= 12'b111010111100;
   43212: result <= 12'b111010111100;
   43213: result <= 12'b111010111100;
   43214: result <= 12'b111010111100;
   43215: result <= 12'b111010111101;
   43216: result <= 12'b111010111101;
   43217: result <= 12'b111010111101;
   43218: result <= 12'b111010111101;
   43219: result <= 12'b111010111101;
   43220: result <= 12'b111010111101;
   43221: result <= 12'b111010111101;
   43222: result <= 12'b111010111101;
   43223: result <= 12'b111010111101;
   43224: result <= 12'b111010111110;
   43225: result <= 12'b111010111110;
   43226: result <= 12'b111010111110;
   43227: result <= 12'b111010111110;
   43228: result <= 12'b111010111110;
   43229: result <= 12'b111010111110;
   43230: result <= 12'b111010111110;
   43231: result <= 12'b111010111110;
   43232: result <= 12'b111010111110;
   43233: result <= 12'b111010111110;
   43234: result <= 12'b111010111111;
   43235: result <= 12'b111010111111;
   43236: result <= 12'b111010111111;
   43237: result <= 12'b111010111111;
   43238: result <= 12'b111010111111;
   43239: result <= 12'b111010111111;
   43240: result <= 12'b111010111111;
   43241: result <= 12'b111010111111;
   43242: result <= 12'b111010111111;
   43243: result <= 12'b111011000000;
   43244: result <= 12'b111011000000;
   43245: result <= 12'b111011000000;
   43246: result <= 12'b111011000000;
   43247: result <= 12'b111011000000;
   43248: result <= 12'b111011000000;
   43249: result <= 12'b111011000000;
   43250: result <= 12'b111011000000;
   43251: result <= 12'b111011000000;
   43252: result <= 12'b111011000000;
   43253: result <= 12'b111011000001;
   43254: result <= 12'b111011000001;
   43255: result <= 12'b111011000001;
   43256: result <= 12'b111011000001;
   43257: result <= 12'b111011000001;
   43258: result <= 12'b111011000001;
   43259: result <= 12'b111011000001;
   43260: result <= 12'b111011000001;
   43261: result <= 12'b111011000001;
   43262: result <= 12'b111011000010;
   43263: result <= 12'b111011000010;
   43264: result <= 12'b111011000010;
   43265: result <= 12'b111011000010;
   43266: result <= 12'b111011000010;
   43267: result <= 12'b111011000010;
   43268: result <= 12'b111011000010;
   43269: result <= 12'b111011000010;
   43270: result <= 12'b111011000010;
   43271: result <= 12'b111011000010;
   43272: result <= 12'b111011000011;
   43273: result <= 12'b111011000011;
   43274: result <= 12'b111011000011;
   43275: result <= 12'b111011000011;
   43276: result <= 12'b111011000011;
   43277: result <= 12'b111011000011;
   43278: result <= 12'b111011000011;
   43279: result <= 12'b111011000011;
   43280: result <= 12'b111011000011;
   43281: result <= 12'b111011000100;
   43282: result <= 12'b111011000100;
   43283: result <= 12'b111011000100;
   43284: result <= 12'b111011000100;
   43285: result <= 12'b111011000100;
   43286: result <= 12'b111011000100;
   43287: result <= 12'b111011000100;
   43288: result <= 12'b111011000100;
   43289: result <= 12'b111011000100;
   43290: result <= 12'b111011000100;
   43291: result <= 12'b111011000101;
   43292: result <= 12'b111011000101;
   43293: result <= 12'b111011000101;
   43294: result <= 12'b111011000101;
   43295: result <= 12'b111011000101;
   43296: result <= 12'b111011000101;
   43297: result <= 12'b111011000101;
   43298: result <= 12'b111011000101;
   43299: result <= 12'b111011000101;
   43300: result <= 12'b111011000110;
   43301: result <= 12'b111011000110;
   43302: result <= 12'b111011000110;
   43303: result <= 12'b111011000110;
   43304: result <= 12'b111011000110;
   43305: result <= 12'b111011000110;
   43306: result <= 12'b111011000110;
   43307: result <= 12'b111011000110;
   43308: result <= 12'b111011000110;
   43309: result <= 12'b111011000110;
   43310: result <= 12'b111011000111;
   43311: result <= 12'b111011000111;
   43312: result <= 12'b111011000111;
   43313: result <= 12'b111011000111;
   43314: result <= 12'b111011000111;
   43315: result <= 12'b111011000111;
   43316: result <= 12'b111011000111;
   43317: result <= 12'b111011000111;
   43318: result <= 12'b111011000111;
   43319: result <= 12'b111011001000;
   43320: result <= 12'b111011001000;
   43321: result <= 12'b111011001000;
   43322: result <= 12'b111011001000;
   43323: result <= 12'b111011001000;
   43324: result <= 12'b111011001000;
   43325: result <= 12'b111011001000;
   43326: result <= 12'b111011001000;
   43327: result <= 12'b111011001000;
   43328: result <= 12'b111011001000;
   43329: result <= 12'b111011001001;
   43330: result <= 12'b111011001001;
   43331: result <= 12'b111011001001;
   43332: result <= 12'b111011001001;
   43333: result <= 12'b111011001001;
   43334: result <= 12'b111011001001;
   43335: result <= 12'b111011001001;
   43336: result <= 12'b111011001001;
   43337: result <= 12'b111011001001;
   43338: result <= 12'b111011001001;
   43339: result <= 12'b111011001010;
   43340: result <= 12'b111011001010;
   43341: result <= 12'b111011001010;
   43342: result <= 12'b111011001010;
   43343: result <= 12'b111011001010;
   43344: result <= 12'b111011001010;
   43345: result <= 12'b111011001010;
   43346: result <= 12'b111011001010;
   43347: result <= 12'b111011001010;
   43348: result <= 12'b111011001011;
   43349: result <= 12'b111011001011;
   43350: result <= 12'b111011001011;
   43351: result <= 12'b111011001011;
   43352: result <= 12'b111011001011;
   43353: result <= 12'b111011001011;
   43354: result <= 12'b111011001011;
   43355: result <= 12'b111011001011;
   43356: result <= 12'b111011001011;
   43357: result <= 12'b111011001011;
   43358: result <= 12'b111011001100;
   43359: result <= 12'b111011001100;
   43360: result <= 12'b111011001100;
   43361: result <= 12'b111011001100;
   43362: result <= 12'b111011001100;
   43363: result <= 12'b111011001100;
   43364: result <= 12'b111011001100;
   43365: result <= 12'b111011001100;
   43366: result <= 12'b111011001100;
   43367: result <= 12'b111011001100;
   43368: result <= 12'b111011001101;
   43369: result <= 12'b111011001101;
   43370: result <= 12'b111011001101;
   43371: result <= 12'b111011001101;
   43372: result <= 12'b111011001101;
   43373: result <= 12'b111011001101;
   43374: result <= 12'b111011001101;
   43375: result <= 12'b111011001101;
   43376: result <= 12'b111011001101;
   43377: result <= 12'b111011001110;
   43378: result <= 12'b111011001110;
   43379: result <= 12'b111011001110;
   43380: result <= 12'b111011001110;
   43381: result <= 12'b111011001110;
   43382: result <= 12'b111011001110;
   43383: result <= 12'b111011001110;
   43384: result <= 12'b111011001110;
   43385: result <= 12'b111011001110;
   43386: result <= 12'b111011001110;
   43387: result <= 12'b111011001111;
   43388: result <= 12'b111011001111;
   43389: result <= 12'b111011001111;
   43390: result <= 12'b111011001111;
   43391: result <= 12'b111011001111;
   43392: result <= 12'b111011001111;
   43393: result <= 12'b111011001111;
   43394: result <= 12'b111011001111;
   43395: result <= 12'b111011001111;
   43396: result <= 12'b111011001111;
   43397: result <= 12'b111011010000;
   43398: result <= 12'b111011010000;
   43399: result <= 12'b111011010000;
   43400: result <= 12'b111011010000;
   43401: result <= 12'b111011010000;
   43402: result <= 12'b111011010000;
   43403: result <= 12'b111011010000;
   43404: result <= 12'b111011010000;
   43405: result <= 12'b111011010000;
   43406: result <= 12'b111011010001;
   43407: result <= 12'b111011010001;
   43408: result <= 12'b111011010001;
   43409: result <= 12'b111011010001;
   43410: result <= 12'b111011010001;
   43411: result <= 12'b111011010001;
   43412: result <= 12'b111011010001;
   43413: result <= 12'b111011010001;
   43414: result <= 12'b111011010001;
   43415: result <= 12'b111011010001;
   43416: result <= 12'b111011010010;
   43417: result <= 12'b111011010010;
   43418: result <= 12'b111011010010;
   43419: result <= 12'b111011010010;
   43420: result <= 12'b111011010010;
   43421: result <= 12'b111011010010;
   43422: result <= 12'b111011010010;
   43423: result <= 12'b111011010010;
   43424: result <= 12'b111011010010;
   43425: result <= 12'b111011010010;
   43426: result <= 12'b111011010011;
   43427: result <= 12'b111011010011;
   43428: result <= 12'b111011010011;
   43429: result <= 12'b111011010011;
   43430: result <= 12'b111011010011;
   43431: result <= 12'b111011010011;
   43432: result <= 12'b111011010011;
   43433: result <= 12'b111011010011;
   43434: result <= 12'b111011010011;
   43435: result <= 12'b111011010011;
   43436: result <= 12'b111011010100;
   43437: result <= 12'b111011010100;
   43438: result <= 12'b111011010100;
   43439: result <= 12'b111011010100;
   43440: result <= 12'b111011010100;
   43441: result <= 12'b111011010100;
   43442: result <= 12'b111011010100;
   43443: result <= 12'b111011010100;
   43444: result <= 12'b111011010100;
   43445: result <= 12'b111011010101;
   43446: result <= 12'b111011010101;
   43447: result <= 12'b111011010101;
   43448: result <= 12'b111011010101;
   43449: result <= 12'b111011010101;
   43450: result <= 12'b111011010101;
   43451: result <= 12'b111011010101;
   43452: result <= 12'b111011010101;
   43453: result <= 12'b111011010101;
   43454: result <= 12'b111011010101;
   43455: result <= 12'b111011010110;
   43456: result <= 12'b111011010110;
   43457: result <= 12'b111011010110;
   43458: result <= 12'b111011010110;
   43459: result <= 12'b111011010110;
   43460: result <= 12'b111011010110;
   43461: result <= 12'b111011010110;
   43462: result <= 12'b111011010110;
   43463: result <= 12'b111011010110;
   43464: result <= 12'b111011010110;
   43465: result <= 12'b111011010111;
   43466: result <= 12'b111011010111;
   43467: result <= 12'b111011010111;
   43468: result <= 12'b111011010111;
   43469: result <= 12'b111011010111;
   43470: result <= 12'b111011010111;
   43471: result <= 12'b111011010111;
   43472: result <= 12'b111011010111;
   43473: result <= 12'b111011010111;
   43474: result <= 12'b111011010111;
   43475: result <= 12'b111011011000;
   43476: result <= 12'b111011011000;
   43477: result <= 12'b111011011000;
   43478: result <= 12'b111011011000;
   43479: result <= 12'b111011011000;
   43480: result <= 12'b111011011000;
   43481: result <= 12'b111011011000;
   43482: result <= 12'b111011011000;
   43483: result <= 12'b111011011000;
   43484: result <= 12'b111011011000;
   43485: result <= 12'b111011011001;
   43486: result <= 12'b111011011001;
   43487: result <= 12'b111011011001;
   43488: result <= 12'b111011011001;
   43489: result <= 12'b111011011001;
   43490: result <= 12'b111011011001;
   43491: result <= 12'b111011011001;
   43492: result <= 12'b111011011001;
   43493: result <= 12'b111011011001;
   43494: result <= 12'b111011011001;
   43495: result <= 12'b111011011010;
   43496: result <= 12'b111011011010;
   43497: result <= 12'b111011011010;
   43498: result <= 12'b111011011010;
   43499: result <= 12'b111011011010;
   43500: result <= 12'b111011011010;
   43501: result <= 12'b111011011010;
   43502: result <= 12'b111011011010;
   43503: result <= 12'b111011011010;
   43504: result <= 12'b111011011011;
   43505: result <= 12'b111011011011;
   43506: result <= 12'b111011011011;
   43507: result <= 12'b111011011011;
   43508: result <= 12'b111011011011;
   43509: result <= 12'b111011011011;
   43510: result <= 12'b111011011011;
   43511: result <= 12'b111011011011;
   43512: result <= 12'b111011011011;
   43513: result <= 12'b111011011011;
   43514: result <= 12'b111011011100;
   43515: result <= 12'b111011011100;
   43516: result <= 12'b111011011100;
   43517: result <= 12'b111011011100;
   43518: result <= 12'b111011011100;
   43519: result <= 12'b111011011100;
   43520: result <= 12'b111011011100;
   43521: result <= 12'b111011011100;
   43522: result <= 12'b111011011100;
   43523: result <= 12'b111011011100;
   43524: result <= 12'b111011011101;
   43525: result <= 12'b111011011101;
   43526: result <= 12'b111011011101;
   43527: result <= 12'b111011011101;
   43528: result <= 12'b111011011101;
   43529: result <= 12'b111011011101;
   43530: result <= 12'b111011011101;
   43531: result <= 12'b111011011101;
   43532: result <= 12'b111011011101;
   43533: result <= 12'b111011011101;
   43534: result <= 12'b111011011110;
   43535: result <= 12'b111011011110;
   43536: result <= 12'b111011011110;
   43537: result <= 12'b111011011110;
   43538: result <= 12'b111011011110;
   43539: result <= 12'b111011011110;
   43540: result <= 12'b111011011110;
   43541: result <= 12'b111011011110;
   43542: result <= 12'b111011011110;
   43543: result <= 12'b111011011110;
   43544: result <= 12'b111011011111;
   43545: result <= 12'b111011011111;
   43546: result <= 12'b111011011111;
   43547: result <= 12'b111011011111;
   43548: result <= 12'b111011011111;
   43549: result <= 12'b111011011111;
   43550: result <= 12'b111011011111;
   43551: result <= 12'b111011011111;
   43552: result <= 12'b111011011111;
   43553: result <= 12'b111011011111;
   43554: result <= 12'b111011100000;
   43555: result <= 12'b111011100000;
   43556: result <= 12'b111011100000;
   43557: result <= 12'b111011100000;
   43558: result <= 12'b111011100000;
   43559: result <= 12'b111011100000;
   43560: result <= 12'b111011100000;
   43561: result <= 12'b111011100000;
   43562: result <= 12'b111011100000;
   43563: result <= 12'b111011100000;
   43564: result <= 12'b111011100001;
   43565: result <= 12'b111011100001;
   43566: result <= 12'b111011100001;
   43567: result <= 12'b111011100001;
   43568: result <= 12'b111011100001;
   43569: result <= 12'b111011100001;
   43570: result <= 12'b111011100001;
   43571: result <= 12'b111011100001;
   43572: result <= 12'b111011100001;
   43573: result <= 12'b111011100001;
   43574: result <= 12'b111011100010;
   43575: result <= 12'b111011100010;
   43576: result <= 12'b111011100010;
   43577: result <= 12'b111011100010;
   43578: result <= 12'b111011100010;
   43579: result <= 12'b111011100010;
   43580: result <= 12'b111011100010;
   43581: result <= 12'b111011100010;
   43582: result <= 12'b111011100010;
   43583: result <= 12'b111011100010;
   43584: result <= 12'b111011100011;
   43585: result <= 12'b111011100011;
   43586: result <= 12'b111011100011;
   43587: result <= 12'b111011100011;
   43588: result <= 12'b111011100011;
   43589: result <= 12'b111011100011;
   43590: result <= 12'b111011100011;
   43591: result <= 12'b111011100011;
   43592: result <= 12'b111011100011;
   43593: result <= 12'b111011100011;
   43594: result <= 12'b111011100100;
   43595: result <= 12'b111011100100;
   43596: result <= 12'b111011100100;
   43597: result <= 12'b111011100100;
   43598: result <= 12'b111011100100;
   43599: result <= 12'b111011100100;
   43600: result <= 12'b111011100100;
   43601: result <= 12'b111011100100;
   43602: result <= 12'b111011100100;
   43603: result <= 12'b111011100100;
   43604: result <= 12'b111011100101;
   43605: result <= 12'b111011100101;
   43606: result <= 12'b111011100101;
   43607: result <= 12'b111011100101;
   43608: result <= 12'b111011100101;
   43609: result <= 12'b111011100101;
   43610: result <= 12'b111011100101;
   43611: result <= 12'b111011100101;
   43612: result <= 12'b111011100101;
   43613: result <= 12'b111011100101;
   43614: result <= 12'b111011100110;
   43615: result <= 12'b111011100110;
   43616: result <= 12'b111011100110;
   43617: result <= 12'b111011100110;
   43618: result <= 12'b111011100110;
   43619: result <= 12'b111011100110;
   43620: result <= 12'b111011100110;
   43621: result <= 12'b111011100110;
   43622: result <= 12'b111011100110;
   43623: result <= 12'b111011100110;
   43624: result <= 12'b111011100111;
   43625: result <= 12'b111011100111;
   43626: result <= 12'b111011100111;
   43627: result <= 12'b111011100111;
   43628: result <= 12'b111011100111;
   43629: result <= 12'b111011100111;
   43630: result <= 12'b111011100111;
   43631: result <= 12'b111011100111;
   43632: result <= 12'b111011100111;
   43633: result <= 12'b111011100111;
   43634: result <= 12'b111011101000;
   43635: result <= 12'b111011101000;
   43636: result <= 12'b111011101000;
   43637: result <= 12'b111011101000;
   43638: result <= 12'b111011101000;
   43639: result <= 12'b111011101000;
   43640: result <= 12'b111011101000;
   43641: result <= 12'b111011101000;
   43642: result <= 12'b111011101000;
   43643: result <= 12'b111011101000;
   43644: result <= 12'b111011101001;
   43645: result <= 12'b111011101001;
   43646: result <= 12'b111011101001;
   43647: result <= 12'b111011101001;
   43648: result <= 12'b111011101001;
   43649: result <= 12'b111011101001;
   43650: result <= 12'b111011101001;
   43651: result <= 12'b111011101001;
   43652: result <= 12'b111011101001;
   43653: result <= 12'b111011101001;
   43654: result <= 12'b111011101010;
   43655: result <= 12'b111011101010;
   43656: result <= 12'b111011101010;
   43657: result <= 12'b111011101010;
   43658: result <= 12'b111011101010;
   43659: result <= 12'b111011101010;
   43660: result <= 12'b111011101010;
   43661: result <= 12'b111011101010;
   43662: result <= 12'b111011101010;
   43663: result <= 12'b111011101010;
   43664: result <= 12'b111011101010;
   43665: result <= 12'b111011101011;
   43666: result <= 12'b111011101011;
   43667: result <= 12'b111011101011;
   43668: result <= 12'b111011101011;
   43669: result <= 12'b111011101011;
   43670: result <= 12'b111011101011;
   43671: result <= 12'b111011101011;
   43672: result <= 12'b111011101011;
   43673: result <= 12'b111011101011;
   43674: result <= 12'b111011101011;
   43675: result <= 12'b111011101100;
   43676: result <= 12'b111011101100;
   43677: result <= 12'b111011101100;
   43678: result <= 12'b111011101100;
   43679: result <= 12'b111011101100;
   43680: result <= 12'b111011101100;
   43681: result <= 12'b111011101100;
   43682: result <= 12'b111011101100;
   43683: result <= 12'b111011101100;
   43684: result <= 12'b111011101100;
   43685: result <= 12'b111011101101;
   43686: result <= 12'b111011101101;
   43687: result <= 12'b111011101101;
   43688: result <= 12'b111011101101;
   43689: result <= 12'b111011101101;
   43690: result <= 12'b111011101101;
   43691: result <= 12'b111011101101;
   43692: result <= 12'b111011101101;
   43693: result <= 12'b111011101101;
   43694: result <= 12'b111011101101;
   43695: result <= 12'b111011101110;
   43696: result <= 12'b111011101110;
   43697: result <= 12'b111011101110;
   43698: result <= 12'b111011101110;
   43699: result <= 12'b111011101110;
   43700: result <= 12'b111011101110;
   43701: result <= 12'b111011101110;
   43702: result <= 12'b111011101110;
   43703: result <= 12'b111011101110;
   43704: result <= 12'b111011101110;
   43705: result <= 12'b111011101111;
   43706: result <= 12'b111011101111;
   43707: result <= 12'b111011101111;
   43708: result <= 12'b111011101111;
   43709: result <= 12'b111011101111;
   43710: result <= 12'b111011101111;
   43711: result <= 12'b111011101111;
   43712: result <= 12'b111011101111;
   43713: result <= 12'b111011101111;
   43714: result <= 12'b111011101111;
   43715: result <= 12'b111011110000;
   43716: result <= 12'b111011110000;
   43717: result <= 12'b111011110000;
   43718: result <= 12'b111011110000;
   43719: result <= 12'b111011110000;
   43720: result <= 12'b111011110000;
   43721: result <= 12'b111011110000;
   43722: result <= 12'b111011110000;
   43723: result <= 12'b111011110000;
   43724: result <= 12'b111011110000;
   43725: result <= 12'b111011110000;
   43726: result <= 12'b111011110001;
   43727: result <= 12'b111011110001;
   43728: result <= 12'b111011110001;
   43729: result <= 12'b111011110001;
   43730: result <= 12'b111011110001;
   43731: result <= 12'b111011110001;
   43732: result <= 12'b111011110001;
   43733: result <= 12'b111011110001;
   43734: result <= 12'b111011110001;
   43735: result <= 12'b111011110001;
   43736: result <= 12'b111011110010;
   43737: result <= 12'b111011110010;
   43738: result <= 12'b111011110010;
   43739: result <= 12'b111011110010;
   43740: result <= 12'b111011110010;
   43741: result <= 12'b111011110010;
   43742: result <= 12'b111011110010;
   43743: result <= 12'b111011110010;
   43744: result <= 12'b111011110010;
   43745: result <= 12'b111011110010;
   43746: result <= 12'b111011110011;
   43747: result <= 12'b111011110011;
   43748: result <= 12'b111011110011;
   43749: result <= 12'b111011110011;
   43750: result <= 12'b111011110011;
   43751: result <= 12'b111011110011;
   43752: result <= 12'b111011110011;
   43753: result <= 12'b111011110011;
   43754: result <= 12'b111011110011;
   43755: result <= 12'b111011110011;
   43756: result <= 12'b111011110011;
   43757: result <= 12'b111011110100;
   43758: result <= 12'b111011110100;
   43759: result <= 12'b111011110100;
   43760: result <= 12'b111011110100;
   43761: result <= 12'b111011110100;
   43762: result <= 12'b111011110100;
   43763: result <= 12'b111011110100;
   43764: result <= 12'b111011110100;
   43765: result <= 12'b111011110100;
   43766: result <= 12'b111011110100;
   43767: result <= 12'b111011110101;
   43768: result <= 12'b111011110101;
   43769: result <= 12'b111011110101;
   43770: result <= 12'b111011110101;
   43771: result <= 12'b111011110101;
   43772: result <= 12'b111011110101;
   43773: result <= 12'b111011110101;
   43774: result <= 12'b111011110101;
   43775: result <= 12'b111011110101;
   43776: result <= 12'b111011110101;
   43777: result <= 12'b111011110110;
   43778: result <= 12'b111011110110;
   43779: result <= 12'b111011110110;
   43780: result <= 12'b111011110110;
   43781: result <= 12'b111011110110;
   43782: result <= 12'b111011110110;
   43783: result <= 12'b111011110110;
   43784: result <= 12'b111011110110;
   43785: result <= 12'b111011110110;
   43786: result <= 12'b111011110110;
   43787: result <= 12'b111011110111;
   43788: result <= 12'b111011110111;
   43789: result <= 12'b111011110111;
   43790: result <= 12'b111011110111;
   43791: result <= 12'b111011110111;
   43792: result <= 12'b111011110111;
   43793: result <= 12'b111011110111;
   43794: result <= 12'b111011110111;
   43795: result <= 12'b111011110111;
   43796: result <= 12'b111011110111;
   43797: result <= 12'b111011110111;
   43798: result <= 12'b111011111000;
   43799: result <= 12'b111011111000;
   43800: result <= 12'b111011111000;
   43801: result <= 12'b111011111000;
   43802: result <= 12'b111011111000;
   43803: result <= 12'b111011111000;
   43804: result <= 12'b111011111000;
   43805: result <= 12'b111011111000;
   43806: result <= 12'b111011111000;
   43807: result <= 12'b111011111000;
   43808: result <= 12'b111011111001;
   43809: result <= 12'b111011111001;
   43810: result <= 12'b111011111001;
   43811: result <= 12'b111011111001;
   43812: result <= 12'b111011111001;
   43813: result <= 12'b111011111001;
   43814: result <= 12'b111011111001;
   43815: result <= 12'b111011111001;
   43816: result <= 12'b111011111001;
   43817: result <= 12'b111011111001;
   43818: result <= 12'b111011111001;
   43819: result <= 12'b111011111010;
   43820: result <= 12'b111011111010;
   43821: result <= 12'b111011111010;
   43822: result <= 12'b111011111010;
   43823: result <= 12'b111011111010;
   43824: result <= 12'b111011111010;
   43825: result <= 12'b111011111010;
   43826: result <= 12'b111011111010;
   43827: result <= 12'b111011111010;
   43828: result <= 12'b111011111010;
   43829: result <= 12'b111011111011;
   43830: result <= 12'b111011111011;
   43831: result <= 12'b111011111011;
   43832: result <= 12'b111011111011;
   43833: result <= 12'b111011111011;
   43834: result <= 12'b111011111011;
   43835: result <= 12'b111011111011;
   43836: result <= 12'b111011111011;
   43837: result <= 12'b111011111011;
   43838: result <= 12'b111011111011;
   43839: result <= 12'b111011111100;
   43840: result <= 12'b111011111100;
   43841: result <= 12'b111011111100;
   43842: result <= 12'b111011111100;
   43843: result <= 12'b111011111100;
   43844: result <= 12'b111011111100;
   43845: result <= 12'b111011111100;
   43846: result <= 12'b111011111100;
   43847: result <= 12'b111011111100;
   43848: result <= 12'b111011111100;
   43849: result <= 12'b111011111100;
   43850: result <= 12'b111011111101;
   43851: result <= 12'b111011111101;
   43852: result <= 12'b111011111101;
   43853: result <= 12'b111011111101;
   43854: result <= 12'b111011111101;
   43855: result <= 12'b111011111101;
   43856: result <= 12'b111011111101;
   43857: result <= 12'b111011111101;
   43858: result <= 12'b111011111101;
   43859: result <= 12'b111011111101;
   43860: result <= 12'b111011111110;
   43861: result <= 12'b111011111110;
   43862: result <= 12'b111011111110;
   43863: result <= 12'b111011111110;
   43864: result <= 12'b111011111110;
   43865: result <= 12'b111011111110;
   43866: result <= 12'b111011111110;
   43867: result <= 12'b111011111110;
   43868: result <= 12'b111011111110;
   43869: result <= 12'b111011111110;
   43870: result <= 12'b111011111110;
   43871: result <= 12'b111011111111;
   43872: result <= 12'b111011111111;
   43873: result <= 12'b111011111111;
   43874: result <= 12'b111011111111;
   43875: result <= 12'b111011111111;
   43876: result <= 12'b111011111111;
   43877: result <= 12'b111011111111;
   43878: result <= 12'b111011111111;
   43879: result <= 12'b111011111111;
   43880: result <= 12'b111011111111;
   43881: result <= 12'b111100000000;
   43882: result <= 12'b111100000000;
   43883: result <= 12'b111100000000;
   43884: result <= 12'b111100000000;
   43885: result <= 12'b111100000000;
   43886: result <= 12'b111100000000;
   43887: result <= 12'b111100000000;
   43888: result <= 12'b111100000000;
   43889: result <= 12'b111100000000;
   43890: result <= 12'b111100000000;
   43891: result <= 12'b111100000000;
   43892: result <= 12'b111100000001;
   43893: result <= 12'b111100000001;
   43894: result <= 12'b111100000001;
   43895: result <= 12'b111100000001;
   43896: result <= 12'b111100000001;
   43897: result <= 12'b111100000001;
   43898: result <= 12'b111100000001;
   43899: result <= 12'b111100000001;
   43900: result <= 12'b111100000001;
   43901: result <= 12'b111100000001;
   43902: result <= 12'b111100000010;
   43903: result <= 12'b111100000010;
   43904: result <= 12'b111100000010;
   43905: result <= 12'b111100000010;
   43906: result <= 12'b111100000010;
   43907: result <= 12'b111100000010;
   43908: result <= 12'b111100000010;
   43909: result <= 12'b111100000010;
   43910: result <= 12'b111100000010;
   43911: result <= 12'b111100000010;
   43912: result <= 12'b111100000010;
   43913: result <= 12'b111100000011;
   43914: result <= 12'b111100000011;
   43915: result <= 12'b111100000011;
   43916: result <= 12'b111100000011;
   43917: result <= 12'b111100000011;
   43918: result <= 12'b111100000011;
   43919: result <= 12'b111100000011;
   43920: result <= 12'b111100000011;
   43921: result <= 12'b111100000011;
   43922: result <= 12'b111100000011;
   43923: result <= 12'b111100000011;
   43924: result <= 12'b111100000100;
   43925: result <= 12'b111100000100;
   43926: result <= 12'b111100000100;
   43927: result <= 12'b111100000100;
   43928: result <= 12'b111100000100;
   43929: result <= 12'b111100000100;
   43930: result <= 12'b111100000100;
   43931: result <= 12'b111100000100;
   43932: result <= 12'b111100000100;
   43933: result <= 12'b111100000100;
   43934: result <= 12'b111100000101;
   43935: result <= 12'b111100000101;
   43936: result <= 12'b111100000101;
   43937: result <= 12'b111100000101;
   43938: result <= 12'b111100000101;
   43939: result <= 12'b111100000101;
   43940: result <= 12'b111100000101;
   43941: result <= 12'b111100000101;
   43942: result <= 12'b111100000101;
   43943: result <= 12'b111100000101;
   43944: result <= 12'b111100000101;
   43945: result <= 12'b111100000110;
   43946: result <= 12'b111100000110;
   43947: result <= 12'b111100000110;
   43948: result <= 12'b111100000110;
   43949: result <= 12'b111100000110;
   43950: result <= 12'b111100000110;
   43951: result <= 12'b111100000110;
   43952: result <= 12'b111100000110;
   43953: result <= 12'b111100000110;
   43954: result <= 12'b111100000110;
   43955: result <= 12'b111100000110;
   43956: result <= 12'b111100000111;
   43957: result <= 12'b111100000111;
   43958: result <= 12'b111100000111;
   43959: result <= 12'b111100000111;
   43960: result <= 12'b111100000111;
   43961: result <= 12'b111100000111;
   43962: result <= 12'b111100000111;
   43963: result <= 12'b111100000111;
   43964: result <= 12'b111100000111;
   43965: result <= 12'b111100000111;
   43966: result <= 12'b111100001000;
   43967: result <= 12'b111100001000;
   43968: result <= 12'b111100001000;
   43969: result <= 12'b111100001000;
   43970: result <= 12'b111100001000;
   43971: result <= 12'b111100001000;
   43972: result <= 12'b111100001000;
   43973: result <= 12'b111100001000;
   43974: result <= 12'b111100001000;
   43975: result <= 12'b111100001000;
   43976: result <= 12'b111100001000;
   43977: result <= 12'b111100001001;
   43978: result <= 12'b111100001001;
   43979: result <= 12'b111100001001;
   43980: result <= 12'b111100001001;
   43981: result <= 12'b111100001001;
   43982: result <= 12'b111100001001;
   43983: result <= 12'b111100001001;
   43984: result <= 12'b111100001001;
   43985: result <= 12'b111100001001;
   43986: result <= 12'b111100001001;
   43987: result <= 12'b111100001001;
   43988: result <= 12'b111100001010;
   43989: result <= 12'b111100001010;
   43990: result <= 12'b111100001010;
   43991: result <= 12'b111100001010;
   43992: result <= 12'b111100001010;
   43993: result <= 12'b111100001010;
   43994: result <= 12'b111100001010;
   43995: result <= 12'b111100001010;
   43996: result <= 12'b111100001010;
   43997: result <= 12'b111100001010;
   43998: result <= 12'b111100001011;
   43999: result <= 12'b111100001011;
   44000: result <= 12'b111100001011;
   44001: result <= 12'b111100001011;
   44002: result <= 12'b111100001011;
   44003: result <= 12'b111100001011;
   44004: result <= 12'b111100001011;
   44005: result <= 12'b111100001011;
   44006: result <= 12'b111100001011;
   44007: result <= 12'b111100001011;
   44008: result <= 12'b111100001011;
   44009: result <= 12'b111100001100;
   44010: result <= 12'b111100001100;
   44011: result <= 12'b111100001100;
   44012: result <= 12'b111100001100;
   44013: result <= 12'b111100001100;
   44014: result <= 12'b111100001100;
   44015: result <= 12'b111100001100;
   44016: result <= 12'b111100001100;
   44017: result <= 12'b111100001100;
   44018: result <= 12'b111100001100;
   44019: result <= 12'b111100001100;
   44020: result <= 12'b111100001101;
   44021: result <= 12'b111100001101;
   44022: result <= 12'b111100001101;
   44023: result <= 12'b111100001101;
   44024: result <= 12'b111100001101;
   44025: result <= 12'b111100001101;
   44026: result <= 12'b111100001101;
   44027: result <= 12'b111100001101;
   44028: result <= 12'b111100001101;
   44029: result <= 12'b111100001101;
   44030: result <= 12'b111100001101;
   44031: result <= 12'b111100001110;
   44032: result <= 12'b111100001110;
   44033: result <= 12'b111100001110;
   44034: result <= 12'b111100001110;
   44035: result <= 12'b111100001110;
   44036: result <= 12'b111100001110;
   44037: result <= 12'b111100001110;
   44038: result <= 12'b111100001110;
   44039: result <= 12'b111100001110;
   44040: result <= 12'b111100001110;
   44041: result <= 12'b111100001111;
   44042: result <= 12'b111100001111;
   44043: result <= 12'b111100001111;
   44044: result <= 12'b111100001111;
   44045: result <= 12'b111100001111;
   44046: result <= 12'b111100001111;
   44047: result <= 12'b111100001111;
   44048: result <= 12'b111100001111;
   44049: result <= 12'b111100001111;
   44050: result <= 12'b111100001111;
   44051: result <= 12'b111100001111;
   44052: result <= 12'b111100010000;
   44053: result <= 12'b111100010000;
   44054: result <= 12'b111100010000;
   44055: result <= 12'b111100010000;
   44056: result <= 12'b111100010000;
   44057: result <= 12'b111100010000;
   44058: result <= 12'b111100010000;
   44059: result <= 12'b111100010000;
   44060: result <= 12'b111100010000;
   44061: result <= 12'b111100010000;
   44062: result <= 12'b111100010000;
   44063: result <= 12'b111100010001;
   44064: result <= 12'b111100010001;
   44065: result <= 12'b111100010001;
   44066: result <= 12'b111100010001;
   44067: result <= 12'b111100010001;
   44068: result <= 12'b111100010001;
   44069: result <= 12'b111100010001;
   44070: result <= 12'b111100010001;
   44071: result <= 12'b111100010001;
   44072: result <= 12'b111100010001;
   44073: result <= 12'b111100010001;
   44074: result <= 12'b111100010010;
   44075: result <= 12'b111100010010;
   44076: result <= 12'b111100010010;
   44077: result <= 12'b111100010010;
   44078: result <= 12'b111100010010;
   44079: result <= 12'b111100010010;
   44080: result <= 12'b111100010010;
   44081: result <= 12'b111100010010;
   44082: result <= 12'b111100010010;
   44083: result <= 12'b111100010010;
   44084: result <= 12'b111100010010;
   44085: result <= 12'b111100010011;
   44086: result <= 12'b111100010011;
   44087: result <= 12'b111100010011;
   44088: result <= 12'b111100010011;
   44089: result <= 12'b111100010011;
   44090: result <= 12'b111100010011;
   44091: result <= 12'b111100010011;
   44092: result <= 12'b111100010011;
   44093: result <= 12'b111100010011;
   44094: result <= 12'b111100010011;
   44095: result <= 12'b111100010011;
   44096: result <= 12'b111100010100;
   44097: result <= 12'b111100010100;
   44098: result <= 12'b111100010100;
   44099: result <= 12'b111100010100;
   44100: result <= 12'b111100010100;
   44101: result <= 12'b111100010100;
   44102: result <= 12'b111100010100;
   44103: result <= 12'b111100010100;
   44104: result <= 12'b111100010100;
   44105: result <= 12'b111100010100;
   44106: result <= 12'b111100010100;
   44107: result <= 12'b111100010101;
   44108: result <= 12'b111100010101;
   44109: result <= 12'b111100010101;
   44110: result <= 12'b111100010101;
   44111: result <= 12'b111100010101;
   44112: result <= 12'b111100010101;
   44113: result <= 12'b111100010101;
   44114: result <= 12'b111100010101;
   44115: result <= 12'b111100010101;
   44116: result <= 12'b111100010101;
   44117: result <= 12'b111100010101;
   44118: result <= 12'b111100010110;
   44119: result <= 12'b111100010110;
   44120: result <= 12'b111100010110;
   44121: result <= 12'b111100010110;
   44122: result <= 12'b111100010110;
   44123: result <= 12'b111100010110;
   44124: result <= 12'b111100010110;
   44125: result <= 12'b111100010110;
   44126: result <= 12'b111100010110;
   44127: result <= 12'b111100010110;
   44128: result <= 12'b111100010110;
   44129: result <= 12'b111100010111;
   44130: result <= 12'b111100010111;
   44131: result <= 12'b111100010111;
   44132: result <= 12'b111100010111;
   44133: result <= 12'b111100010111;
   44134: result <= 12'b111100010111;
   44135: result <= 12'b111100010111;
   44136: result <= 12'b111100010111;
   44137: result <= 12'b111100010111;
   44138: result <= 12'b111100010111;
   44139: result <= 12'b111100010111;
   44140: result <= 12'b111100011000;
   44141: result <= 12'b111100011000;
   44142: result <= 12'b111100011000;
   44143: result <= 12'b111100011000;
   44144: result <= 12'b111100011000;
   44145: result <= 12'b111100011000;
   44146: result <= 12'b111100011000;
   44147: result <= 12'b111100011000;
   44148: result <= 12'b111100011000;
   44149: result <= 12'b111100011000;
   44150: result <= 12'b111100011000;
   44151: result <= 12'b111100011001;
   44152: result <= 12'b111100011001;
   44153: result <= 12'b111100011001;
   44154: result <= 12'b111100011001;
   44155: result <= 12'b111100011001;
   44156: result <= 12'b111100011001;
   44157: result <= 12'b111100011001;
   44158: result <= 12'b111100011001;
   44159: result <= 12'b111100011001;
   44160: result <= 12'b111100011001;
   44161: result <= 12'b111100011001;
   44162: result <= 12'b111100011010;
   44163: result <= 12'b111100011010;
   44164: result <= 12'b111100011010;
   44165: result <= 12'b111100011010;
   44166: result <= 12'b111100011010;
   44167: result <= 12'b111100011010;
   44168: result <= 12'b111100011010;
   44169: result <= 12'b111100011010;
   44170: result <= 12'b111100011010;
   44171: result <= 12'b111100011010;
   44172: result <= 12'b111100011010;
   44173: result <= 12'b111100011011;
   44174: result <= 12'b111100011011;
   44175: result <= 12'b111100011011;
   44176: result <= 12'b111100011011;
   44177: result <= 12'b111100011011;
   44178: result <= 12'b111100011011;
   44179: result <= 12'b111100011011;
   44180: result <= 12'b111100011011;
   44181: result <= 12'b111100011011;
   44182: result <= 12'b111100011011;
   44183: result <= 12'b111100011011;
   44184: result <= 12'b111100011100;
   44185: result <= 12'b111100011100;
   44186: result <= 12'b111100011100;
   44187: result <= 12'b111100011100;
   44188: result <= 12'b111100011100;
   44189: result <= 12'b111100011100;
   44190: result <= 12'b111100011100;
   44191: result <= 12'b111100011100;
   44192: result <= 12'b111100011100;
   44193: result <= 12'b111100011100;
   44194: result <= 12'b111100011100;
   44195: result <= 12'b111100011101;
   44196: result <= 12'b111100011101;
   44197: result <= 12'b111100011101;
   44198: result <= 12'b111100011101;
   44199: result <= 12'b111100011101;
   44200: result <= 12'b111100011101;
   44201: result <= 12'b111100011101;
   44202: result <= 12'b111100011101;
   44203: result <= 12'b111100011101;
   44204: result <= 12'b111100011101;
   44205: result <= 12'b111100011101;
   44206: result <= 12'b111100011110;
   44207: result <= 12'b111100011110;
   44208: result <= 12'b111100011110;
   44209: result <= 12'b111100011110;
   44210: result <= 12'b111100011110;
   44211: result <= 12'b111100011110;
   44212: result <= 12'b111100011110;
   44213: result <= 12'b111100011110;
   44214: result <= 12'b111100011110;
   44215: result <= 12'b111100011110;
   44216: result <= 12'b111100011110;
   44217: result <= 12'b111100011111;
   44218: result <= 12'b111100011111;
   44219: result <= 12'b111100011111;
   44220: result <= 12'b111100011111;
   44221: result <= 12'b111100011111;
   44222: result <= 12'b111100011111;
   44223: result <= 12'b111100011111;
   44224: result <= 12'b111100011111;
   44225: result <= 12'b111100011111;
   44226: result <= 12'b111100011111;
   44227: result <= 12'b111100011111;
   44228: result <= 12'b111100011111;
   44229: result <= 12'b111100100000;
   44230: result <= 12'b111100100000;
   44231: result <= 12'b111100100000;
   44232: result <= 12'b111100100000;
   44233: result <= 12'b111100100000;
   44234: result <= 12'b111100100000;
   44235: result <= 12'b111100100000;
   44236: result <= 12'b111100100000;
   44237: result <= 12'b111100100000;
   44238: result <= 12'b111100100000;
   44239: result <= 12'b111100100000;
   44240: result <= 12'b111100100001;
   44241: result <= 12'b111100100001;
   44242: result <= 12'b111100100001;
   44243: result <= 12'b111100100001;
   44244: result <= 12'b111100100001;
   44245: result <= 12'b111100100001;
   44246: result <= 12'b111100100001;
   44247: result <= 12'b111100100001;
   44248: result <= 12'b111100100001;
   44249: result <= 12'b111100100001;
   44250: result <= 12'b111100100001;
   44251: result <= 12'b111100100010;
   44252: result <= 12'b111100100010;
   44253: result <= 12'b111100100010;
   44254: result <= 12'b111100100010;
   44255: result <= 12'b111100100010;
   44256: result <= 12'b111100100010;
   44257: result <= 12'b111100100010;
   44258: result <= 12'b111100100010;
   44259: result <= 12'b111100100010;
   44260: result <= 12'b111100100010;
   44261: result <= 12'b111100100010;
   44262: result <= 12'b111100100011;
   44263: result <= 12'b111100100011;
   44264: result <= 12'b111100100011;
   44265: result <= 12'b111100100011;
   44266: result <= 12'b111100100011;
   44267: result <= 12'b111100100011;
   44268: result <= 12'b111100100011;
   44269: result <= 12'b111100100011;
   44270: result <= 12'b111100100011;
   44271: result <= 12'b111100100011;
   44272: result <= 12'b111100100011;
   44273: result <= 12'b111100100011;
   44274: result <= 12'b111100100100;
   44275: result <= 12'b111100100100;
   44276: result <= 12'b111100100100;
   44277: result <= 12'b111100100100;
   44278: result <= 12'b111100100100;
   44279: result <= 12'b111100100100;
   44280: result <= 12'b111100100100;
   44281: result <= 12'b111100100100;
   44282: result <= 12'b111100100100;
   44283: result <= 12'b111100100100;
   44284: result <= 12'b111100100100;
   44285: result <= 12'b111100100101;
   44286: result <= 12'b111100100101;
   44287: result <= 12'b111100100101;
   44288: result <= 12'b111100100101;
   44289: result <= 12'b111100100101;
   44290: result <= 12'b111100100101;
   44291: result <= 12'b111100100101;
   44292: result <= 12'b111100100101;
   44293: result <= 12'b111100100101;
   44294: result <= 12'b111100100101;
   44295: result <= 12'b111100100101;
   44296: result <= 12'b111100100110;
   44297: result <= 12'b111100100110;
   44298: result <= 12'b111100100110;
   44299: result <= 12'b111100100110;
   44300: result <= 12'b111100100110;
   44301: result <= 12'b111100100110;
   44302: result <= 12'b111100100110;
   44303: result <= 12'b111100100110;
   44304: result <= 12'b111100100110;
   44305: result <= 12'b111100100110;
   44306: result <= 12'b111100100110;
   44307: result <= 12'b111100100110;
   44308: result <= 12'b111100100111;
   44309: result <= 12'b111100100111;
   44310: result <= 12'b111100100111;
   44311: result <= 12'b111100100111;
   44312: result <= 12'b111100100111;
   44313: result <= 12'b111100100111;
   44314: result <= 12'b111100100111;
   44315: result <= 12'b111100100111;
   44316: result <= 12'b111100100111;
   44317: result <= 12'b111100100111;
   44318: result <= 12'b111100100111;
   44319: result <= 12'b111100101000;
   44320: result <= 12'b111100101000;
   44321: result <= 12'b111100101000;
   44322: result <= 12'b111100101000;
   44323: result <= 12'b111100101000;
   44324: result <= 12'b111100101000;
   44325: result <= 12'b111100101000;
   44326: result <= 12'b111100101000;
   44327: result <= 12'b111100101000;
   44328: result <= 12'b111100101000;
   44329: result <= 12'b111100101000;
   44330: result <= 12'b111100101001;
   44331: result <= 12'b111100101001;
   44332: result <= 12'b111100101001;
   44333: result <= 12'b111100101001;
   44334: result <= 12'b111100101001;
   44335: result <= 12'b111100101001;
   44336: result <= 12'b111100101001;
   44337: result <= 12'b111100101001;
   44338: result <= 12'b111100101001;
   44339: result <= 12'b111100101001;
   44340: result <= 12'b111100101001;
   44341: result <= 12'b111100101001;
   44342: result <= 12'b111100101010;
   44343: result <= 12'b111100101010;
   44344: result <= 12'b111100101010;
   44345: result <= 12'b111100101010;
   44346: result <= 12'b111100101010;
   44347: result <= 12'b111100101010;
   44348: result <= 12'b111100101010;
   44349: result <= 12'b111100101010;
   44350: result <= 12'b111100101010;
   44351: result <= 12'b111100101010;
   44352: result <= 12'b111100101010;
   44353: result <= 12'b111100101011;
   44354: result <= 12'b111100101011;
   44355: result <= 12'b111100101011;
   44356: result <= 12'b111100101011;
   44357: result <= 12'b111100101011;
   44358: result <= 12'b111100101011;
   44359: result <= 12'b111100101011;
   44360: result <= 12'b111100101011;
   44361: result <= 12'b111100101011;
   44362: result <= 12'b111100101011;
   44363: result <= 12'b111100101011;
   44364: result <= 12'b111100101011;
   44365: result <= 12'b111100101100;
   44366: result <= 12'b111100101100;
   44367: result <= 12'b111100101100;
   44368: result <= 12'b111100101100;
   44369: result <= 12'b111100101100;
   44370: result <= 12'b111100101100;
   44371: result <= 12'b111100101100;
   44372: result <= 12'b111100101100;
   44373: result <= 12'b111100101100;
   44374: result <= 12'b111100101100;
   44375: result <= 12'b111100101100;
   44376: result <= 12'b111100101101;
   44377: result <= 12'b111100101101;
   44378: result <= 12'b111100101101;
   44379: result <= 12'b111100101101;
   44380: result <= 12'b111100101101;
   44381: result <= 12'b111100101101;
   44382: result <= 12'b111100101101;
   44383: result <= 12'b111100101101;
   44384: result <= 12'b111100101101;
   44385: result <= 12'b111100101101;
   44386: result <= 12'b111100101101;
   44387: result <= 12'b111100101101;
   44388: result <= 12'b111100101110;
   44389: result <= 12'b111100101110;
   44390: result <= 12'b111100101110;
   44391: result <= 12'b111100101110;
   44392: result <= 12'b111100101110;
   44393: result <= 12'b111100101110;
   44394: result <= 12'b111100101110;
   44395: result <= 12'b111100101110;
   44396: result <= 12'b111100101110;
   44397: result <= 12'b111100101110;
   44398: result <= 12'b111100101110;
   44399: result <= 12'b111100101111;
   44400: result <= 12'b111100101111;
   44401: result <= 12'b111100101111;
   44402: result <= 12'b111100101111;
   44403: result <= 12'b111100101111;
   44404: result <= 12'b111100101111;
   44405: result <= 12'b111100101111;
   44406: result <= 12'b111100101111;
   44407: result <= 12'b111100101111;
   44408: result <= 12'b111100101111;
   44409: result <= 12'b111100101111;
   44410: result <= 12'b111100101111;
   44411: result <= 12'b111100110000;
   44412: result <= 12'b111100110000;
   44413: result <= 12'b111100110000;
   44414: result <= 12'b111100110000;
   44415: result <= 12'b111100110000;
   44416: result <= 12'b111100110000;
   44417: result <= 12'b111100110000;
   44418: result <= 12'b111100110000;
   44419: result <= 12'b111100110000;
   44420: result <= 12'b111100110000;
   44421: result <= 12'b111100110000;
   44422: result <= 12'b111100110001;
   44423: result <= 12'b111100110001;
   44424: result <= 12'b111100110001;
   44425: result <= 12'b111100110001;
   44426: result <= 12'b111100110001;
   44427: result <= 12'b111100110001;
   44428: result <= 12'b111100110001;
   44429: result <= 12'b111100110001;
   44430: result <= 12'b111100110001;
   44431: result <= 12'b111100110001;
   44432: result <= 12'b111100110001;
   44433: result <= 12'b111100110001;
   44434: result <= 12'b111100110010;
   44435: result <= 12'b111100110010;
   44436: result <= 12'b111100110010;
   44437: result <= 12'b111100110010;
   44438: result <= 12'b111100110010;
   44439: result <= 12'b111100110010;
   44440: result <= 12'b111100110010;
   44441: result <= 12'b111100110010;
   44442: result <= 12'b111100110010;
   44443: result <= 12'b111100110010;
   44444: result <= 12'b111100110010;
   44445: result <= 12'b111100110010;
   44446: result <= 12'b111100110011;
   44447: result <= 12'b111100110011;
   44448: result <= 12'b111100110011;
   44449: result <= 12'b111100110011;
   44450: result <= 12'b111100110011;
   44451: result <= 12'b111100110011;
   44452: result <= 12'b111100110011;
   44453: result <= 12'b111100110011;
   44454: result <= 12'b111100110011;
   44455: result <= 12'b111100110011;
   44456: result <= 12'b111100110011;
   44457: result <= 12'b111100110100;
   44458: result <= 12'b111100110100;
   44459: result <= 12'b111100110100;
   44460: result <= 12'b111100110100;
   44461: result <= 12'b111100110100;
   44462: result <= 12'b111100110100;
   44463: result <= 12'b111100110100;
   44464: result <= 12'b111100110100;
   44465: result <= 12'b111100110100;
   44466: result <= 12'b111100110100;
   44467: result <= 12'b111100110100;
   44468: result <= 12'b111100110100;
   44469: result <= 12'b111100110101;
   44470: result <= 12'b111100110101;
   44471: result <= 12'b111100110101;
   44472: result <= 12'b111100110101;
   44473: result <= 12'b111100110101;
   44474: result <= 12'b111100110101;
   44475: result <= 12'b111100110101;
   44476: result <= 12'b111100110101;
   44477: result <= 12'b111100110101;
   44478: result <= 12'b111100110101;
   44479: result <= 12'b111100110101;
   44480: result <= 12'b111100110101;
   44481: result <= 12'b111100110110;
   44482: result <= 12'b111100110110;
   44483: result <= 12'b111100110110;
   44484: result <= 12'b111100110110;
   44485: result <= 12'b111100110110;
   44486: result <= 12'b111100110110;
   44487: result <= 12'b111100110110;
   44488: result <= 12'b111100110110;
   44489: result <= 12'b111100110110;
   44490: result <= 12'b111100110110;
   44491: result <= 12'b111100110110;
   44492: result <= 12'b111100110110;
   44493: result <= 12'b111100110111;
   44494: result <= 12'b111100110111;
   44495: result <= 12'b111100110111;
   44496: result <= 12'b111100110111;
   44497: result <= 12'b111100110111;
   44498: result <= 12'b111100110111;
   44499: result <= 12'b111100110111;
   44500: result <= 12'b111100110111;
   44501: result <= 12'b111100110111;
   44502: result <= 12'b111100110111;
   44503: result <= 12'b111100110111;
   44504: result <= 12'b111100110111;
   44505: result <= 12'b111100111000;
   44506: result <= 12'b111100111000;
   44507: result <= 12'b111100111000;
   44508: result <= 12'b111100111000;
   44509: result <= 12'b111100111000;
   44510: result <= 12'b111100111000;
   44511: result <= 12'b111100111000;
   44512: result <= 12'b111100111000;
   44513: result <= 12'b111100111000;
   44514: result <= 12'b111100111000;
   44515: result <= 12'b111100111000;
   44516: result <= 12'b111100111001;
   44517: result <= 12'b111100111001;
   44518: result <= 12'b111100111001;
   44519: result <= 12'b111100111001;
   44520: result <= 12'b111100111001;
   44521: result <= 12'b111100111001;
   44522: result <= 12'b111100111001;
   44523: result <= 12'b111100111001;
   44524: result <= 12'b111100111001;
   44525: result <= 12'b111100111001;
   44526: result <= 12'b111100111001;
   44527: result <= 12'b111100111001;
   44528: result <= 12'b111100111010;
   44529: result <= 12'b111100111010;
   44530: result <= 12'b111100111010;
   44531: result <= 12'b111100111010;
   44532: result <= 12'b111100111010;
   44533: result <= 12'b111100111010;
   44534: result <= 12'b111100111010;
   44535: result <= 12'b111100111010;
   44536: result <= 12'b111100111010;
   44537: result <= 12'b111100111010;
   44538: result <= 12'b111100111010;
   44539: result <= 12'b111100111010;
   44540: result <= 12'b111100111011;
   44541: result <= 12'b111100111011;
   44542: result <= 12'b111100111011;
   44543: result <= 12'b111100111011;
   44544: result <= 12'b111100111011;
   44545: result <= 12'b111100111011;
   44546: result <= 12'b111100111011;
   44547: result <= 12'b111100111011;
   44548: result <= 12'b111100111011;
   44549: result <= 12'b111100111011;
   44550: result <= 12'b111100111011;
   44551: result <= 12'b111100111011;
   44552: result <= 12'b111100111100;
   44553: result <= 12'b111100111100;
   44554: result <= 12'b111100111100;
   44555: result <= 12'b111100111100;
   44556: result <= 12'b111100111100;
   44557: result <= 12'b111100111100;
   44558: result <= 12'b111100111100;
   44559: result <= 12'b111100111100;
   44560: result <= 12'b111100111100;
   44561: result <= 12'b111100111100;
   44562: result <= 12'b111100111100;
   44563: result <= 12'b111100111100;
   44564: result <= 12'b111100111101;
   44565: result <= 12'b111100111101;
   44566: result <= 12'b111100111101;
   44567: result <= 12'b111100111101;
   44568: result <= 12'b111100111101;
   44569: result <= 12'b111100111101;
   44570: result <= 12'b111100111101;
   44571: result <= 12'b111100111101;
   44572: result <= 12'b111100111101;
   44573: result <= 12'b111100111101;
   44574: result <= 12'b111100111101;
   44575: result <= 12'b111100111101;
   44576: result <= 12'b111100111110;
   44577: result <= 12'b111100111110;
   44578: result <= 12'b111100111110;
   44579: result <= 12'b111100111110;
   44580: result <= 12'b111100111110;
   44581: result <= 12'b111100111110;
   44582: result <= 12'b111100111110;
   44583: result <= 12'b111100111110;
   44584: result <= 12'b111100111110;
   44585: result <= 12'b111100111110;
   44586: result <= 12'b111100111110;
   44587: result <= 12'b111100111110;
   44588: result <= 12'b111100111111;
   44589: result <= 12'b111100111111;
   44590: result <= 12'b111100111111;
   44591: result <= 12'b111100111111;
   44592: result <= 12'b111100111111;
   44593: result <= 12'b111100111111;
   44594: result <= 12'b111100111111;
   44595: result <= 12'b111100111111;
   44596: result <= 12'b111100111111;
   44597: result <= 12'b111100111111;
   44598: result <= 12'b111100111111;
   44599: result <= 12'b111100111111;
   44600: result <= 12'b111101000000;
   44601: result <= 12'b111101000000;
   44602: result <= 12'b111101000000;
   44603: result <= 12'b111101000000;
   44604: result <= 12'b111101000000;
   44605: result <= 12'b111101000000;
   44606: result <= 12'b111101000000;
   44607: result <= 12'b111101000000;
   44608: result <= 12'b111101000000;
   44609: result <= 12'b111101000000;
   44610: result <= 12'b111101000000;
   44611: result <= 12'b111101000000;
   44612: result <= 12'b111101000001;
   44613: result <= 12'b111101000001;
   44614: result <= 12'b111101000001;
   44615: result <= 12'b111101000001;
   44616: result <= 12'b111101000001;
   44617: result <= 12'b111101000001;
   44618: result <= 12'b111101000001;
   44619: result <= 12'b111101000001;
   44620: result <= 12'b111101000001;
   44621: result <= 12'b111101000001;
   44622: result <= 12'b111101000001;
   44623: result <= 12'b111101000001;
   44624: result <= 12'b111101000010;
   44625: result <= 12'b111101000010;
   44626: result <= 12'b111101000010;
   44627: result <= 12'b111101000010;
   44628: result <= 12'b111101000010;
   44629: result <= 12'b111101000010;
   44630: result <= 12'b111101000010;
   44631: result <= 12'b111101000010;
   44632: result <= 12'b111101000010;
   44633: result <= 12'b111101000010;
   44634: result <= 12'b111101000010;
   44635: result <= 12'b111101000010;
   44636: result <= 12'b111101000011;
   44637: result <= 12'b111101000011;
   44638: result <= 12'b111101000011;
   44639: result <= 12'b111101000011;
   44640: result <= 12'b111101000011;
   44641: result <= 12'b111101000011;
   44642: result <= 12'b111101000011;
   44643: result <= 12'b111101000011;
   44644: result <= 12'b111101000011;
   44645: result <= 12'b111101000011;
   44646: result <= 12'b111101000011;
   44647: result <= 12'b111101000011;
   44648: result <= 12'b111101000100;
   44649: result <= 12'b111101000100;
   44650: result <= 12'b111101000100;
   44651: result <= 12'b111101000100;
   44652: result <= 12'b111101000100;
   44653: result <= 12'b111101000100;
   44654: result <= 12'b111101000100;
   44655: result <= 12'b111101000100;
   44656: result <= 12'b111101000100;
   44657: result <= 12'b111101000100;
   44658: result <= 12'b111101000100;
   44659: result <= 12'b111101000100;
   44660: result <= 12'b111101000100;
   44661: result <= 12'b111101000101;
   44662: result <= 12'b111101000101;
   44663: result <= 12'b111101000101;
   44664: result <= 12'b111101000101;
   44665: result <= 12'b111101000101;
   44666: result <= 12'b111101000101;
   44667: result <= 12'b111101000101;
   44668: result <= 12'b111101000101;
   44669: result <= 12'b111101000101;
   44670: result <= 12'b111101000101;
   44671: result <= 12'b111101000101;
   44672: result <= 12'b111101000101;
   44673: result <= 12'b111101000110;
   44674: result <= 12'b111101000110;
   44675: result <= 12'b111101000110;
   44676: result <= 12'b111101000110;
   44677: result <= 12'b111101000110;
   44678: result <= 12'b111101000110;
   44679: result <= 12'b111101000110;
   44680: result <= 12'b111101000110;
   44681: result <= 12'b111101000110;
   44682: result <= 12'b111101000110;
   44683: result <= 12'b111101000110;
   44684: result <= 12'b111101000110;
   44685: result <= 12'b111101000111;
   44686: result <= 12'b111101000111;
   44687: result <= 12'b111101000111;
   44688: result <= 12'b111101000111;
   44689: result <= 12'b111101000111;
   44690: result <= 12'b111101000111;
   44691: result <= 12'b111101000111;
   44692: result <= 12'b111101000111;
   44693: result <= 12'b111101000111;
   44694: result <= 12'b111101000111;
   44695: result <= 12'b111101000111;
   44696: result <= 12'b111101000111;
   44697: result <= 12'b111101001000;
   44698: result <= 12'b111101001000;
   44699: result <= 12'b111101001000;
   44700: result <= 12'b111101001000;
   44701: result <= 12'b111101001000;
   44702: result <= 12'b111101001000;
   44703: result <= 12'b111101001000;
   44704: result <= 12'b111101001000;
   44705: result <= 12'b111101001000;
   44706: result <= 12'b111101001000;
   44707: result <= 12'b111101001000;
   44708: result <= 12'b111101001000;
   44709: result <= 12'b111101001000;
   44710: result <= 12'b111101001001;
   44711: result <= 12'b111101001001;
   44712: result <= 12'b111101001001;
   44713: result <= 12'b111101001001;
   44714: result <= 12'b111101001001;
   44715: result <= 12'b111101001001;
   44716: result <= 12'b111101001001;
   44717: result <= 12'b111101001001;
   44718: result <= 12'b111101001001;
   44719: result <= 12'b111101001001;
   44720: result <= 12'b111101001001;
   44721: result <= 12'b111101001001;
   44722: result <= 12'b111101001010;
   44723: result <= 12'b111101001010;
   44724: result <= 12'b111101001010;
   44725: result <= 12'b111101001010;
   44726: result <= 12'b111101001010;
   44727: result <= 12'b111101001010;
   44728: result <= 12'b111101001010;
   44729: result <= 12'b111101001010;
   44730: result <= 12'b111101001010;
   44731: result <= 12'b111101001010;
   44732: result <= 12'b111101001010;
   44733: result <= 12'b111101001010;
   44734: result <= 12'b111101001011;
   44735: result <= 12'b111101001011;
   44736: result <= 12'b111101001011;
   44737: result <= 12'b111101001011;
   44738: result <= 12'b111101001011;
   44739: result <= 12'b111101001011;
   44740: result <= 12'b111101001011;
   44741: result <= 12'b111101001011;
   44742: result <= 12'b111101001011;
   44743: result <= 12'b111101001011;
   44744: result <= 12'b111101001011;
   44745: result <= 12'b111101001011;
   44746: result <= 12'b111101001011;
   44747: result <= 12'b111101001100;
   44748: result <= 12'b111101001100;
   44749: result <= 12'b111101001100;
   44750: result <= 12'b111101001100;
   44751: result <= 12'b111101001100;
   44752: result <= 12'b111101001100;
   44753: result <= 12'b111101001100;
   44754: result <= 12'b111101001100;
   44755: result <= 12'b111101001100;
   44756: result <= 12'b111101001100;
   44757: result <= 12'b111101001100;
   44758: result <= 12'b111101001100;
   44759: result <= 12'b111101001101;
   44760: result <= 12'b111101001101;
   44761: result <= 12'b111101001101;
   44762: result <= 12'b111101001101;
   44763: result <= 12'b111101001101;
   44764: result <= 12'b111101001101;
   44765: result <= 12'b111101001101;
   44766: result <= 12'b111101001101;
   44767: result <= 12'b111101001101;
   44768: result <= 12'b111101001101;
   44769: result <= 12'b111101001101;
   44770: result <= 12'b111101001101;
   44771: result <= 12'b111101001101;
   44772: result <= 12'b111101001110;
   44773: result <= 12'b111101001110;
   44774: result <= 12'b111101001110;
   44775: result <= 12'b111101001110;
   44776: result <= 12'b111101001110;
   44777: result <= 12'b111101001110;
   44778: result <= 12'b111101001110;
   44779: result <= 12'b111101001110;
   44780: result <= 12'b111101001110;
   44781: result <= 12'b111101001110;
   44782: result <= 12'b111101001110;
   44783: result <= 12'b111101001110;
   44784: result <= 12'b111101001111;
   44785: result <= 12'b111101001111;
   44786: result <= 12'b111101001111;
   44787: result <= 12'b111101001111;
   44788: result <= 12'b111101001111;
   44789: result <= 12'b111101001111;
   44790: result <= 12'b111101001111;
   44791: result <= 12'b111101001111;
   44792: result <= 12'b111101001111;
   44793: result <= 12'b111101001111;
   44794: result <= 12'b111101001111;
   44795: result <= 12'b111101001111;
   44796: result <= 12'b111101001111;
   44797: result <= 12'b111101010000;
   44798: result <= 12'b111101010000;
   44799: result <= 12'b111101010000;
   44800: result <= 12'b111101010000;
   44801: result <= 12'b111101010000;
   44802: result <= 12'b111101010000;
   44803: result <= 12'b111101010000;
   44804: result <= 12'b111101010000;
   44805: result <= 12'b111101010000;
   44806: result <= 12'b111101010000;
   44807: result <= 12'b111101010000;
   44808: result <= 12'b111101010000;
   44809: result <= 12'b111101010001;
   44810: result <= 12'b111101010001;
   44811: result <= 12'b111101010001;
   44812: result <= 12'b111101010001;
   44813: result <= 12'b111101010001;
   44814: result <= 12'b111101010001;
   44815: result <= 12'b111101010001;
   44816: result <= 12'b111101010001;
   44817: result <= 12'b111101010001;
   44818: result <= 12'b111101010001;
   44819: result <= 12'b111101010001;
   44820: result <= 12'b111101010001;
   44821: result <= 12'b111101010001;
   44822: result <= 12'b111101010010;
   44823: result <= 12'b111101010010;
   44824: result <= 12'b111101010010;
   44825: result <= 12'b111101010010;
   44826: result <= 12'b111101010010;
   44827: result <= 12'b111101010010;
   44828: result <= 12'b111101010010;
   44829: result <= 12'b111101010010;
   44830: result <= 12'b111101010010;
   44831: result <= 12'b111101010010;
   44832: result <= 12'b111101010010;
   44833: result <= 12'b111101010010;
   44834: result <= 12'b111101010010;
   44835: result <= 12'b111101010011;
   44836: result <= 12'b111101010011;
   44837: result <= 12'b111101010011;
   44838: result <= 12'b111101010011;
   44839: result <= 12'b111101010011;
   44840: result <= 12'b111101010011;
   44841: result <= 12'b111101010011;
   44842: result <= 12'b111101010011;
   44843: result <= 12'b111101010011;
   44844: result <= 12'b111101010011;
   44845: result <= 12'b111101010011;
   44846: result <= 12'b111101010011;
   44847: result <= 12'b111101010100;
   44848: result <= 12'b111101010100;
   44849: result <= 12'b111101010100;
   44850: result <= 12'b111101010100;
   44851: result <= 12'b111101010100;
   44852: result <= 12'b111101010100;
   44853: result <= 12'b111101010100;
   44854: result <= 12'b111101010100;
   44855: result <= 12'b111101010100;
   44856: result <= 12'b111101010100;
   44857: result <= 12'b111101010100;
   44858: result <= 12'b111101010100;
   44859: result <= 12'b111101010100;
   44860: result <= 12'b111101010101;
   44861: result <= 12'b111101010101;
   44862: result <= 12'b111101010101;
   44863: result <= 12'b111101010101;
   44864: result <= 12'b111101010101;
   44865: result <= 12'b111101010101;
   44866: result <= 12'b111101010101;
   44867: result <= 12'b111101010101;
   44868: result <= 12'b111101010101;
   44869: result <= 12'b111101010101;
   44870: result <= 12'b111101010101;
   44871: result <= 12'b111101010101;
   44872: result <= 12'b111101010101;
   44873: result <= 12'b111101010110;
   44874: result <= 12'b111101010110;
   44875: result <= 12'b111101010110;
   44876: result <= 12'b111101010110;
   44877: result <= 12'b111101010110;
   44878: result <= 12'b111101010110;
   44879: result <= 12'b111101010110;
   44880: result <= 12'b111101010110;
   44881: result <= 12'b111101010110;
   44882: result <= 12'b111101010110;
   44883: result <= 12'b111101010110;
   44884: result <= 12'b111101010110;
   44885: result <= 12'b111101010111;
   44886: result <= 12'b111101010111;
   44887: result <= 12'b111101010111;
   44888: result <= 12'b111101010111;
   44889: result <= 12'b111101010111;
   44890: result <= 12'b111101010111;
   44891: result <= 12'b111101010111;
   44892: result <= 12'b111101010111;
   44893: result <= 12'b111101010111;
   44894: result <= 12'b111101010111;
   44895: result <= 12'b111101010111;
   44896: result <= 12'b111101010111;
   44897: result <= 12'b111101010111;
   44898: result <= 12'b111101011000;
   44899: result <= 12'b111101011000;
   44900: result <= 12'b111101011000;
   44901: result <= 12'b111101011000;
   44902: result <= 12'b111101011000;
   44903: result <= 12'b111101011000;
   44904: result <= 12'b111101011000;
   44905: result <= 12'b111101011000;
   44906: result <= 12'b111101011000;
   44907: result <= 12'b111101011000;
   44908: result <= 12'b111101011000;
   44909: result <= 12'b111101011000;
   44910: result <= 12'b111101011000;
   44911: result <= 12'b111101011001;
   44912: result <= 12'b111101011001;
   44913: result <= 12'b111101011001;
   44914: result <= 12'b111101011001;
   44915: result <= 12'b111101011001;
   44916: result <= 12'b111101011001;
   44917: result <= 12'b111101011001;
   44918: result <= 12'b111101011001;
   44919: result <= 12'b111101011001;
   44920: result <= 12'b111101011001;
   44921: result <= 12'b111101011001;
   44922: result <= 12'b111101011001;
   44923: result <= 12'b111101011001;
   44924: result <= 12'b111101011010;
   44925: result <= 12'b111101011010;
   44926: result <= 12'b111101011010;
   44927: result <= 12'b111101011010;
   44928: result <= 12'b111101011010;
   44929: result <= 12'b111101011010;
   44930: result <= 12'b111101011010;
   44931: result <= 12'b111101011010;
   44932: result <= 12'b111101011010;
   44933: result <= 12'b111101011010;
   44934: result <= 12'b111101011010;
   44935: result <= 12'b111101011010;
   44936: result <= 12'b111101011010;
   44937: result <= 12'b111101011011;
   44938: result <= 12'b111101011011;
   44939: result <= 12'b111101011011;
   44940: result <= 12'b111101011011;
   44941: result <= 12'b111101011011;
   44942: result <= 12'b111101011011;
   44943: result <= 12'b111101011011;
   44944: result <= 12'b111101011011;
   44945: result <= 12'b111101011011;
   44946: result <= 12'b111101011011;
   44947: result <= 12'b111101011011;
   44948: result <= 12'b111101011011;
   44949: result <= 12'b111101011011;
   44950: result <= 12'b111101011100;
   44951: result <= 12'b111101011100;
   44952: result <= 12'b111101011100;
   44953: result <= 12'b111101011100;
   44954: result <= 12'b111101011100;
   44955: result <= 12'b111101011100;
   44956: result <= 12'b111101011100;
   44957: result <= 12'b111101011100;
   44958: result <= 12'b111101011100;
   44959: result <= 12'b111101011100;
   44960: result <= 12'b111101011100;
   44961: result <= 12'b111101011100;
   44962: result <= 12'b111101011100;
   44963: result <= 12'b111101011101;
   44964: result <= 12'b111101011101;
   44965: result <= 12'b111101011101;
   44966: result <= 12'b111101011101;
   44967: result <= 12'b111101011101;
   44968: result <= 12'b111101011101;
   44969: result <= 12'b111101011101;
   44970: result <= 12'b111101011101;
   44971: result <= 12'b111101011101;
   44972: result <= 12'b111101011101;
   44973: result <= 12'b111101011101;
   44974: result <= 12'b111101011101;
   44975: result <= 12'b111101011101;
   44976: result <= 12'b111101011110;
   44977: result <= 12'b111101011110;
   44978: result <= 12'b111101011110;
   44979: result <= 12'b111101011110;
   44980: result <= 12'b111101011110;
   44981: result <= 12'b111101011110;
   44982: result <= 12'b111101011110;
   44983: result <= 12'b111101011110;
   44984: result <= 12'b111101011110;
   44985: result <= 12'b111101011110;
   44986: result <= 12'b111101011110;
   44987: result <= 12'b111101011110;
   44988: result <= 12'b111101011110;
   44989: result <= 12'b111101011111;
   44990: result <= 12'b111101011111;
   44991: result <= 12'b111101011111;
   44992: result <= 12'b111101011111;
   44993: result <= 12'b111101011111;
   44994: result <= 12'b111101011111;
   44995: result <= 12'b111101011111;
   44996: result <= 12'b111101011111;
   44997: result <= 12'b111101011111;
   44998: result <= 12'b111101011111;
   44999: result <= 12'b111101011111;
   45000: result <= 12'b111101011111;
   45001: result <= 12'b111101011111;
   45002: result <= 12'b111101100000;
   45003: result <= 12'b111101100000;
   45004: result <= 12'b111101100000;
   45005: result <= 12'b111101100000;
   45006: result <= 12'b111101100000;
   45007: result <= 12'b111101100000;
   45008: result <= 12'b111101100000;
   45009: result <= 12'b111101100000;
   45010: result <= 12'b111101100000;
   45011: result <= 12'b111101100000;
   45012: result <= 12'b111101100000;
   45013: result <= 12'b111101100000;
   45014: result <= 12'b111101100000;
   45015: result <= 12'b111101100001;
   45016: result <= 12'b111101100001;
   45017: result <= 12'b111101100001;
   45018: result <= 12'b111101100001;
   45019: result <= 12'b111101100001;
   45020: result <= 12'b111101100001;
   45021: result <= 12'b111101100001;
   45022: result <= 12'b111101100001;
   45023: result <= 12'b111101100001;
   45024: result <= 12'b111101100001;
   45025: result <= 12'b111101100001;
   45026: result <= 12'b111101100001;
   45027: result <= 12'b111101100001;
   45028: result <= 12'b111101100001;
   45029: result <= 12'b111101100010;
   45030: result <= 12'b111101100010;
   45031: result <= 12'b111101100010;
   45032: result <= 12'b111101100010;
   45033: result <= 12'b111101100010;
   45034: result <= 12'b111101100010;
   45035: result <= 12'b111101100010;
   45036: result <= 12'b111101100010;
   45037: result <= 12'b111101100010;
   45038: result <= 12'b111101100010;
   45039: result <= 12'b111101100010;
   45040: result <= 12'b111101100010;
   45041: result <= 12'b111101100010;
   45042: result <= 12'b111101100011;
   45043: result <= 12'b111101100011;
   45044: result <= 12'b111101100011;
   45045: result <= 12'b111101100011;
   45046: result <= 12'b111101100011;
   45047: result <= 12'b111101100011;
   45048: result <= 12'b111101100011;
   45049: result <= 12'b111101100011;
   45050: result <= 12'b111101100011;
   45051: result <= 12'b111101100011;
   45052: result <= 12'b111101100011;
   45053: result <= 12'b111101100011;
   45054: result <= 12'b111101100011;
   45055: result <= 12'b111101100100;
   45056: result <= 12'b111101100100;
   45057: result <= 12'b111101100100;
   45058: result <= 12'b111101100100;
   45059: result <= 12'b111101100100;
   45060: result <= 12'b111101100100;
   45061: result <= 12'b111101100100;
   45062: result <= 12'b111101100100;
   45063: result <= 12'b111101100100;
   45064: result <= 12'b111101100100;
   45065: result <= 12'b111101100100;
   45066: result <= 12'b111101100100;
   45067: result <= 12'b111101100100;
   45068: result <= 12'b111101100101;
   45069: result <= 12'b111101100101;
   45070: result <= 12'b111101100101;
   45071: result <= 12'b111101100101;
   45072: result <= 12'b111101100101;
   45073: result <= 12'b111101100101;
   45074: result <= 12'b111101100101;
   45075: result <= 12'b111101100101;
   45076: result <= 12'b111101100101;
   45077: result <= 12'b111101100101;
   45078: result <= 12'b111101100101;
   45079: result <= 12'b111101100101;
   45080: result <= 12'b111101100101;
   45081: result <= 12'b111101100101;
   45082: result <= 12'b111101100110;
   45083: result <= 12'b111101100110;
   45084: result <= 12'b111101100110;
   45085: result <= 12'b111101100110;
   45086: result <= 12'b111101100110;
   45087: result <= 12'b111101100110;
   45088: result <= 12'b111101100110;
   45089: result <= 12'b111101100110;
   45090: result <= 12'b111101100110;
   45091: result <= 12'b111101100110;
   45092: result <= 12'b111101100110;
   45093: result <= 12'b111101100110;
   45094: result <= 12'b111101100110;
   45095: result <= 12'b111101100111;
   45096: result <= 12'b111101100111;
   45097: result <= 12'b111101100111;
   45098: result <= 12'b111101100111;
   45099: result <= 12'b111101100111;
   45100: result <= 12'b111101100111;
   45101: result <= 12'b111101100111;
   45102: result <= 12'b111101100111;
   45103: result <= 12'b111101100111;
   45104: result <= 12'b111101100111;
   45105: result <= 12'b111101100111;
   45106: result <= 12'b111101100111;
   45107: result <= 12'b111101100111;
   45108: result <= 12'b111101100111;
   45109: result <= 12'b111101101000;
   45110: result <= 12'b111101101000;
   45111: result <= 12'b111101101000;
   45112: result <= 12'b111101101000;
   45113: result <= 12'b111101101000;
   45114: result <= 12'b111101101000;
   45115: result <= 12'b111101101000;
   45116: result <= 12'b111101101000;
   45117: result <= 12'b111101101000;
   45118: result <= 12'b111101101000;
   45119: result <= 12'b111101101000;
   45120: result <= 12'b111101101000;
   45121: result <= 12'b111101101000;
   45122: result <= 12'b111101101001;
   45123: result <= 12'b111101101001;
   45124: result <= 12'b111101101001;
   45125: result <= 12'b111101101001;
   45126: result <= 12'b111101101001;
   45127: result <= 12'b111101101001;
   45128: result <= 12'b111101101001;
   45129: result <= 12'b111101101001;
   45130: result <= 12'b111101101001;
   45131: result <= 12'b111101101001;
   45132: result <= 12'b111101101001;
   45133: result <= 12'b111101101001;
   45134: result <= 12'b111101101001;
   45135: result <= 12'b111101101001;
   45136: result <= 12'b111101101010;
   45137: result <= 12'b111101101010;
   45138: result <= 12'b111101101010;
   45139: result <= 12'b111101101010;
   45140: result <= 12'b111101101010;
   45141: result <= 12'b111101101010;
   45142: result <= 12'b111101101010;
   45143: result <= 12'b111101101010;
   45144: result <= 12'b111101101010;
   45145: result <= 12'b111101101010;
   45146: result <= 12'b111101101010;
   45147: result <= 12'b111101101010;
   45148: result <= 12'b111101101010;
   45149: result <= 12'b111101101011;
   45150: result <= 12'b111101101011;
   45151: result <= 12'b111101101011;
   45152: result <= 12'b111101101011;
   45153: result <= 12'b111101101011;
   45154: result <= 12'b111101101011;
   45155: result <= 12'b111101101011;
   45156: result <= 12'b111101101011;
   45157: result <= 12'b111101101011;
   45158: result <= 12'b111101101011;
   45159: result <= 12'b111101101011;
   45160: result <= 12'b111101101011;
   45161: result <= 12'b111101101011;
   45162: result <= 12'b111101101011;
   45163: result <= 12'b111101101100;
   45164: result <= 12'b111101101100;
   45165: result <= 12'b111101101100;
   45166: result <= 12'b111101101100;
   45167: result <= 12'b111101101100;
   45168: result <= 12'b111101101100;
   45169: result <= 12'b111101101100;
   45170: result <= 12'b111101101100;
   45171: result <= 12'b111101101100;
   45172: result <= 12'b111101101100;
   45173: result <= 12'b111101101100;
   45174: result <= 12'b111101101100;
   45175: result <= 12'b111101101100;
   45176: result <= 12'b111101101100;
   45177: result <= 12'b111101101101;
   45178: result <= 12'b111101101101;
   45179: result <= 12'b111101101101;
   45180: result <= 12'b111101101101;
   45181: result <= 12'b111101101101;
   45182: result <= 12'b111101101101;
   45183: result <= 12'b111101101101;
   45184: result <= 12'b111101101101;
   45185: result <= 12'b111101101101;
   45186: result <= 12'b111101101101;
   45187: result <= 12'b111101101101;
   45188: result <= 12'b111101101101;
   45189: result <= 12'b111101101101;
   45190: result <= 12'b111101101110;
   45191: result <= 12'b111101101110;
   45192: result <= 12'b111101101110;
   45193: result <= 12'b111101101110;
   45194: result <= 12'b111101101110;
   45195: result <= 12'b111101101110;
   45196: result <= 12'b111101101110;
   45197: result <= 12'b111101101110;
   45198: result <= 12'b111101101110;
   45199: result <= 12'b111101101110;
   45200: result <= 12'b111101101110;
   45201: result <= 12'b111101101110;
   45202: result <= 12'b111101101110;
   45203: result <= 12'b111101101110;
   45204: result <= 12'b111101101111;
   45205: result <= 12'b111101101111;
   45206: result <= 12'b111101101111;
   45207: result <= 12'b111101101111;
   45208: result <= 12'b111101101111;
   45209: result <= 12'b111101101111;
   45210: result <= 12'b111101101111;
   45211: result <= 12'b111101101111;
   45212: result <= 12'b111101101111;
   45213: result <= 12'b111101101111;
   45214: result <= 12'b111101101111;
   45215: result <= 12'b111101101111;
   45216: result <= 12'b111101101111;
   45217: result <= 12'b111101101111;
   45218: result <= 12'b111101110000;
   45219: result <= 12'b111101110000;
   45220: result <= 12'b111101110000;
   45221: result <= 12'b111101110000;
   45222: result <= 12'b111101110000;
   45223: result <= 12'b111101110000;
   45224: result <= 12'b111101110000;
   45225: result <= 12'b111101110000;
   45226: result <= 12'b111101110000;
   45227: result <= 12'b111101110000;
   45228: result <= 12'b111101110000;
   45229: result <= 12'b111101110000;
   45230: result <= 12'b111101110000;
   45231: result <= 12'b111101110000;
   45232: result <= 12'b111101110001;
   45233: result <= 12'b111101110001;
   45234: result <= 12'b111101110001;
   45235: result <= 12'b111101110001;
   45236: result <= 12'b111101110001;
   45237: result <= 12'b111101110001;
   45238: result <= 12'b111101110001;
   45239: result <= 12'b111101110001;
   45240: result <= 12'b111101110001;
   45241: result <= 12'b111101110001;
   45242: result <= 12'b111101110001;
   45243: result <= 12'b111101110001;
   45244: result <= 12'b111101110001;
   45245: result <= 12'b111101110001;
   45246: result <= 12'b111101110010;
   45247: result <= 12'b111101110010;
   45248: result <= 12'b111101110010;
   45249: result <= 12'b111101110010;
   45250: result <= 12'b111101110010;
   45251: result <= 12'b111101110010;
   45252: result <= 12'b111101110010;
   45253: result <= 12'b111101110010;
   45254: result <= 12'b111101110010;
   45255: result <= 12'b111101110010;
   45256: result <= 12'b111101110010;
   45257: result <= 12'b111101110010;
   45258: result <= 12'b111101110010;
   45259: result <= 12'b111101110010;
   45260: result <= 12'b111101110011;
   45261: result <= 12'b111101110011;
   45262: result <= 12'b111101110011;
   45263: result <= 12'b111101110011;
   45264: result <= 12'b111101110011;
   45265: result <= 12'b111101110011;
   45266: result <= 12'b111101110011;
   45267: result <= 12'b111101110011;
   45268: result <= 12'b111101110011;
   45269: result <= 12'b111101110011;
   45270: result <= 12'b111101110011;
   45271: result <= 12'b111101110011;
   45272: result <= 12'b111101110011;
   45273: result <= 12'b111101110011;
   45274: result <= 12'b111101110100;
   45275: result <= 12'b111101110100;
   45276: result <= 12'b111101110100;
   45277: result <= 12'b111101110100;
   45278: result <= 12'b111101110100;
   45279: result <= 12'b111101110100;
   45280: result <= 12'b111101110100;
   45281: result <= 12'b111101110100;
   45282: result <= 12'b111101110100;
   45283: result <= 12'b111101110100;
   45284: result <= 12'b111101110100;
   45285: result <= 12'b111101110100;
   45286: result <= 12'b111101110100;
   45287: result <= 12'b111101110100;
   45288: result <= 12'b111101110101;
   45289: result <= 12'b111101110101;
   45290: result <= 12'b111101110101;
   45291: result <= 12'b111101110101;
   45292: result <= 12'b111101110101;
   45293: result <= 12'b111101110101;
   45294: result <= 12'b111101110101;
   45295: result <= 12'b111101110101;
   45296: result <= 12'b111101110101;
   45297: result <= 12'b111101110101;
   45298: result <= 12'b111101110101;
   45299: result <= 12'b111101110101;
   45300: result <= 12'b111101110101;
   45301: result <= 12'b111101110101;
   45302: result <= 12'b111101110110;
   45303: result <= 12'b111101110110;
   45304: result <= 12'b111101110110;
   45305: result <= 12'b111101110110;
   45306: result <= 12'b111101110110;
   45307: result <= 12'b111101110110;
   45308: result <= 12'b111101110110;
   45309: result <= 12'b111101110110;
   45310: result <= 12'b111101110110;
   45311: result <= 12'b111101110110;
   45312: result <= 12'b111101110110;
   45313: result <= 12'b111101110110;
   45314: result <= 12'b111101110110;
   45315: result <= 12'b111101110110;
   45316: result <= 12'b111101110111;
   45317: result <= 12'b111101110111;
   45318: result <= 12'b111101110111;
   45319: result <= 12'b111101110111;
   45320: result <= 12'b111101110111;
   45321: result <= 12'b111101110111;
   45322: result <= 12'b111101110111;
   45323: result <= 12'b111101110111;
   45324: result <= 12'b111101110111;
   45325: result <= 12'b111101110111;
   45326: result <= 12'b111101110111;
   45327: result <= 12'b111101110111;
   45328: result <= 12'b111101110111;
   45329: result <= 12'b111101110111;
   45330: result <= 12'b111101111000;
   45331: result <= 12'b111101111000;
   45332: result <= 12'b111101111000;
   45333: result <= 12'b111101111000;
   45334: result <= 12'b111101111000;
   45335: result <= 12'b111101111000;
   45336: result <= 12'b111101111000;
   45337: result <= 12'b111101111000;
   45338: result <= 12'b111101111000;
   45339: result <= 12'b111101111000;
   45340: result <= 12'b111101111000;
   45341: result <= 12'b111101111000;
   45342: result <= 12'b111101111000;
   45343: result <= 12'b111101111000;
   45344: result <= 12'b111101111001;
   45345: result <= 12'b111101111001;
   45346: result <= 12'b111101111001;
   45347: result <= 12'b111101111001;
   45348: result <= 12'b111101111001;
   45349: result <= 12'b111101111001;
   45350: result <= 12'b111101111001;
   45351: result <= 12'b111101111001;
   45352: result <= 12'b111101111001;
   45353: result <= 12'b111101111001;
   45354: result <= 12'b111101111001;
   45355: result <= 12'b111101111001;
   45356: result <= 12'b111101111001;
   45357: result <= 12'b111101111001;
   45358: result <= 12'b111101111010;
   45359: result <= 12'b111101111010;
   45360: result <= 12'b111101111010;
   45361: result <= 12'b111101111010;
   45362: result <= 12'b111101111010;
   45363: result <= 12'b111101111010;
   45364: result <= 12'b111101111010;
   45365: result <= 12'b111101111010;
   45366: result <= 12'b111101111010;
   45367: result <= 12'b111101111010;
   45368: result <= 12'b111101111010;
   45369: result <= 12'b111101111010;
   45370: result <= 12'b111101111010;
   45371: result <= 12'b111101111010;
   45372: result <= 12'b111101111010;
   45373: result <= 12'b111101111011;
   45374: result <= 12'b111101111011;
   45375: result <= 12'b111101111011;
   45376: result <= 12'b111101111011;
   45377: result <= 12'b111101111011;
   45378: result <= 12'b111101111011;
   45379: result <= 12'b111101111011;
   45380: result <= 12'b111101111011;
   45381: result <= 12'b111101111011;
   45382: result <= 12'b111101111011;
   45383: result <= 12'b111101111011;
   45384: result <= 12'b111101111011;
   45385: result <= 12'b111101111011;
   45386: result <= 12'b111101111011;
   45387: result <= 12'b111101111100;
   45388: result <= 12'b111101111100;
   45389: result <= 12'b111101111100;
   45390: result <= 12'b111101111100;
   45391: result <= 12'b111101111100;
   45392: result <= 12'b111101111100;
   45393: result <= 12'b111101111100;
   45394: result <= 12'b111101111100;
   45395: result <= 12'b111101111100;
   45396: result <= 12'b111101111100;
   45397: result <= 12'b111101111100;
   45398: result <= 12'b111101111100;
   45399: result <= 12'b111101111100;
   45400: result <= 12'b111101111100;
   45401: result <= 12'b111101111100;
   45402: result <= 12'b111101111101;
   45403: result <= 12'b111101111101;
   45404: result <= 12'b111101111101;
   45405: result <= 12'b111101111101;
   45406: result <= 12'b111101111101;
   45407: result <= 12'b111101111101;
   45408: result <= 12'b111101111101;
   45409: result <= 12'b111101111101;
   45410: result <= 12'b111101111101;
   45411: result <= 12'b111101111101;
   45412: result <= 12'b111101111101;
   45413: result <= 12'b111101111101;
   45414: result <= 12'b111101111101;
   45415: result <= 12'b111101111101;
   45416: result <= 12'b111101111110;
   45417: result <= 12'b111101111110;
   45418: result <= 12'b111101111110;
   45419: result <= 12'b111101111110;
   45420: result <= 12'b111101111110;
   45421: result <= 12'b111101111110;
   45422: result <= 12'b111101111110;
   45423: result <= 12'b111101111110;
   45424: result <= 12'b111101111110;
   45425: result <= 12'b111101111110;
   45426: result <= 12'b111101111110;
   45427: result <= 12'b111101111110;
   45428: result <= 12'b111101111110;
   45429: result <= 12'b111101111110;
   45430: result <= 12'b111101111110;
   45431: result <= 12'b111101111111;
   45432: result <= 12'b111101111111;
   45433: result <= 12'b111101111111;
   45434: result <= 12'b111101111111;
   45435: result <= 12'b111101111111;
   45436: result <= 12'b111101111111;
   45437: result <= 12'b111101111111;
   45438: result <= 12'b111101111111;
   45439: result <= 12'b111101111111;
   45440: result <= 12'b111101111111;
   45441: result <= 12'b111101111111;
   45442: result <= 12'b111101111111;
   45443: result <= 12'b111101111111;
   45444: result <= 12'b111101111111;
   45445: result <= 12'b111110000000;
   45446: result <= 12'b111110000000;
   45447: result <= 12'b111110000000;
   45448: result <= 12'b111110000000;
   45449: result <= 12'b111110000000;
   45450: result <= 12'b111110000000;
   45451: result <= 12'b111110000000;
   45452: result <= 12'b111110000000;
   45453: result <= 12'b111110000000;
   45454: result <= 12'b111110000000;
   45455: result <= 12'b111110000000;
   45456: result <= 12'b111110000000;
   45457: result <= 12'b111110000000;
   45458: result <= 12'b111110000000;
   45459: result <= 12'b111110000000;
   45460: result <= 12'b111110000001;
   45461: result <= 12'b111110000001;
   45462: result <= 12'b111110000001;
   45463: result <= 12'b111110000001;
   45464: result <= 12'b111110000001;
   45465: result <= 12'b111110000001;
   45466: result <= 12'b111110000001;
   45467: result <= 12'b111110000001;
   45468: result <= 12'b111110000001;
   45469: result <= 12'b111110000001;
   45470: result <= 12'b111110000001;
   45471: result <= 12'b111110000001;
   45472: result <= 12'b111110000001;
   45473: result <= 12'b111110000001;
   45474: result <= 12'b111110000001;
   45475: result <= 12'b111110000010;
   45476: result <= 12'b111110000010;
   45477: result <= 12'b111110000010;
   45478: result <= 12'b111110000010;
   45479: result <= 12'b111110000010;
   45480: result <= 12'b111110000010;
   45481: result <= 12'b111110000010;
   45482: result <= 12'b111110000010;
   45483: result <= 12'b111110000010;
   45484: result <= 12'b111110000010;
   45485: result <= 12'b111110000010;
   45486: result <= 12'b111110000010;
   45487: result <= 12'b111110000010;
   45488: result <= 12'b111110000010;
   45489: result <= 12'b111110000011;
   45490: result <= 12'b111110000011;
   45491: result <= 12'b111110000011;
   45492: result <= 12'b111110000011;
   45493: result <= 12'b111110000011;
   45494: result <= 12'b111110000011;
   45495: result <= 12'b111110000011;
   45496: result <= 12'b111110000011;
   45497: result <= 12'b111110000011;
   45498: result <= 12'b111110000011;
   45499: result <= 12'b111110000011;
   45500: result <= 12'b111110000011;
   45501: result <= 12'b111110000011;
   45502: result <= 12'b111110000011;
   45503: result <= 12'b111110000011;
   45504: result <= 12'b111110000100;
   45505: result <= 12'b111110000100;
   45506: result <= 12'b111110000100;
   45507: result <= 12'b111110000100;
   45508: result <= 12'b111110000100;
   45509: result <= 12'b111110000100;
   45510: result <= 12'b111110000100;
   45511: result <= 12'b111110000100;
   45512: result <= 12'b111110000100;
   45513: result <= 12'b111110000100;
   45514: result <= 12'b111110000100;
   45515: result <= 12'b111110000100;
   45516: result <= 12'b111110000100;
   45517: result <= 12'b111110000100;
   45518: result <= 12'b111110000100;
   45519: result <= 12'b111110000101;
   45520: result <= 12'b111110000101;
   45521: result <= 12'b111110000101;
   45522: result <= 12'b111110000101;
   45523: result <= 12'b111110000101;
   45524: result <= 12'b111110000101;
   45525: result <= 12'b111110000101;
   45526: result <= 12'b111110000101;
   45527: result <= 12'b111110000101;
   45528: result <= 12'b111110000101;
   45529: result <= 12'b111110000101;
   45530: result <= 12'b111110000101;
   45531: result <= 12'b111110000101;
   45532: result <= 12'b111110000101;
   45533: result <= 12'b111110000101;
   45534: result <= 12'b111110000110;
   45535: result <= 12'b111110000110;
   45536: result <= 12'b111110000110;
   45537: result <= 12'b111110000110;
   45538: result <= 12'b111110000110;
   45539: result <= 12'b111110000110;
   45540: result <= 12'b111110000110;
   45541: result <= 12'b111110000110;
   45542: result <= 12'b111110000110;
   45543: result <= 12'b111110000110;
   45544: result <= 12'b111110000110;
   45545: result <= 12'b111110000110;
   45546: result <= 12'b111110000110;
   45547: result <= 12'b111110000110;
   45548: result <= 12'b111110000110;
   45549: result <= 12'b111110000111;
   45550: result <= 12'b111110000111;
   45551: result <= 12'b111110000111;
   45552: result <= 12'b111110000111;
   45553: result <= 12'b111110000111;
   45554: result <= 12'b111110000111;
   45555: result <= 12'b111110000111;
   45556: result <= 12'b111110000111;
   45557: result <= 12'b111110000111;
   45558: result <= 12'b111110000111;
   45559: result <= 12'b111110000111;
   45560: result <= 12'b111110000111;
   45561: result <= 12'b111110000111;
   45562: result <= 12'b111110000111;
   45563: result <= 12'b111110000111;
   45564: result <= 12'b111110001000;
   45565: result <= 12'b111110001000;
   45566: result <= 12'b111110001000;
   45567: result <= 12'b111110001000;
   45568: result <= 12'b111110001000;
   45569: result <= 12'b111110001000;
   45570: result <= 12'b111110001000;
   45571: result <= 12'b111110001000;
   45572: result <= 12'b111110001000;
   45573: result <= 12'b111110001000;
   45574: result <= 12'b111110001000;
   45575: result <= 12'b111110001000;
   45576: result <= 12'b111110001000;
   45577: result <= 12'b111110001000;
   45578: result <= 12'b111110001000;
   45579: result <= 12'b111110001001;
   45580: result <= 12'b111110001001;
   45581: result <= 12'b111110001001;
   45582: result <= 12'b111110001001;
   45583: result <= 12'b111110001001;
   45584: result <= 12'b111110001001;
   45585: result <= 12'b111110001001;
   45586: result <= 12'b111110001001;
   45587: result <= 12'b111110001001;
   45588: result <= 12'b111110001001;
   45589: result <= 12'b111110001001;
   45590: result <= 12'b111110001001;
   45591: result <= 12'b111110001001;
   45592: result <= 12'b111110001001;
   45593: result <= 12'b111110001001;
   45594: result <= 12'b111110001001;
   45595: result <= 12'b111110001010;
   45596: result <= 12'b111110001010;
   45597: result <= 12'b111110001010;
   45598: result <= 12'b111110001010;
   45599: result <= 12'b111110001010;
   45600: result <= 12'b111110001010;
   45601: result <= 12'b111110001010;
   45602: result <= 12'b111110001010;
   45603: result <= 12'b111110001010;
   45604: result <= 12'b111110001010;
   45605: result <= 12'b111110001010;
   45606: result <= 12'b111110001010;
   45607: result <= 12'b111110001010;
   45608: result <= 12'b111110001010;
   45609: result <= 12'b111110001010;
   45610: result <= 12'b111110001011;
   45611: result <= 12'b111110001011;
   45612: result <= 12'b111110001011;
   45613: result <= 12'b111110001011;
   45614: result <= 12'b111110001011;
   45615: result <= 12'b111110001011;
   45616: result <= 12'b111110001011;
   45617: result <= 12'b111110001011;
   45618: result <= 12'b111110001011;
   45619: result <= 12'b111110001011;
   45620: result <= 12'b111110001011;
   45621: result <= 12'b111110001011;
   45622: result <= 12'b111110001011;
   45623: result <= 12'b111110001011;
   45624: result <= 12'b111110001011;
   45625: result <= 12'b111110001100;
   45626: result <= 12'b111110001100;
   45627: result <= 12'b111110001100;
   45628: result <= 12'b111110001100;
   45629: result <= 12'b111110001100;
   45630: result <= 12'b111110001100;
   45631: result <= 12'b111110001100;
   45632: result <= 12'b111110001100;
   45633: result <= 12'b111110001100;
   45634: result <= 12'b111110001100;
   45635: result <= 12'b111110001100;
   45636: result <= 12'b111110001100;
   45637: result <= 12'b111110001100;
   45638: result <= 12'b111110001100;
   45639: result <= 12'b111110001100;
   45640: result <= 12'b111110001100;
   45641: result <= 12'b111110001101;
   45642: result <= 12'b111110001101;
   45643: result <= 12'b111110001101;
   45644: result <= 12'b111110001101;
   45645: result <= 12'b111110001101;
   45646: result <= 12'b111110001101;
   45647: result <= 12'b111110001101;
   45648: result <= 12'b111110001101;
   45649: result <= 12'b111110001101;
   45650: result <= 12'b111110001101;
   45651: result <= 12'b111110001101;
   45652: result <= 12'b111110001101;
   45653: result <= 12'b111110001101;
   45654: result <= 12'b111110001101;
   45655: result <= 12'b111110001101;
   45656: result <= 12'b111110001110;
   45657: result <= 12'b111110001110;
   45658: result <= 12'b111110001110;
   45659: result <= 12'b111110001110;
   45660: result <= 12'b111110001110;
   45661: result <= 12'b111110001110;
   45662: result <= 12'b111110001110;
   45663: result <= 12'b111110001110;
   45664: result <= 12'b111110001110;
   45665: result <= 12'b111110001110;
   45666: result <= 12'b111110001110;
   45667: result <= 12'b111110001110;
   45668: result <= 12'b111110001110;
   45669: result <= 12'b111110001110;
   45670: result <= 12'b111110001110;
   45671: result <= 12'b111110001111;
   45672: result <= 12'b111110001111;
   45673: result <= 12'b111110001111;
   45674: result <= 12'b111110001111;
   45675: result <= 12'b111110001111;
   45676: result <= 12'b111110001111;
   45677: result <= 12'b111110001111;
   45678: result <= 12'b111110001111;
   45679: result <= 12'b111110001111;
   45680: result <= 12'b111110001111;
   45681: result <= 12'b111110001111;
   45682: result <= 12'b111110001111;
   45683: result <= 12'b111110001111;
   45684: result <= 12'b111110001111;
   45685: result <= 12'b111110001111;
   45686: result <= 12'b111110001111;
   45687: result <= 12'b111110010000;
   45688: result <= 12'b111110010000;
   45689: result <= 12'b111110010000;
   45690: result <= 12'b111110010000;
   45691: result <= 12'b111110010000;
   45692: result <= 12'b111110010000;
   45693: result <= 12'b111110010000;
   45694: result <= 12'b111110010000;
   45695: result <= 12'b111110010000;
   45696: result <= 12'b111110010000;
   45697: result <= 12'b111110010000;
   45698: result <= 12'b111110010000;
   45699: result <= 12'b111110010000;
   45700: result <= 12'b111110010000;
   45701: result <= 12'b111110010000;
   45702: result <= 12'b111110010000;
   45703: result <= 12'b111110010001;
   45704: result <= 12'b111110010001;
   45705: result <= 12'b111110010001;
   45706: result <= 12'b111110010001;
   45707: result <= 12'b111110010001;
   45708: result <= 12'b111110010001;
   45709: result <= 12'b111110010001;
   45710: result <= 12'b111110010001;
   45711: result <= 12'b111110010001;
   45712: result <= 12'b111110010001;
   45713: result <= 12'b111110010001;
   45714: result <= 12'b111110010001;
   45715: result <= 12'b111110010001;
   45716: result <= 12'b111110010001;
   45717: result <= 12'b111110010001;
   45718: result <= 12'b111110010010;
   45719: result <= 12'b111110010010;
   45720: result <= 12'b111110010010;
   45721: result <= 12'b111110010010;
   45722: result <= 12'b111110010010;
   45723: result <= 12'b111110010010;
   45724: result <= 12'b111110010010;
   45725: result <= 12'b111110010010;
   45726: result <= 12'b111110010010;
   45727: result <= 12'b111110010010;
   45728: result <= 12'b111110010010;
   45729: result <= 12'b111110010010;
   45730: result <= 12'b111110010010;
   45731: result <= 12'b111110010010;
   45732: result <= 12'b111110010010;
   45733: result <= 12'b111110010010;
   45734: result <= 12'b111110010011;
   45735: result <= 12'b111110010011;
   45736: result <= 12'b111110010011;
   45737: result <= 12'b111110010011;
   45738: result <= 12'b111110010011;
   45739: result <= 12'b111110010011;
   45740: result <= 12'b111110010011;
   45741: result <= 12'b111110010011;
   45742: result <= 12'b111110010011;
   45743: result <= 12'b111110010011;
   45744: result <= 12'b111110010011;
   45745: result <= 12'b111110010011;
   45746: result <= 12'b111110010011;
   45747: result <= 12'b111110010011;
   45748: result <= 12'b111110010011;
   45749: result <= 12'b111110010011;
   45750: result <= 12'b111110010100;
   45751: result <= 12'b111110010100;
   45752: result <= 12'b111110010100;
   45753: result <= 12'b111110010100;
   45754: result <= 12'b111110010100;
   45755: result <= 12'b111110010100;
   45756: result <= 12'b111110010100;
   45757: result <= 12'b111110010100;
   45758: result <= 12'b111110010100;
   45759: result <= 12'b111110010100;
   45760: result <= 12'b111110010100;
   45761: result <= 12'b111110010100;
   45762: result <= 12'b111110010100;
   45763: result <= 12'b111110010100;
   45764: result <= 12'b111110010100;
   45765: result <= 12'b111110010100;
   45766: result <= 12'b111110010101;
   45767: result <= 12'b111110010101;
   45768: result <= 12'b111110010101;
   45769: result <= 12'b111110010101;
   45770: result <= 12'b111110010101;
   45771: result <= 12'b111110010101;
   45772: result <= 12'b111110010101;
   45773: result <= 12'b111110010101;
   45774: result <= 12'b111110010101;
   45775: result <= 12'b111110010101;
   45776: result <= 12'b111110010101;
   45777: result <= 12'b111110010101;
   45778: result <= 12'b111110010101;
   45779: result <= 12'b111110010101;
   45780: result <= 12'b111110010101;
   45781: result <= 12'b111110010101;
   45782: result <= 12'b111110010110;
   45783: result <= 12'b111110010110;
   45784: result <= 12'b111110010110;
   45785: result <= 12'b111110010110;
   45786: result <= 12'b111110010110;
   45787: result <= 12'b111110010110;
   45788: result <= 12'b111110010110;
   45789: result <= 12'b111110010110;
   45790: result <= 12'b111110010110;
   45791: result <= 12'b111110010110;
   45792: result <= 12'b111110010110;
   45793: result <= 12'b111110010110;
   45794: result <= 12'b111110010110;
   45795: result <= 12'b111110010110;
   45796: result <= 12'b111110010110;
   45797: result <= 12'b111110010110;
   45798: result <= 12'b111110010111;
   45799: result <= 12'b111110010111;
   45800: result <= 12'b111110010111;
   45801: result <= 12'b111110010111;
   45802: result <= 12'b111110010111;
   45803: result <= 12'b111110010111;
   45804: result <= 12'b111110010111;
   45805: result <= 12'b111110010111;
   45806: result <= 12'b111110010111;
   45807: result <= 12'b111110010111;
   45808: result <= 12'b111110010111;
   45809: result <= 12'b111110010111;
   45810: result <= 12'b111110010111;
   45811: result <= 12'b111110010111;
   45812: result <= 12'b111110010111;
   45813: result <= 12'b111110010111;
   45814: result <= 12'b111110011000;
   45815: result <= 12'b111110011000;
   45816: result <= 12'b111110011000;
   45817: result <= 12'b111110011000;
   45818: result <= 12'b111110011000;
   45819: result <= 12'b111110011000;
   45820: result <= 12'b111110011000;
   45821: result <= 12'b111110011000;
   45822: result <= 12'b111110011000;
   45823: result <= 12'b111110011000;
   45824: result <= 12'b111110011000;
   45825: result <= 12'b111110011000;
   45826: result <= 12'b111110011000;
   45827: result <= 12'b111110011000;
   45828: result <= 12'b111110011000;
   45829: result <= 12'b111110011000;
   45830: result <= 12'b111110011001;
   45831: result <= 12'b111110011001;
   45832: result <= 12'b111110011001;
   45833: result <= 12'b111110011001;
   45834: result <= 12'b111110011001;
   45835: result <= 12'b111110011001;
   45836: result <= 12'b111110011001;
   45837: result <= 12'b111110011001;
   45838: result <= 12'b111110011001;
   45839: result <= 12'b111110011001;
   45840: result <= 12'b111110011001;
   45841: result <= 12'b111110011001;
   45842: result <= 12'b111110011001;
   45843: result <= 12'b111110011001;
   45844: result <= 12'b111110011001;
   45845: result <= 12'b111110011001;
   45846: result <= 12'b111110011001;
   45847: result <= 12'b111110011010;
   45848: result <= 12'b111110011010;
   45849: result <= 12'b111110011010;
   45850: result <= 12'b111110011010;
   45851: result <= 12'b111110011010;
   45852: result <= 12'b111110011010;
   45853: result <= 12'b111110011010;
   45854: result <= 12'b111110011010;
   45855: result <= 12'b111110011010;
   45856: result <= 12'b111110011010;
   45857: result <= 12'b111110011010;
   45858: result <= 12'b111110011010;
   45859: result <= 12'b111110011010;
   45860: result <= 12'b111110011010;
   45861: result <= 12'b111110011010;
   45862: result <= 12'b111110011010;
   45863: result <= 12'b111110011011;
   45864: result <= 12'b111110011011;
   45865: result <= 12'b111110011011;
   45866: result <= 12'b111110011011;
   45867: result <= 12'b111110011011;
   45868: result <= 12'b111110011011;
   45869: result <= 12'b111110011011;
   45870: result <= 12'b111110011011;
   45871: result <= 12'b111110011011;
   45872: result <= 12'b111110011011;
   45873: result <= 12'b111110011011;
   45874: result <= 12'b111110011011;
   45875: result <= 12'b111110011011;
   45876: result <= 12'b111110011011;
   45877: result <= 12'b111110011011;
   45878: result <= 12'b111110011011;
   45879: result <= 12'b111110011011;
   45880: result <= 12'b111110011100;
   45881: result <= 12'b111110011100;
   45882: result <= 12'b111110011100;
   45883: result <= 12'b111110011100;
   45884: result <= 12'b111110011100;
   45885: result <= 12'b111110011100;
   45886: result <= 12'b111110011100;
   45887: result <= 12'b111110011100;
   45888: result <= 12'b111110011100;
   45889: result <= 12'b111110011100;
   45890: result <= 12'b111110011100;
   45891: result <= 12'b111110011100;
   45892: result <= 12'b111110011100;
   45893: result <= 12'b111110011100;
   45894: result <= 12'b111110011100;
   45895: result <= 12'b111110011100;
   45896: result <= 12'b111110011101;
   45897: result <= 12'b111110011101;
   45898: result <= 12'b111110011101;
   45899: result <= 12'b111110011101;
   45900: result <= 12'b111110011101;
   45901: result <= 12'b111110011101;
   45902: result <= 12'b111110011101;
   45903: result <= 12'b111110011101;
   45904: result <= 12'b111110011101;
   45905: result <= 12'b111110011101;
   45906: result <= 12'b111110011101;
   45907: result <= 12'b111110011101;
   45908: result <= 12'b111110011101;
   45909: result <= 12'b111110011101;
   45910: result <= 12'b111110011101;
   45911: result <= 12'b111110011101;
   45912: result <= 12'b111110011101;
   45913: result <= 12'b111110011110;
   45914: result <= 12'b111110011110;
   45915: result <= 12'b111110011110;
   45916: result <= 12'b111110011110;
   45917: result <= 12'b111110011110;
   45918: result <= 12'b111110011110;
   45919: result <= 12'b111110011110;
   45920: result <= 12'b111110011110;
   45921: result <= 12'b111110011110;
   45922: result <= 12'b111110011110;
   45923: result <= 12'b111110011110;
   45924: result <= 12'b111110011110;
   45925: result <= 12'b111110011110;
   45926: result <= 12'b111110011110;
   45927: result <= 12'b111110011110;
   45928: result <= 12'b111110011110;
   45929: result <= 12'b111110011111;
   45930: result <= 12'b111110011111;
   45931: result <= 12'b111110011111;
   45932: result <= 12'b111110011111;
   45933: result <= 12'b111110011111;
   45934: result <= 12'b111110011111;
   45935: result <= 12'b111110011111;
   45936: result <= 12'b111110011111;
   45937: result <= 12'b111110011111;
   45938: result <= 12'b111110011111;
   45939: result <= 12'b111110011111;
   45940: result <= 12'b111110011111;
   45941: result <= 12'b111110011111;
   45942: result <= 12'b111110011111;
   45943: result <= 12'b111110011111;
   45944: result <= 12'b111110011111;
   45945: result <= 12'b111110011111;
   45946: result <= 12'b111110100000;
   45947: result <= 12'b111110100000;
   45948: result <= 12'b111110100000;
   45949: result <= 12'b111110100000;
   45950: result <= 12'b111110100000;
   45951: result <= 12'b111110100000;
   45952: result <= 12'b111110100000;
   45953: result <= 12'b111110100000;
   45954: result <= 12'b111110100000;
   45955: result <= 12'b111110100000;
   45956: result <= 12'b111110100000;
   45957: result <= 12'b111110100000;
   45958: result <= 12'b111110100000;
   45959: result <= 12'b111110100000;
   45960: result <= 12'b111110100000;
   45961: result <= 12'b111110100000;
   45962: result <= 12'b111110100000;
   45963: result <= 12'b111110100001;
   45964: result <= 12'b111110100001;
   45965: result <= 12'b111110100001;
   45966: result <= 12'b111110100001;
   45967: result <= 12'b111110100001;
   45968: result <= 12'b111110100001;
   45969: result <= 12'b111110100001;
   45970: result <= 12'b111110100001;
   45971: result <= 12'b111110100001;
   45972: result <= 12'b111110100001;
   45973: result <= 12'b111110100001;
   45974: result <= 12'b111110100001;
   45975: result <= 12'b111110100001;
   45976: result <= 12'b111110100001;
   45977: result <= 12'b111110100001;
   45978: result <= 12'b111110100001;
   45979: result <= 12'b111110100001;
   45980: result <= 12'b111110100010;
   45981: result <= 12'b111110100010;
   45982: result <= 12'b111110100010;
   45983: result <= 12'b111110100010;
   45984: result <= 12'b111110100010;
   45985: result <= 12'b111110100010;
   45986: result <= 12'b111110100010;
   45987: result <= 12'b111110100010;
   45988: result <= 12'b111110100010;
   45989: result <= 12'b111110100010;
   45990: result <= 12'b111110100010;
   45991: result <= 12'b111110100010;
   45992: result <= 12'b111110100010;
   45993: result <= 12'b111110100010;
   45994: result <= 12'b111110100010;
   45995: result <= 12'b111110100010;
   45996: result <= 12'b111110100010;
   45997: result <= 12'b111110100011;
   45998: result <= 12'b111110100011;
   45999: result <= 12'b111110100011;
   46000: result <= 12'b111110100011;
   46001: result <= 12'b111110100011;
   46002: result <= 12'b111110100011;
   46003: result <= 12'b111110100011;
   46004: result <= 12'b111110100011;
   46005: result <= 12'b111110100011;
   46006: result <= 12'b111110100011;
   46007: result <= 12'b111110100011;
   46008: result <= 12'b111110100011;
   46009: result <= 12'b111110100011;
   46010: result <= 12'b111110100011;
   46011: result <= 12'b111110100011;
   46012: result <= 12'b111110100011;
   46013: result <= 12'b111110100011;
   46014: result <= 12'b111110100100;
   46015: result <= 12'b111110100100;
   46016: result <= 12'b111110100100;
   46017: result <= 12'b111110100100;
   46018: result <= 12'b111110100100;
   46019: result <= 12'b111110100100;
   46020: result <= 12'b111110100100;
   46021: result <= 12'b111110100100;
   46022: result <= 12'b111110100100;
   46023: result <= 12'b111110100100;
   46024: result <= 12'b111110100100;
   46025: result <= 12'b111110100100;
   46026: result <= 12'b111110100100;
   46027: result <= 12'b111110100100;
   46028: result <= 12'b111110100100;
   46029: result <= 12'b111110100100;
   46030: result <= 12'b111110100100;
   46031: result <= 12'b111110100100;
   46032: result <= 12'b111110100101;
   46033: result <= 12'b111110100101;
   46034: result <= 12'b111110100101;
   46035: result <= 12'b111110100101;
   46036: result <= 12'b111110100101;
   46037: result <= 12'b111110100101;
   46038: result <= 12'b111110100101;
   46039: result <= 12'b111110100101;
   46040: result <= 12'b111110100101;
   46041: result <= 12'b111110100101;
   46042: result <= 12'b111110100101;
   46043: result <= 12'b111110100101;
   46044: result <= 12'b111110100101;
   46045: result <= 12'b111110100101;
   46046: result <= 12'b111110100101;
   46047: result <= 12'b111110100101;
   46048: result <= 12'b111110100101;
   46049: result <= 12'b111110100110;
   46050: result <= 12'b111110100110;
   46051: result <= 12'b111110100110;
   46052: result <= 12'b111110100110;
   46053: result <= 12'b111110100110;
   46054: result <= 12'b111110100110;
   46055: result <= 12'b111110100110;
   46056: result <= 12'b111110100110;
   46057: result <= 12'b111110100110;
   46058: result <= 12'b111110100110;
   46059: result <= 12'b111110100110;
   46060: result <= 12'b111110100110;
   46061: result <= 12'b111110100110;
   46062: result <= 12'b111110100110;
   46063: result <= 12'b111110100110;
   46064: result <= 12'b111110100110;
   46065: result <= 12'b111110100110;
   46066: result <= 12'b111110100111;
   46067: result <= 12'b111110100111;
   46068: result <= 12'b111110100111;
   46069: result <= 12'b111110100111;
   46070: result <= 12'b111110100111;
   46071: result <= 12'b111110100111;
   46072: result <= 12'b111110100111;
   46073: result <= 12'b111110100111;
   46074: result <= 12'b111110100111;
   46075: result <= 12'b111110100111;
   46076: result <= 12'b111110100111;
   46077: result <= 12'b111110100111;
   46078: result <= 12'b111110100111;
   46079: result <= 12'b111110100111;
   46080: result <= 12'b111110100111;
   46081: result <= 12'b111110100111;
   46082: result <= 12'b111110100111;
   46083: result <= 12'b111110100111;
   46084: result <= 12'b111110101000;
   46085: result <= 12'b111110101000;
   46086: result <= 12'b111110101000;
   46087: result <= 12'b111110101000;
   46088: result <= 12'b111110101000;
   46089: result <= 12'b111110101000;
   46090: result <= 12'b111110101000;
   46091: result <= 12'b111110101000;
   46092: result <= 12'b111110101000;
   46093: result <= 12'b111110101000;
   46094: result <= 12'b111110101000;
   46095: result <= 12'b111110101000;
   46096: result <= 12'b111110101000;
   46097: result <= 12'b111110101000;
   46098: result <= 12'b111110101000;
   46099: result <= 12'b111110101000;
   46100: result <= 12'b111110101000;
   46101: result <= 12'b111110101001;
   46102: result <= 12'b111110101001;
   46103: result <= 12'b111110101001;
   46104: result <= 12'b111110101001;
   46105: result <= 12'b111110101001;
   46106: result <= 12'b111110101001;
   46107: result <= 12'b111110101001;
   46108: result <= 12'b111110101001;
   46109: result <= 12'b111110101001;
   46110: result <= 12'b111110101001;
   46111: result <= 12'b111110101001;
   46112: result <= 12'b111110101001;
   46113: result <= 12'b111110101001;
   46114: result <= 12'b111110101001;
   46115: result <= 12'b111110101001;
   46116: result <= 12'b111110101001;
   46117: result <= 12'b111110101001;
   46118: result <= 12'b111110101001;
   46119: result <= 12'b111110101010;
   46120: result <= 12'b111110101010;
   46121: result <= 12'b111110101010;
   46122: result <= 12'b111110101010;
   46123: result <= 12'b111110101010;
   46124: result <= 12'b111110101010;
   46125: result <= 12'b111110101010;
   46126: result <= 12'b111110101010;
   46127: result <= 12'b111110101010;
   46128: result <= 12'b111110101010;
   46129: result <= 12'b111110101010;
   46130: result <= 12'b111110101010;
   46131: result <= 12'b111110101010;
   46132: result <= 12'b111110101010;
   46133: result <= 12'b111110101010;
   46134: result <= 12'b111110101010;
   46135: result <= 12'b111110101010;
   46136: result <= 12'b111110101010;
   46137: result <= 12'b111110101011;
   46138: result <= 12'b111110101011;
   46139: result <= 12'b111110101011;
   46140: result <= 12'b111110101011;
   46141: result <= 12'b111110101011;
   46142: result <= 12'b111110101011;
   46143: result <= 12'b111110101011;
   46144: result <= 12'b111110101011;
   46145: result <= 12'b111110101011;
   46146: result <= 12'b111110101011;
   46147: result <= 12'b111110101011;
   46148: result <= 12'b111110101011;
   46149: result <= 12'b111110101011;
   46150: result <= 12'b111110101011;
   46151: result <= 12'b111110101011;
   46152: result <= 12'b111110101011;
   46153: result <= 12'b111110101011;
   46154: result <= 12'b111110101011;
   46155: result <= 12'b111110101100;
   46156: result <= 12'b111110101100;
   46157: result <= 12'b111110101100;
   46158: result <= 12'b111110101100;
   46159: result <= 12'b111110101100;
   46160: result <= 12'b111110101100;
   46161: result <= 12'b111110101100;
   46162: result <= 12'b111110101100;
   46163: result <= 12'b111110101100;
   46164: result <= 12'b111110101100;
   46165: result <= 12'b111110101100;
   46166: result <= 12'b111110101100;
   46167: result <= 12'b111110101100;
   46168: result <= 12'b111110101100;
   46169: result <= 12'b111110101100;
   46170: result <= 12'b111110101100;
   46171: result <= 12'b111110101100;
   46172: result <= 12'b111110101100;
   46173: result <= 12'b111110101101;
   46174: result <= 12'b111110101101;
   46175: result <= 12'b111110101101;
   46176: result <= 12'b111110101101;
   46177: result <= 12'b111110101101;
   46178: result <= 12'b111110101101;
   46179: result <= 12'b111110101101;
   46180: result <= 12'b111110101101;
   46181: result <= 12'b111110101101;
   46182: result <= 12'b111110101101;
   46183: result <= 12'b111110101101;
   46184: result <= 12'b111110101101;
   46185: result <= 12'b111110101101;
   46186: result <= 12'b111110101101;
   46187: result <= 12'b111110101101;
   46188: result <= 12'b111110101101;
   46189: result <= 12'b111110101101;
   46190: result <= 12'b111110101101;
   46191: result <= 12'b111110101110;
   46192: result <= 12'b111110101110;
   46193: result <= 12'b111110101110;
   46194: result <= 12'b111110101110;
   46195: result <= 12'b111110101110;
   46196: result <= 12'b111110101110;
   46197: result <= 12'b111110101110;
   46198: result <= 12'b111110101110;
   46199: result <= 12'b111110101110;
   46200: result <= 12'b111110101110;
   46201: result <= 12'b111110101110;
   46202: result <= 12'b111110101110;
   46203: result <= 12'b111110101110;
   46204: result <= 12'b111110101110;
   46205: result <= 12'b111110101110;
   46206: result <= 12'b111110101110;
   46207: result <= 12'b111110101110;
   46208: result <= 12'b111110101110;
   46209: result <= 12'b111110101111;
   46210: result <= 12'b111110101111;
   46211: result <= 12'b111110101111;
   46212: result <= 12'b111110101111;
   46213: result <= 12'b111110101111;
   46214: result <= 12'b111110101111;
   46215: result <= 12'b111110101111;
   46216: result <= 12'b111110101111;
   46217: result <= 12'b111110101111;
   46218: result <= 12'b111110101111;
   46219: result <= 12'b111110101111;
   46220: result <= 12'b111110101111;
   46221: result <= 12'b111110101111;
   46222: result <= 12'b111110101111;
   46223: result <= 12'b111110101111;
   46224: result <= 12'b111110101111;
   46225: result <= 12'b111110101111;
   46226: result <= 12'b111110101111;
   46227: result <= 12'b111110101111;
   46228: result <= 12'b111110110000;
   46229: result <= 12'b111110110000;
   46230: result <= 12'b111110110000;
   46231: result <= 12'b111110110000;
   46232: result <= 12'b111110110000;
   46233: result <= 12'b111110110000;
   46234: result <= 12'b111110110000;
   46235: result <= 12'b111110110000;
   46236: result <= 12'b111110110000;
   46237: result <= 12'b111110110000;
   46238: result <= 12'b111110110000;
   46239: result <= 12'b111110110000;
   46240: result <= 12'b111110110000;
   46241: result <= 12'b111110110000;
   46242: result <= 12'b111110110000;
   46243: result <= 12'b111110110000;
   46244: result <= 12'b111110110000;
   46245: result <= 12'b111110110000;
   46246: result <= 12'b111110110001;
   46247: result <= 12'b111110110001;
   46248: result <= 12'b111110110001;
   46249: result <= 12'b111110110001;
   46250: result <= 12'b111110110001;
   46251: result <= 12'b111110110001;
   46252: result <= 12'b111110110001;
   46253: result <= 12'b111110110001;
   46254: result <= 12'b111110110001;
   46255: result <= 12'b111110110001;
   46256: result <= 12'b111110110001;
   46257: result <= 12'b111110110001;
   46258: result <= 12'b111110110001;
   46259: result <= 12'b111110110001;
   46260: result <= 12'b111110110001;
   46261: result <= 12'b111110110001;
   46262: result <= 12'b111110110001;
   46263: result <= 12'b111110110001;
   46264: result <= 12'b111110110001;
   46265: result <= 12'b111110110010;
   46266: result <= 12'b111110110010;
   46267: result <= 12'b111110110010;
   46268: result <= 12'b111110110010;
   46269: result <= 12'b111110110010;
   46270: result <= 12'b111110110010;
   46271: result <= 12'b111110110010;
   46272: result <= 12'b111110110010;
   46273: result <= 12'b111110110010;
   46274: result <= 12'b111110110010;
   46275: result <= 12'b111110110010;
   46276: result <= 12'b111110110010;
   46277: result <= 12'b111110110010;
   46278: result <= 12'b111110110010;
   46279: result <= 12'b111110110010;
   46280: result <= 12'b111110110010;
   46281: result <= 12'b111110110010;
   46282: result <= 12'b111110110010;
   46283: result <= 12'b111110110011;
   46284: result <= 12'b111110110011;
   46285: result <= 12'b111110110011;
   46286: result <= 12'b111110110011;
   46287: result <= 12'b111110110011;
   46288: result <= 12'b111110110011;
   46289: result <= 12'b111110110011;
   46290: result <= 12'b111110110011;
   46291: result <= 12'b111110110011;
   46292: result <= 12'b111110110011;
   46293: result <= 12'b111110110011;
   46294: result <= 12'b111110110011;
   46295: result <= 12'b111110110011;
   46296: result <= 12'b111110110011;
   46297: result <= 12'b111110110011;
   46298: result <= 12'b111110110011;
   46299: result <= 12'b111110110011;
   46300: result <= 12'b111110110011;
   46301: result <= 12'b111110110011;
   46302: result <= 12'b111110110100;
   46303: result <= 12'b111110110100;
   46304: result <= 12'b111110110100;
   46305: result <= 12'b111110110100;
   46306: result <= 12'b111110110100;
   46307: result <= 12'b111110110100;
   46308: result <= 12'b111110110100;
   46309: result <= 12'b111110110100;
   46310: result <= 12'b111110110100;
   46311: result <= 12'b111110110100;
   46312: result <= 12'b111110110100;
   46313: result <= 12'b111110110100;
   46314: result <= 12'b111110110100;
   46315: result <= 12'b111110110100;
   46316: result <= 12'b111110110100;
   46317: result <= 12'b111110110100;
   46318: result <= 12'b111110110100;
   46319: result <= 12'b111110110100;
   46320: result <= 12'b111110110100;
   46321: result <= 12'b111110110101;
   46322: result <= 12'b111110110101;
   46323: result <= 12'b111110110101;
   46324: result <= 12'b111110110101;
   46325: result <= 12'b111110110101;
   46326: result <= 12'b111110110101;
   46327: result <= 12'b111110110101;
   46328: result <= 12'b111110110101;
   46329: result <= 12'b111110110101;
   46330: result <= 12'b111110110101;
   46331: result <= 12'b111110110101;
   46332: result <= 12'b111110110101;
   46333: result <= 12'b111110110101;
   46334: result <= 12'b111110110101;
   46335: result <= 12'b111110110101;
   46336: result <= 12'b111110110101;
   46337: result <= 12'b111110110101;
   46338: result <= 12'b111110110101;
   46339: result <= 12'b111110110101;
   46340: result <= 12'b111110110110;
   46341: result <= 12'b111110110110;
   46342: result <= 12'b111110110110;
   46343: result <= 12'b111110110110;
   46344: result <= 12'b111110110110;
   46345: result <= 12'b111110110110;
   46346: result <= 12'b111110110110;
   46347: result <= 12'b111110110110;
   46348: result <= 12'b111110110110;
   46349: result <= 12'b111110110110;
   46350: result <= 12'b111110110110;
   46351: result <= 12'b111110110110;
   46352: result <= 12'b111110110110;
   46353: result <= 12'b111110110110;
   46354: result <= 12'b111110110110;
   46355: result <= 12'b111110110110;
   46356: result <= 12'b111110110110;
   46357: result <= 12'b111110110110;
   46358: result <= 12'b111110110110;
   46359: result <= 12'b111110110111;
   46360: result <= 12'b111110110111;
   46361: result <= 12'b111110110111;
   46362: result <= 12'b111110110111;
   46363: result <= 12'b111110110111;
   46364: result <= 12'b111110110111;
   46365: result <= 12'b111110110111;
   46366: result <= 12'b111110110111;
   46367: result <= 12'b111110110111;
   46368: result <= 12'b111110110111;
   46369: result <= 12'b111110110111;
   46370: result <= 12'b111110110111;
   46371: result <= 12'b111110110111;
   46372: result <= 12'b111110110111;
   46373: result <= 12'b111110110111;
   46374: result <= 12'b111110110111;
   46375: result <= 12'b111110110111;
   46376: result <= 12'b111110110111;
   46377: result <= 12'b111110110111;
   46378: result <= 12'b111110110111;
   46379: result <= 12'b111110111000;
   46380: result <= 12'b111110111000;
   46381: result <= 12'b111110111000;
   46382: result <= 12'b111110111000;
   46383: result <= 12'b111110111000;
   46384: result <= 12'b111110111000;
   46385: result <= 12'b111110111000;
   46386: result <= 12'b111110111000;
   46387: result <= 12'b111110111000;
   46388: result <= 12'b111110111000;
   46389: result <= 12'b111110111000;
   46390: result <= 12'b111110111000;
   46391: result <= 12'b111110111000;
   46392: result <= 12'b111110111000;
   46393: result <= 12'b111110111000;
   46394: result <= 12'b111110111000;
   46395: result <= 12'b111110111000;
   46396: result <= 12'b111110111000;
   46397: result <= 12'b111110111000;
   46398: result <= 12'b111110111001;
   46399: result <= 12'b111110111001;
   46400: result <= 12'b111110111001;
   46401: result <= 12'b111110111001;
   46402: result <= 12'b111110111001;
   46403: result <= 12'b111110111001;
   46404: result <= 12'b111110111001;
   46405: result <= 12'b111110111001;
   46406: result <= 12'b111110111001;
   46407: result <= 12'b111110111001;
   46408: result <= 12'b111110111001;
   46409: result <= 12'b111110111001;
   46410: result <= 12'b111110111001;
   46411: result <= 12'b111110111001;
   46412: result <= 12'b111110111001;
   46413: result <= 12'b111110111001;
   46414: result <= 12'b111110111001;
   46415: result <= 12'b111110111001;
   46416: result <= 12'b111110111001;
   46417: result <= 12'b111110111001;
   46418: result <= 12'b111110111010;
   46419: result <= 12'b111110111010;
   46420: result <= 12'b111110111010;
   46421: result <= 12'b111110111010;
   46422: result <= 12'b111110111010;
   46423: result <= 12'b111110111010;
   46424: result <= 12'b111110111010;
   46425: result <= 12'b111110111010;
   46426: result <= 12'b111110111010;
   46427: result <= 12'b111110111010;
   46428: result <= 12'b111110111010;
   46429: result <= 12'b111110111010;
   46430: result <= 12'b111110111010;
   46431: result <= 12'b111110111010;
   46432: result <= 12'b111110111010;
   46433: result <= 12'b111110111010;
   46434: result <= 12'b111110111010;
   46435: result <= 12'b111110111010;
   46436: result <= 12'b111110111010;
   46437: result <= 12'b111110111011;
   46438: result <= 12'b111110111011;
   46439: result <= 12'b111110111011;
   46440: result <= 12'b111110111011;
   46441: result <= 12'b111110111011;
   46442: result <= 12'b111110111011;
   46443: result <= 12'b111110111011;
   46444: result <= 12'b111110111011;
   46445: result <= 12'b111110111011;
   46446: result <= 12'b111110111011;
   46447: result <= 12'b111110111011;
   46448: result <= 12'b111110111011;
   46449: result <= 12'b111110111011;
   46450: result <= 12'b111110111011;
   46451: result <= 12'b111110111011;
   46452: result <= 12'b111110111011;
   46453: result <= 12'b111110111011;
   46454: result <= 12'b111110111011;
   46455: result <= 12'b111110111011;
   46456: result <= 12'b111110111011;
   46457: result <= 12'b111110111100;
   46458: result <= 12'b111110111100;
   46459: result <= 12'b111110111100;
   46460: result <= 12'b111110111100;
   46461: result <= 12'b111110111100;
   46462: result <= 12'b111110111100;
   46463: result <= 12'b111110111100;
   46464: result <= 12'b111110111100;
   46465: result <= 12'b111110111100;
   46466: result <= 12'b111110111100;
   46467: result <= 12'b111110111100;
   46468: result <= 12'b111110111100;
   46469: result <= 12'b111110111100;
   46470: result <= 12'b111110111100;
   46471: result <= 12'b111110111100;
   46472: result <= 12'b111110111100;
   46473: result <= 12'b111110111100;
   46474: result <= 12'b111110111100;
   46475: result <= 12'b111110111100;
   46476: result <= 12'b111110111100;
   46477: result <= 12'b111110111101;
   46478: result <= 12'b111110111101;
   46479: result <= 12'b111110111101;
   46480: result <= 12'b111110111101;
   46481: result <= 12'b111110111101;
   46482: result <= 12'b111110111101;
   46483: result <= 12'b111110111101;
   46484: result <= 12'b111110111101;
   46485: result <= 12'b111110111101;
   46486: result <= 12'b111110111101;
   46487: result <= 12'b111110111101;
   46488: result <= 12'b111110111101;
   46489: result <= 12'b111110111101;
   46490: result <= 12'b111110111101;
   46491: result <= 12'b111110111101;
   46492: result <= 12'b111110111101;
   46493: result <= 12'b111110111101;
   46494: result <= 12'b111110111101;
   46495: result <= 12'b111110111101;
   46496: result <= 12'b111110111101;
   46497: result <= 12'b111110111110;
   46498: result <= 12'b111110111110;
   46499: result <= 12'b111110111110;
   46500: result <= 12'b111110111110;
   46501: result <= 12'b111110111110;
   46502: result <= 12'b111110111110;
   46503: result <= 12'b111110111110;
   46504: result <= 12'b111110111110;
   46505: result <= 12'b111110111110;
   46506: result <= 12'b111110111110;
   46507: result <= 12'b111110111110;
   46508: result <= 12'b111110111110;
   46509: result <= 12'b111110111110;
   46510: result <= 12'b111110111110;
   46511: result <= 12'b111110111110;
   46512: result <= 12'b111110111110;
   46513: result <= 12'b111110111110;
   46514: result <= 12'b111110111110;
   46515: result <= 12'b111110111110;
   46516: result <= 12'b111110111110;
   46517: result <= 12'b111110111110;
   46518: result <= 12'b111110111111;
   46519: result <= 12'b111110111111;
   46520: result <= 12'b111110111111;
   46521: result <= 12'b111110111111;
   46522: result <= 12'b111110111111;
   46523: result <= 12'b111110111111;
   46524: result <= 12'b111110111111;
   46525: result <= 12'b111110111111;
   46526: result <= 12'b111110111111;
   46527: result <= 12'b111110111111;
   46528: result <= 12'b111110111111;
   46529: result <= 12'b111110111111;
   46530: result <= 12'b111110111111;
   46531: result <= 12'b111110111111;
   46532: result <= 12'b111110111111;
   46533: result <= 12'b111110111111;
   46534: result <= 12'b111110111111;
   46535: result <= 12'b111110111111;
   46536: result <= 12'b111110111111;
   46537: result <= 12'b111110111111;
   46538: result <= 12'b111111000000;
   46539: result <= 12'b111111000000;
   46540: result <= 12'b111111000000;
   46541: result <= 12'b111111000000;
   46542: result <= 12'b111111000000;
   46543: result <= 12'b111111000000;
   46544: result <= 12'b111111000000;
   46545: result <= 12'b111111000000;
   46546: result <= 12'b111111000000;
   46547: result <= 12'b111111000000;
   46548: result <= 12'b111111000000;
   46549: result <= 12'b111111000000;
   46550: result <= 12'b111111000000;
   46551: result <= 12'b111111000000;
   46552: result <= 12'b111111000000;
   46553: result <= 12'b111111000000;
   46554: result <= 12'b111111000000;
   46555: result <= 12'b111111000000;
   46556: result <= 12'b111111000000;
   46557: result <= 12'b111111000000;
   46558: result <= 12'b111111000000;
   46559: result <= 12'b111111000001;
   46560: result <= 12'b111111000001;
   46561: result <= 12'b111111000001;
   46562: result <= 12'b111111000001;
   46563: result <= 12'b111111000001;
   46564: result <= 12'b111111000001;
   46565: result <= 12'b111111000001;
   46566: result <= 12'b111111000001;
   46567: result <= 12'b111111000001;
   46568: result <= 12'b111111000001;
   46569: result <= 12'b111111000001;
   46570: result <= 12'b111111000001;
   46571: result <= 12'b111111000001;
   46572: result <= 12'b111111000001;
   46573: result <= 12'b111111000001;
   46574: result <= 12'b111111000001;
   46575: result <= 12'b111111000001;
   46576: result <= 12'b111111000001;
   46577: result <= 12'b111111000001;
   46578: result <= 12'b111111000001;
   46579: result <= 12'b111111000010;
   46580: result <= 12'b111111000010;
   46581: result <= 12'b111111000010;
   46582: result <= 12'b111111000010;
   46583: result <= 12'b111111000010;
   46584: result <= 12'b111111000010;
   46585: result <= 12'b111111000010;
   46586: result <= 12'b111111000010;
   46587: result <= 12'b111111000010;
   46588: result <= 12'b111111000010;
   46589: result <= 12'b111111000010;
   46590: result <= 12'b111111000010;
   46591: result <= 12'b111111000010;
   46592: result <= 12'b111111000010;
   46593: result <= 12'b111111000010;
   46594: result <= 12'b111111000010;
   46595: result <= 12'b111111000010;
   46596: result <= 12'b111111000010;
   46597: result <= 12'b111111000010;
   46598: result <= 12'b111111000010;
   46599: result <= 12'b111111000010;
   46600: result <= 12'b111111000011;
   46601: result <= 12'b111111000011;
   46602: result <= 12'b111111000011;
   46603: result <= 12'b111111000011;
   46604: result <= 12'b111111000011;
   46605: result <= 12'b111111000011;
   46606: result <= 12'b111111000011;
   46607: result <= 12'b111111000011;
   46608: result <= 12'b111111000011;
   46609: result <= 12'b111111000011;
   46610: result <= 12'b111111000011;
   46611: result <= 12'b111111000011;
   46612: result <= 12'b111111000011;
   46613: result <= 12'b111111000011;
   46614: result <= 12'b111111000011;
   46615: result <= 12'b111111000011;
   46616: result <= 12'b111111000011;
   46617: result <= 12'b111111000011;
   46618: result <= 12'b111111000011;
   46619: result <= 12'b111111000011;
   46620: result <= 12'b111111000011;
   46621: result <= 12'b111111000011;
   46622: result <= 12'b111111000100;
   46623: result <= 12'b111111000100;
   46624: result <= 12'b111111000100;
   46625: result <= 12'b111111000100;
   46626: result <= 12'b111111000100;
   46627: result <= 12'b111111000100;
   46628: result <= 12'b111111000100;
   46629: result <= 12'b111111000100;
   46630: result <= 12'b111111000100;
   46631: result <= 12'b111111000100;
   46632: result <= 12'b111111000100;
   46633: result <= 12'b111111000100;
   46634: result <= 12'b111111000100;
   46635: result <= 12'b111111000100;
   46636: result <= 12'b111111000100;
   46637: result <= 12'b111111000100;
   46638: result <= 12'b111111000100;
   46639: result <= 12'b111111000100;
   46640: result <= 12'b111111000100;
   46641: result <= 12'b111111000100;
   46642: result <= 12'b111111000100;
   46643: result <= 12'b111111000101;
   46644: result <= 12'b111111000101;
   46645: result <= 12'b111111000101;
   46646: result <= 12'b111111000101;
   46647: result <= 12'b111111000101;
   46648: result <= 12'b111111000101;
   46649: result <= 12'b111111000101;
   46650: result <= 12'b111111000101;
   46651: result <= 12'b111111000101;
   46652: result <= 12'b111111000101;
   46653: result <= 12'b111111000101;
   46654: result <= 12'b111111000101;
   46655: result <= 12'b111111000101;
   46656: result <= 12'b111111000101;
   46657: result <= 12'b111111000101;
   46658: result <= 12'b111111000101;
   46659: result <= 12'b111111000101;
   46660: result <= 12'b111111000101;
   46661: result <= 12'b111111000101;
   46662: result <= 12'b111111000101;
   46663: result <= 12'b111111000101;
   46664: result <= 12'b111111000110;
   46665: result <= 12'b111111000110;
   46666: result <= 12'b111111000110;
   46667: result <= 12'b111111000110;
   46668: result <= 12'b111111000110;
   46669: result <= 12'b111111000110;
   46670: result <= 12'b111111000110;
   46671: result <= 12'b111111000110;
   46672: result <= 12'b111111000110;
   46673: result <= 12'b111111000110;
   46674: result <= 12'b111111000110;
   46675: result <= 12'b111111000110;
   46676: result <= 12'b111111000110;
   46677: result <= 12'b111111000110;
   46678: result <= 12'b111111000110;
   46679: result <= 12'b111111000110;
   46680: result <= 12'b111111000110;
   46681: result <= 12'b111111000110;
   46682: result <= 12'b111111000110;
   46683: result <= 12'b111111000110;
   46684: result <= 12'b111111000110;
   46685: result <= 12'b111111000110;
   46686: result <= 12'b111111000111;
   46687: result <= 12'b111111000111;
   46688: result <= 12'b111111000111;
   46689: result <= 12'b111111000111;
   46690: result <= 12'b111111000111;
   46691: result <= 12'b111111000111;
   46692: result <= 12'b111111000111;
   46693: result <= 12'b111111000111;
   46694: result <= 12'b111111000111;
   46695: result <= 12'b111111000111;
   46696: result <= 12'b111111000111;
   46697: result <= 12'b111111000111;
   46698: result <= 12'b111111000111;
   46699: result <= 12'b111111000111;
   46700: result <= 12'b111111000111;
   46701: result <= 12'b111111000111;
   46702: result <= 12'b111111000111;
   46703: result <= 12'b111111000111;
   46704: result <= 12'b111111000111;
   46705: result <= 12'b111111000111;
   46706: result <= 12'b111111000111;
   46707: result <= 12'b111111000111;
   46708: result <= 12'b111111001000;
   46709: result <= 12'b111111001000;
   46710: result <= 12'b111111001000;
   46711: result <= 12'b111111001000;
   46712: result <= 12'b111111001000;
   46713: result <= 12'b111111001000;
   46714: result <= 12'b111111001000;
   46715: result <= 12'b111111001000;
   46716: result <= 12'b111111001000;
   46717: result <= 12'b111111001000;
   46718: result <= 12'b111111001000;
   46719: result <= 12'b111111001000;
   46720: result <= 12'b111111001000;
   46721: result <= 12'b111111001000;
   46722: result <= 12'b111111001000;
   46723: result <= 12'b111111001000;
   46724: result <= 12'b111111001000;
   46725: result <= 12'b111111001000;
   46726: result <= 12'b111111001000;
   46727: result <= 12'b111111001000;
   46728: result <= 12'b111111001000;
   46729: result <= 12'b111111001000;
   46730: result <= 12'b111111001001;
   46731: result <= 12'b111111001001;
   46732: result <= 12'b111111001001;
   46733: result <= 12'b111111001001;
   46734: result <= 12'b111111001001;
   46735: result <= 12'b111111001001;
   46736: result <= 12'b111111001001;
   46737: result <= 12'b111111001001;
   46738: result <= 12'b111111001001;
   46739: result <= 12'b111111001001;
   46740: result <= 12'b111111001001;
   46741: result <= 12'b111111001001;
   46742: result <= 12'b111111001001;
   46743: result <= 12'b111111001001;
   46744: result <= 12'b111111001001;
   46745: result <= 12'b111111001001;
   46746: result <= 12'b111111001001;
   46747: result <= 12'b111111001001;
   46748: result <= 12'b111111001001;
   46749: result <= 12'b111111001001;
   46750: result <= 12'b111111001001;
   46751: result <= 12'b111111001001;
   46752: result <= 12'b111111001010;
   46753: result <= 12'b111111001010;
   46754: result <= 12'b111111001010;
   46755: result <= 12'b111111001010;
   46756: result <= 12'b111111001010;
   46757: result <= 12'b111111001010;
   46758: result <= 12'b111111001010;
   46759: result <= 12'b111111001010;
   46760: result <= 12'b111111001010;
   46761: result <= 12'b111111001010;
   46762: result <= 12'b111111001010;
   46763: result <= 12'b111111001010;
   46764: result <= 12'b111111001010;
   46765: result <= 12'b111111001010;
   46766: result <= 12'b111111001010;
   46767: result <= 12'b111111001010;
   46768: result <= 12'b111111001010;
   46769: result <= 12'b111111001010;
   46770: result <= 12'b111111001010;
   46771: result <= 12'b111111001010;
   46772: result <= 12'b111111001010;
   46773: result <= 12'b111111001010;
   46774: result <= 12'b111111001011;
   46775: result <= 12'b111111001011;
   46776: result <= 12'b111111001011;
   46777: result <= 12'b111111001011;
   46778: result <= 12'b111111001011;
   46779: result <= 12'b111111001011;
   46780: result <= 12'b111111001011;
   46781: result <= 12'b111111001011;
   46782: result <= 12'b111111001011;
   46783: result <= 12'b111111001011;
   46784: result <= 12'b111111001011;
   46785: result <= 12'b111111001011;
   46786: result <= 12'b111111001011;
   46787: result <= 12'b111111001011;
   46788: result <= 12'b111111001011;
   46789: result <= 12'b111111001011;
   46790: result <= 12'b111111001011;
   46791: result <= 12'b111111001011;
   46792: result <= 12'b111111001011;
   46793: result <= 12'b111111001011;
   46794: result <= 12'b111111001011;
   46795: result <= 12'b111111001011;
   46796: result <= 12'b111111001011;
   46797: result <= 12'b111111001100;
   46798: result <= 12'b111111001100;
   46799: result <= 12'b111111001100;
   46800: result <= 12'b111111001100;
   46801: result <= 12'b111111001100;
   46802: result <= 12'b111111001100;
   46803: result <= 12'b111111001100;
   46804: result <= 12'b111111001100;
   46805: result <= 12'b111111001100;
   46806: result <= 12'b111111001100;
   46807: result <= 12'b111111001100;
   46808: result <= 12'b111111001100;
   46809: result <= 12'b111111001100;
   46810: result <= 12'b111111001100;
   46811: result <= 12'b111111001100;
   46812: result <= 12'b111111001100;
   46813: result <= 12'b111111001100;
   46814: result <= 12'b111111001100;
   46815: result <= 12'b111111001100;
   46816: result <= 12'b111111001100;
   46817: result <= 12'b111111001100;
   46818: result <= 12'b111111001100;
   46819: result <= 12'b111111001100;
   46820: result <= 12'b111111001101;
   46821: result <= 12'b111111001101;
   46822: result <= 12'b111111001101;
   46823: result <= 12'b111111001101;
   46824: result <= 12'b111111001101;
   46825: result <= 12'b111111001101;
   46826: result <= 12'b111111001101;
   46827: result <= 12'b111111001101;
   46828: result <= 12'b111111001101;
   46829: result <= 12'b111111001101;
   46830: result <= 12'b111111001101;
   46831: result <= 12'b111111001101;
   46832: result <= 12'b111111001101;
   46833: result <= 12'b111111001101;
   46834: result <= 12'b111111001101;
   46835: result <= 12'b111111001101;
   46836: result <= 12'b111111001101;
   46837: result <= 12'b111111001101;
   46838: result <= 12'b111111001101;
   46839: result <= 12'b111111001101;
   46840: result <= 12'b111111001101;
   46841: result <= 12'b111111001101;
   46842: result <= 12'b111111001101;
   46843: result <= 12'b111111001110;
   46844: result <= 12'b111111001110;
   46845: result <= 12'b111111001110;
   46846: result <= 12'b111111001110;
   46847: result <= 12'b111111001110;
   46848: result <= 12'b111111001110;
   46849: result <= 12'b111111001110;
   46850: result <= 12'b111111001110;
   46851: result <= 12'b111111001110;
   46852: result <= 12'b111111001110;
   46853: result <= 12'b111111001110;
   46854: result <= 12'b111111001110;
   46855: result <= 12'b111111001110;
   46856: result <= 12'b111111001110;
   46857: result <= 12'b111111001110;
   46858: result <= 12'b111111001110;
   46859: result <= 12'b111111001110;
   46860: result <= 12'b111111001110;
   46861: result <= 12'b111111001110;
   46862: result <= 12'b111111001110;
   46863: result <= 12'b111111001110;
   46864: result <= 12'b111111001110;
   46865: result <= 12'b111111001110;
   46866: result <= 12'b111111001111;
   46867: result <= 12'b111111001111;
   46868: result <= 12'b111111001111;
   46869: result <= 12'b111111001111;
   46870: result <= 12'b111111001111;
   46871: result <= 12'b111111001111;
   46872: result <= 12'b111111001111;
   46873: result <= 12'b111111001111;
   46874: result <= 12'b111111001111;
   46875: result <= 12'b111111001111;
   46876: result <= 12'b111111001111;
   46877: result <= 12'b111111001111;
   46878: result <= 12'b111111001111;
   46879: result <= 12'b111111001111;
   46880: result <= 12'b111111001111;
   46881: result <= 12'b111111001111;
   46882: result <= 12'b111111001111;
   46883: result <= 12'b111111001111;
   46884: result <= 12'b111111001111;
   46885: result <= 12'b111111001111;
   46886: result <= 12'b111111001111;
   46887: result <= 12'b111111001111;
   46888: result <= 12'b111111001111;
   46889: result <= 12'b111111001111;
   46890: result <= 12'b111111010000;
   46891: result <= 12'b111111010000;
   46892: result <= 12'b111111010000;
   46893: result <= 12'b111111010000;
   46894: result <= 12'b111111010000;
   46895: result <= 12'b111111010000;
   46896: result <= 12'b111111010000;
   46897: result <= 12'b111111010000;
   46898: result <= 12'b111111010000;
   46899: result <= 12'b111111010000;
   46900: result <= 12'b111111010000;
   46901: result <= 12'b111111010000;
   46902: result <= 12'b111111010000;
   46903: result <= 12'b111111010000;
   46904: result <= 12'b111111010000;
   46905: result <= 12'b111111010000;
   46906: result <= 12'b111111010000;
   46907: result <= 12'b111111010000;
   46908: result <= 12'b111111010000;
   46909: result <= 12'b111111010000;
   46910: result <= 12'b111111010000;
   46911: result <= 12'b111111010000;
   46912: result <= 12'b111111010000;
   46913: result <= 12'b111111010000;
   46914: result <= 12'b111111010001;
   46915: result <= 12'b111111010001;
   46916: result <= 12'b111111010001;
   46917: result <= 12'b111111010001;
   46918: result <= 12'b111111010001;
   46919: result <= 12'b111111010001;
   46920: result <= 12'b111111010001;
   46921: result <= 12'b111111010001;
   46922: result <= 12'b111111010001;
   46923: result <= 12'b111111010001;
   46924: result <= 12'b111111010001;
   46925: result <= 12'b111111010001;
   46926: result <= 12'b111111010001;
   46927: result <= 12'b111111010001;
   46928: result <= 12'b111111010001;
   46929: result <= 12'b111111010001;
   46930: result <= 12'b111111010001;
   46931: result <= 12'b111111010001;
   46932: result <= 12'b111111010001;
   46933: result <= 12'b111111010001;
   46934: result <= 12'b111111010001;
   46935: result <= 12'b111111010001;
   46936: result <= 12'b111111010001;
   46937: result <= 12'b111111010001;
   46938: result <= 12'b111111010010;
   46939: result <= 12'b111111010010;
   46940: result <= 12'b111111010010;
   46941: result <= 12'b111111010010;
   46942: result <= 12'b111111010010;
   46943: result <= 12'b111111010010;
   46944: result <= 12'b111111010010;
   46945: result <= 12'b111111010010;
   46946: result <= 12'b111111010010;
   46947: result <= 12'b111111010010;
   46948: result <= 12'b111111010010;
   46949: result <= 12'b111111010010;
   46950: result <= 12'b111111010010;
   46951: result <= 12'b111111010010;
   46952: result <= 12'b111111010010;
   46953: result <= 12'b111111010010;
   46954: result <= 12'b111111010010;
   46955: result <= 12'b111111010010;
   46956: result <= 12'b111111010010;
   46957: result <= 12'b111111010010;
   46958: result <= 12'b111111010010;
   46959: result <= 12'b111111010010;
   46960: result <= 12'b111111010010;
   46961: result <= 12'b111111010010;
   46962: result <= 12'b111111010011;
   46963: result <= 12'b111111010011;
   46964: result <= 12'b111111010011;
   46965: result <= 12'b111111010011;
   46966: result <= 12'b111111010011;
   46967: result <= 12'b111111010011;
   46968: result <= 12'b111111010011;
   46969: result <= 12'b111111010011;
   46970: result <= 12'b111111010011;
   46971: result <= 12'b111111010011;
   46972: result <= 12'b111111010011;
   46973: result <= 12'b111111010011;
   46974: result <= 12'b111111010011;
   46975: result <= 12'b111111010011;
   46976: result <= 12'b111111010011;
   46977: result <= 12'b111111010011;
   46978: result <= 12'b111111010011;
   46979: result <= 12'b111111010011;
   46980: result <= 12'b111111010011;
   46981: result <= 12'b111111010011;
   46982: result <= 12'b111111010011;
   46983: result <= 12'b111111010011;
   46984: result <= 12'b111111010011;
   46985: result <= 12'b111111010011;
   46986: result <= 12'b111111010011;
   46987: result <= 12'b111111010100;
   46988: result <= 12'b111111010100;
   46989: result <= 12'b111111010100;
   46990: result <= 12'b111111010100;
   46991: result <= 12'b111111010100;
   46992: result <= 12'b111111010100;
   46993: result <= 12'b111111010100;
   46994: result <= 12'b111111010100;
   46995: result <= 12'b111111010100;
   46996: result <= 12'b111111010100;
   46997: result <= 12'b111111010100;
   46998: result <= 12'b111111010100;
   46999: result <= 12'b111111010100;
   47000: result <= 12'b111111010100;
   47001: result <= 12'b111111010100;
   47002: result <= 12'b111111010100;
   47003: result <= 12'b111111010100;
   47004: result <= 12'b111111010100;
   47005: result <= 12'b111111010100;
   47006: result <= 12'b111111010100;
   47007: result <= 12'b111111010100;
   47008: result <= 12'b111111010100;
   47009: result <= 12'b111111010100;
   47010: result <= 12'b111111010100;
   47011: result <= 12'b111111010101;
   47012: result <= 12'b111111010101;
   47013: result <= 12'b111111010101;
   47014: result <= 12'b111111010101;
   47015: result <= 12'b111111010101;
   47016: result <= 12'b111111010101;
   47017: result <= 12'b111111010101;
   47018: result <= 12'b111111010101;
   47019: result <= 12'b111111010101;
   47020: result <= 12'b111111010101;
   47021: result <= 12'b111111010101;
   47022: result <= 12'b111111010101;
   47023: result <= 12'b111111010101;
   47024: result <= 12'b111111010101;
   47025: result <= 12'b111111010101;
   47026: result <= 12'b111111010101;
   47027: result <= 12'b111111010101;
   47028: result <= 12'b111111010101;
   47029: result <= 12'b111111010101;
   47030: result <= 12'b111111010101;
   47031: result <= 12'b111111010101;
   47032: result <= 12'b111111010101;
   47033: result <= 12'b111111010101;
   47034: result <= 12'b111111010101;
   47035: result <= 12'b111111010101;
   47036: result <= 12'b111111010110;
   47037: result <= 12'b111111010110;
   47038: result <= 12'b111111010110;
   47039: result <= 12'b111111010110;
   47040: result <= 12'b111111010110;
   47041: result <= 12'b111111010110;
   47042: result <= 12'b111111010110;
   47043: result <= 12'b111111010110;
   47044: result <= 12'b111111010110;
   47045: result <= 12'b111111010110;
   47046: result <= 12'b111111010110;
   47047: result <= 12'b111111010110;
   47048: result <= 12'b111111010110;
   47049: result <= 12'b111111010110;
   47050: result <= 12'b111111010110;
   47051: result <= 12'b111111010110;
   47052: result <= 12'b111111010110;
   47053: result <= 12'b111111010110;
   47054: result <= 12'b111111010110;
   47055: result <= 12'b111111010110;
   47056: result <= 12'b111111010110;
   47057: result <= 12'b111111010110;
   47058: result <= 12'b111111010110;
   47059: result <= 12'b111111010110;
   47060: result <= 12'b111111010110;
   47061: result <= 12'b111111010110;
   47062: result <= 12'b111111010111;
   47063: result <= 12'b111111010111;
   47064: result <= 12'b111111010111;
   47065: result <= 12'b111111010111;
   47066: result <= 12'b111111010111;
   47067: result <= 12'b111111010111;
   47068: result <= 12'b111111010111;
   47069: result <= 12'b111111010111;
   47070: result <= 12'b111111010111;
   47071: result <= 12'b111111010111;
   47072: result <= 12'b111111010111;
   47073: result <= 12'b111111010111;
   47074: result <= 12'b111111010111;
   47075: result <= 12'b111111010111;
   47076: result <= 12'b111111010111;
   47077: result <= 12'b111111010111;
   47078: result <= 12'b111111010111;
   47079: result <= 12'b111111010111;
   47080: result <= 12'b111111010111;
   47081: result <= 12'b111111010111;
   47082: result <= 12'b111111010111;
   47083: result <= 12'b111111010111;
   47084: result <= 12'b111111010111;
   47085: result <= 12'b111111010111;
   47086: result <= 12'b111111010111;
   47087: result <= 12'b111111010111;
   47088: result <= 12'b111111011000;
   47089: result <= 12'b111111011000;
   47090: result <= 12'b111111011000;
   47091: result <= 12'b111111011000;
   47092: result <= 12'b111111011000;
   47093: result <= 12'b111111011000;
   47094: result <= 12'b111111011000;
   47095: result <= 12'b111111011000;
   47096: result <= 12'b111111011000;
   47097: result <= 12'b111111011000;
   47098: result <= 12'b111111011000;
   47099: result <= 12'b111111011000;
   47100: result <= 12'b111111011000;
   47101: result <= 12'b111111011000;
   47102: result <= 12'b111111011000;
   47103: result <= 12'b111111011000;
   47104: result <= 12'b111111011000;
   47105: result <= 12'b111111011000;
   47106: result <= 12'b111111011000;
   47107: result <= 12'b111111011000;
   47108: result <= 12'b111111011000;
   47109: result <= 12'b111111011000;
   47110: result <= 12'b111111011000;
   47111: result <= 12'b111111011000;
   47112: result <= 12'b111111011000;
   47113: result <= 12'b111111011000;
   47114: result <= 12'b111111011001;
   47115: result <= 12'b111111011001;
   47116: result <= 12'b111111011001;
   47117: result <= 12'b111111011001;
   47118: result <= 12'b111111011001;
   47119: result <= 12'b111111011001;
   47120: result <= 12'b111111011001;
   47121: result <= 12'b111111011001;
   47122: result <= 12'b111111011001;
   47123: result <= 12'b111111011001;
   47124: result <= 12'b111111011001;
   47125: result <= 12'b111111011001;
   47126: result <= 12'b111111011001;
   47127: result <= 12'b111111011001;
   47128: result <= 12'b111111011001;
   47129: result <= 12'b111111011001;
   47130: result <= 12'b111111011001;
   47131: result <= 12'b111111011001;
   47132: result <= 12'b111111011001;
   47133: result <= 12'b111111011001;
   47134: result <= 12'b111111011001;
   47135: result <= 12'b111111011001;
   47136: result <= 12'b111111011001;
   47137: result <= 12'b111111011001;
   47138: result <= 12'b111111011001;
   47139: result <= 12'b111111011001;
   47140: result <= 12'b111111011010;
   47141: result <= 12'b111111011010;
   47142: result <= 12'b111111011010;
   47143: result <= 12'b111111011010;
   47144: result <= 12'b111111011010;
   47145: result <= 12'b111111011010;
   47146: result <= 12'b111111011010;
   47147: result <= 12'b111111011010;
   47148: result <= 12'b111111011010;
   47149: result <= 12'b111111011010;
   47150: result <= 12'b111111011010;
   47151: result <= 12'b111111011010;
   47152: result <= 12'b111111011010;
   47153: result <= 12'b111111011010;
   47154: result <= 12'b111111011010;
   47155: result <= 12'b111111011010;
   47156: result <= 12'b111111011010;
   47157: result <= 12'b111111011010;
   47158: result <= 12'b111111011010;
   47159: result <= 12'b111111011010;
   47160: result <= 12'b111111011010;
   47161: result <= 12'b111111011010;
   47162: result <= 12'b111111011010;
   47163: result <= 12'b111111011010;
   47164: result <= 12'b111111011010;
   47165: result <= 12'b111111011010;
   47166: result <= 12'b111111011010;
   47167: result <= 12'b111111011011;
   47168: result <= 12'b111111011011;
   47169: result <= 12'b111111011011;
   47170: result <= 12'b111111011011;
   47171: result <= 12'b111111011011;
   47172: result <= 12'b111111011011;
   47173: result <= 12'b111111011011;
   47174: result <= 12'b111111011011;
   47175: result <= 12'b111111011011;
   47176: result <= 12'b111111011011;
   47177: result <= 12'b111111011011;
   47178: result <= 12'b111111011011;
   47179: result <= 12'b111111011011;
   47180: result <= 12'b111111011011;
   47181: result <= 12'b111111011011;
   47182: result <= 12'b111111011011;
   47183: result <= 12'b111111011011;
   47184: result <= 12'b111111011011;
   47185: result <= 12'b111111011011;
   47186: result <= 12'b111111011011;
   47187: result <= 12'b111111011011;
   47188: result <= 12'b111111011011;
   47189: result <= 12'b111111011011;
   47190: result <= 12'b111111011011;
   47191: result <= 12'b111111011011;
   47192: result <= 12'b111111011011;
   47193: result <= 12'b111111011011;
   47194: result <= 12'b111111011100;
   47195: result <= 12'b111111011100;
   47196: result <= 12'b111111011100;
   47197: result <= 12'b111111011100;
   47198: result <= 12'b111111011100;
   47199: result <= 12'b111111011100;
   47200: result <= 12'b111111011100;
   47201: result <= 12'b111111011100;
   47202: result <= 12'b111111011100;
   47203: result <= 12'b111111011100;
   47204: result <= 12'b111111011100;
   47205: result <= 12'b111111011100;
   47206: result <= 12'b111111011100;
   47207: result <= 12'b111111011100;
   47208: result <= 12'b111111011100;
   47209: result <= 12'b111111011100;
   47210: result <= 12'b111111011100;
   47211: result <= 12'b111111011100;
   47212: result <= 12'b111111011100;
   47213: result <= 12'b111111011100;
   47214: result <= 12'b111111011100;
   47215: result <= 12'b111111011100;
   47216: result <= 12'b111111011100;
   47217: result <= 12'b111111011100;
   47218: result <= 12'b111111011100;
   47219: result <= 12'b111111011100;
   47220: result <= 12'b111111011100;
   47221: result <= 12'b111111011101;
   47222: result <= 12'b111111011101;
   47223: result <= 12'b111111011101;
   47224: result <= 12'b111111011101;
   47225: result <= 12'b111111011101;
   47226: result <= 12'b111111011101;
   47227: result <= 12'b111111011101;
   47228: result <= 12'b111111011101;
   47229: result <= 12'b111111011101;
   47230: result <= 12'b111111011101;
   47231: result <= 12'b111111011101;
   47232: result <= 12'b111111011101;
   47233: result <= 12'b111111011101;
   47234: result <= 12'b111111011101;
   47235: result <= 12'b111111011101;
   47236: result <= 12'b111111011101;
   47237: result <= 12'b111111011101;
   47238: result <= 12'b111111011101;
   47239: result <= 12'b111111011101;
   47240: result <= 12'b111111011101;
   47241: result <= 12'b111111011101;
   47242: result <= 12'b111111011101;
   47243: result <= 12'b111111011101;
   47244: result <= 12'b111111011101;
   47245: result <= 12'b111111011101;
   47246: result <= 12'b111111011101;
   47247: result <= 12'b111111011101;
   47248: result <= 12'b111111011101;
   47249: result <= 12'b111111011110;
   47250: result <= 12'b111111011110;
   47251: result <= 12'b111111011110;
   47252: result <= 12'b111111011110;
   47253: result <= 12'b111111011110;
   47254: result <= 12'b111111011110;
   47255: result <= 12'b111111011110;
   47256: result <= 12'b111111011110;
   47257: result <= 12'b111111011110;
   47258: result <= 12'b111111011110;
   47259: result <= 12'b111111011110;
   47260: result <= 12'b111111011110;
   47261: result <= 12'b111111011110;
   47262: result <= 12'b111111011110;
   47263: result <= 12'b111111011110;
   47264: result <= 12'b111111011110;
   47265: result <= 12'b111111011110;
   47266: result <= 12'b111111011110;
   47267: result <= 12'b111111011110;
   47268: result <= 12'b111111011110;
   47269: result <= 12'b111111011110;
   47270: result <= 12'b111111011110;
   47271: result <= 12'b111111011110;
   47272: result <= 12'b111111011110;
   47273: result <= 12'b111111011110;
   47274: result <= 12'b111111011110;
   47275: result <= 12'b111111011110;
   47276: result <= 12'b111111011110;
   47277: result <= 12'b111111011110;
   47278: result <= 12'b111111011111;
   47279: result <= 12'b111111011111;
   47280: result <= 12'b111111011111;
   47281: result <= 12'b111111011111;
   47282: result <= 12'b111111011111;
   47283: result <= 12'b111111011111;
   47284: result <= 12'b111111011111;
   47285: result <= 12'b111111011111;
   47286: result <= 12'b111111011111;
   47287: result <= 12'b111111011111;
   47288: result <= 12'b111111011111;
   47289: result <= 12'b111111011111;
   47290: result <= 12'b111111011111;
   47291: result <= 12'b111111011111;
   47292: result <= 12'b111111011111;
   47293: result <= 12'b111111011111;
   47294: result <= 12'b111111011111;
   47295: result <= 12'b111111011111;
   47296: result <= 12'b111111011111;
   47297: result <= 12'b111111011111;
   47298: result <= 12'b111111011111;
   47299: result <= 12'b111111011111;
   47300: result <= 12'b111111011111;
   47301: result <= 12'b111111011111;
   47302: result <= 12'b111111011111;
   47303: result <= 12'b111111011111;
   47304: result <= 12'b111111011111;
   47305: result <= 12'b111111011111;
   47306: result <= 12'b111111100000;
   47307: result <= 12'b111111100000;
   47308: result <= 12'b111111100000;
   47309: result <= 12'b111111100000;
   47310: result <= 12'b111111100000;
   47311: result <= 12'b111111100000;
   47312: result <= 12'b111111100000;
   47313: result <= 12'b111111100000;
   47314: result <= 12'b111111100000;
   47315: result <= 12'b111111100000;
   47316: result <= 12'b111111100000;
   47317: result <= 12'b111111100000;
   47318: result <= 12'b111111100000;
   47319: result <= 12'b111111100000;
   47320: result <= 12'b111111100000;
   47321: result <= 12'b111111100000;
   47322: result <= 12'b111111100000;
   47323: result <= 12'b111111100000;
   47324: result <= 12'b111111100000;
   47325: result <= 12'b111111100000;
   47326: result <= 12'b111111100000;
   47327: result <= 12'b111111100000;
   47328: result <= 12'b111111100000;
   47329: result <= 12'b111111100000;
   47330: result <= 12'b111111100000;
   47331: result <= 12'b111111100000;
   47332: result <= 12'b111111100000;
   47333: result <= 12'b111111100000;
   47334: result <= 12'b111111100000;
   47335: result <= 12'b111111100001;
   47336: result <= 12'b111111100001;
   47337: result <= 12'b111111100001;
   47338: result <= 12'b111111100001;
   47339: result <= 12'b111111100001;
   47340: result <= 12'b111111100001;
   47341: result <= 12'b111111100001;
   47342: result <= 12'b111111100001;
   47343: result <= 12'b111111100001;
   47344: result <= 12'b111111100001;
   47345: result <= 12'b111111100001;
   47346: result <= 12'b111111100001;
   47347: result <= 12'b111111100001;
   47348: result <= 12'b111111100001;
   47349: result <= 12'b111111100001;
   47350: result <= 12'b111111100001;
   47351: result <= 12'b111111100001;
   47352: result <= 12'b111111100001;
   47353: result <= 12'b111111100001;
   47354: result <= 12'b111111100001;
   47355: result <= 12'b111111100001;
   47356: result <= 12'b111111100001;
   47357: result <= 12'b111111100001;
   47358: result <= 12'b111111100001;
   47359: result <= 12'b111111100001;
   47360: result <= 12'b111111100001;
   47361: result <= 12'b111111100001;
   47362: result <= 12'b111111100001;
   47363: result <= 12'b111111100001;
   47364: result <= 12'b111111100001;
   47365: result <= 12'b111111100010;
   47366: result <= 12'b111111100010;
   47367: result <= 12'b111111100010;
   47368: result <= 12'b111111100010;
   47369: result <= 12'b111111100010;
   47370: result <= 12'b111111100010;
   47371: result <= 12'b111111100010;
   47372: result <= 12'b111111100010;
   47373: result <= 12'b111111100010;
   47374: result <= 12'b111111100010;
   47375: result <= 12'b111111100010;
   47376: result <= 12'b111111100010;
   47377: result <= 12'b111111100010;
   47378: result <= 12'b111111100010;
   47379: result <= 12'b111111100010;
   47380: result <= 12'b111111100010;
   47381: result <= 12'b111111100010;
   47382: result <= 12'b111111100010;
   47383: result <= 12'b111111100010;
   47384: result <= 12'b111111100010;
   47385: result <= 12'b111111100010;
   47386: result <= 12'b111111100010;
   47387: result <= 12'b111111100010;
   47388: result <= 12'b111111100010;
   47389: result <= 12'b111111100010;
   47390: result <= 12'b111111100010;
   47391: result <= 12'b111111100010;
   47392: result <= 12'b111111100010;
   47393: result <= 12'b111111100010;
   47394: result <= 12'b111111100010;
   47395: result <= 12'b111111100011;
   47396: result <= 12'b111111100011;
   47397: result <= 12'b111111100011;
   47398: result <= 12'b111111100011;
   47399: result <= 12'b111111100011;
   47400: result <= 12'b111111100011;
   47401: result <= 12'b111111100011;
   47402: result <= 12'b111111100011;
   47403: result <= 12'b111111100011;
   47404: result <= 12'b111111100011;
   47405: result <= 12'b111111100011;
   47406: result <= 12'b111111100011;
   47407: result <= 12'b111111100011;
   47408: result <= 12'b111111100011;
   47409: result <= 12'b111111100011;
   47410: result <= 12'b111111100011;
   47411: result <= 12'b111111100011;
   47412: result <= 12'b111111100011;
   47413: result <= 12'b111111100011;
   47414: result <= 12'b111111100011;
   47415: result <= 12'b111111100011;
   47416: result <= 12'b111111100011;
   47417: result <= 12'b111111100011;
   47418: result <= 12'b111111100011;
   47419: result <= 12'b111111100011;
   47420: result <= 12'b111111100011;
   47421: result <= 12'b111111100011;
   47422: result <= 12'b111111100011;
   47423: result <= 12'b111111100011;
   47424: result <= 12'b111111100011;
   47425: result <= 12'b111111100011;
   47426: result <= 12'b111111100100;
   47427: result <= 12'b111111100100;
   47428: result <= 12'b111111100100;
   47429: result <= 12'b111111100100;
   47430: result <= 12'b111111100100;
   47431: result <= 12'b111111100100;
   47432: result <= 12'b111111100100;
   47433: result <= 12'b111111100100;
   47434: result <= 12'b111111100100;
   47435: result <= 12'b111111100100;
   47436: result <= 12'b111111100100;
   47437: result <= 12'b111111100100;
   47438: result <= 12'b111111100100;
   47439: result <= 12'b111111100100;
   47440: result <= 12'b111111100100;
   47441: result <= 12'b111111100100;
   47442: result <= 12'b111111100100;
   47443: result <= 12'b111111100100;
   47444: result <= 12'b111111100100;
   47445: result <= 12'b111111100100;
   47446: result <= 12'b111111100100;
   47447: result <= 12'b111111100100;
   47448: result <= 12'b111111100100;
   47449: result <= 12'b111111100100;
   47450: result <= 12'b111111100100;
   47451: result <= 12'b111111100100;
   47452: result <= 12'b111111100100;
   47453: result <= 12'b111111100100;
   47454: result <= 12'b111111100100;
   47455: result <= 12'b111111100100;
   47456: result <= 12'b111111100100;
   47457: result <= 12'b111111100101;
   47458: result <= 12'b111111100101;
   47459: result <= 12'b111111100101;
   47460: result <= 12'b111111100101;
   47461: result <= 12'b111111100101;
   47462: result <= 12'b111111100101;
   47463: result <= 12'b111111100101;
   47464: result <= 12'b111111100101;
   47465: result <= 12'b111111100101;
   47466: result <= 12'b111111100101;
   47467: result <= 12'b111111100101;
   47468: result <= 12'b111111100101;
   47469: result <= 12'b111111100101;
   47470: result <= 12'b111111100101;
   47471: result <= 12'b111111100101;
   47472: result <= 12'b111111100101;
   47473: result <= 12'b111111100101;
   47474: result <= 12'b111111100101;
   47475: result <= 12'b111111100101;
   47476: result <= 12'b111111100101;
   47477: result <= 12'b111111100101;
   47478: result <= 12'b111111100101;
   47479: result <= 12'b111111100101;
   47480: result <= 12'b111111100101;
   47481: result <= 12'b111111100101;
   47482: result <= 12'b111111100101;
   47483: result <= 12'b111111100101;
   47484: result <= 12'b111111100101;
   47485: result <= 12'b111111100101;
   47486: result <= 12'b111111100101;
   47487: result <= 12'b111111100101;
   47488: result <= 12'b111111100101;
   47489: result <= 12'b111111100110;
   47490: result <= 12'b111111100110;
   47491: result <= 12'b111111100110;
   47492: result <= 12'b111111100110;
   47493: result <= 12'b111111100110;
   47494: result <= 12'b111111100110;
   47495: result <= 12'b111111100110;
   47496: result <= 12'b111111100110;
   47497: result <= 12'b111111100110;
   47498: result <= 12'b111111100110;
   47499: result <= 12'b111111100110;
   47500: result <= 12'b111111100110;
   47501: result <= 12'b111111100110;
   47502: result <= 12'b111111100110;
   47503: result <= 12'b111111100110;
   47504: result <= 12'b111111100110;
   47505: result <= 12'b111111100110;
   47506: result <= 12'b111111100110;
   47507: result <= 12'b111111100110;
   47508: result <= 12'b111111100110;
   47509: result <= 12'b111111100110;
   47510: result <= 12'b111111100110;
   47511: result <= 12'b111111100110;
   47512: result <= 12'b111111100110;
   47513: result <= 12'b111111100110;
   47514: result <= 12'b111111100110;
   47515: result <= 12'b111111100110;
   47516: result <= 12'b111111100110;
   47517: result <= 12'b111111100110;
   47518: result <= 12'b111111100110;
   47519: result <= 12'b111111100110;
   47520: result <= 12'b111111100110;
   47521: result <= 12'b111111100111;
   47522: result <= 12'b111111100111;
   47523: result <= 12'b111111100111;
   47524: result <= 12'b111111100111;
   47525: result <= 12'b111111100111;
   47526: result <= 12'b111111100111;
   47527: result <= 12'b111111100111;
   47528: result <= 12'b111111100111;
   47529: result <= 12'b111111100111;
   47530: result <= 12'b111111100111;
   47531: result <= 12'b111111100111;
   47532: result <= 12'b111111100111;
   47533: result <= 12'b111111100111;
   47534: result <= 12'b111111100111;
   47535: result <= 12'b111111100111;
   47536: result <= 12'b111111100111;
   47537: result <= 12'b111111100111;
   47538: result <= 12'b111111100111;
   47539: result <= 12'b111111100111;
   47540: result <= 12'b111111100111;
   47541: result <= 12'b111111100111;
   47542: result <= 12'b111111100111;
   47543: result <= 12'b111111100111;
   47544: result <= 12'b111111100111;
   47545: result <= 12'b111111100111;
   47546: result <= 12'b111111100111;
   47547: result <= 12'b111111100111;
   47548: result <= 12'b111111100111;
   47549: result <= 12'b111111100111;
   47550: result <= 12'b111111100111;
   47551: result <= 12'b111111100111;
   47552: result <= 12'b111111100111;
   47553: result <= 12'b111111100111;
   47554: result <= 12'b111111101000;
   47555: result <= 12'b111111101000;
   47556: result <= 12'b111111101000;
   47557: result <= 12'b111111101000;
   47558: result <= 12'b111111101000;
   47559: result <= 12'b111111101000;
   47560: result <= 12'b111111101000;
   47561: result <= 12'b111111101000;
   47562: result <= 12'b111111101000;
   47563: result <= 12'b111111101000;
   47564: result <= 12'b111111101000;
   47565: result <= 12'b111111101000;
   47566: result <= 12'b111111101000;
   47567: result <= 12'b111111101000;
   47568: result <= 12'b111111101000;
   47569: result <= 12'b111111101000;
   47570: result <= 12'b111111101000;
   47571: result <= 12'b111111101000;
   47572: result <= 12'b111111101000;
   47573: result <= 12'b111111101000;
   47574: result <= 12'b111111101000;
   47575: result <= 12'b111111101000;
   47576: result <= 12'b111111101000;
   47577: result <= 12'b111111101000;
   47578: result <= 12'b111111101000;
   47579: result <= 12'b111111101000;
   47580: result <= 12'b111111101000;
   47581: result <= 12'b111111101000;
   47582: result <= 12'b111111101000;
   47583: result <= 12'b111111101000;
   47584: result <= 12'b111111101000;
   47585: result <= 12'b111111101000;
   47586: result <= 12'b111111101000;
   47587: result <= 12'b111111101000;
   47588: result <= 12'b111111101001;
   47589: result <= 12'b111111101001;
   47590: result <= 12'b111111101001;
   47591: result <= 12'b111111101001;
   47592: result <= 12'b111111101001;
   47593: result <= 12'b111111101001;
   47594: result <= 12'b111111101001;
   47595: result <= 12'b111111101001;
   47596: result <= 12'b111111101001;
   47597: result <= 12'b111111101001;
   47598: result <= 12'b111111101001;
   47599: result <= 12'b111111101001;
   47600: result <= 12'b111111101001;
   47601: result <= 12'b111111101001;
   47602: result <= 12'b111111101001;
   47603: result <= 12'b111111101001;
   47604: result <= 12'b111111101001;
   47605: result <= 12'b111111101001;
   47606: result <= 12'b111111101001;
   47607: result <= 12'b111111101001;
   47608: result <= 12'b111111101001;
   47609: result <= 12'b111111101001;
   47610: result <= 12'b111111101001;
   47611: result <= 12'b111111101001;
   47612: result <= 12'b111111101001;
   47613: result <= 12'b111111101001;
   47614: result <= 12'b111111101001;
   47615: result <= 12'b111111101001;
   47616: result <= 12'b111111101001;
   47617: result <= 12'b111111101001;
   47618: result <= 12'b111111101001;
   47619: result <= 12'b111111101001;
   47620: result <= 12'b111111101001;
   47621: result <= 12'b111111101001;
   47622: result <= 12'b111111101010;
   47623: result <= 12'b111111101010;
   47624: result <= 12'b111111101010;
   47625: result <= 12'b111111101010;
   47626: result <= 12'b111111101010;
   47627: result <= 12'b111111101010;
   47628: result <= 12'b111111101010;
   47629: result <= 12'b111111101010;
   47630: result <= 12'b111111101010;
   47631: result <= 12'b111111101010;
   47632: result <= 12'b111111101010;
   47633: result <= 12'b111111101010;
   47634: result <= 12'b111111101010;
   47635: result <= 12'b111111101010;
   47636: result <= 12'b111111101010;
   47637: result <= 12'b111111101010;
   47638: result <= 12'b111111101010;
   47639: result <= 12'b111111101010;
   47640: result <= 12'b111111101010;
   47641: result <= 12'b111111101010;
   47642: result <= 12'b111111101010;
   47643: result <= 12'b111111101010;
   47644: result <= 12'b111111101010;
   47645: result <= 12'b111111101010;
   47646: result <= 12'b111111101010;
   47647: result <= 12'b111111101010;
   47648: result <= 12'b111111101010;
   47649: result <= 12'b111111101010;
   47650: result <= 12'b111111101010;
   47651: result <= 12'b111111101010;
   47652: result <= 12'b111111101010;
   47653: result <= 12'b111111101010;
   47654: result <= 12'b111111101010;
   47655: result <= 12'b111111101010;
   47656: result <= 12'b111111101010;
   47657: result <= 12'b111111101010;
   47658: result <= 12'b111111101011;
   47659: result <= 12'b111111101011;
   47660: result <= 12'b111111101011;
   47661: result <= 12'b111111101011;
   47662: result <= 12'b111111101011;
   47663: result <= 12'b111111101011;
   47664: result <= 12'b111111101011;
   47665: result <= 12'b111111101011;
   47666: result <= 12'b111111101011;
   47667: result <= 12'b111111101011;
   47668: result <= 12'b111111101011;
   47669: result <= 12'b111111101011;
   47670: result <= 12'b111111101011;
   47671: result <= 12'b111111101011;
   47672: result <= 12'b111111101011;
   47673: result <= 12'b111111101011;
   47674: result <= 12'b111111101011;
   47675: result <= 12'b111111101011;
   47676: result <= 12'b111111101011;
   47677: result <= 12'b111111101011;
   47678: result <= 12'b111111101011;
   47679: result <= 12'b111111101011;
   47680: result <= 12'b111111101011;
   47681: result <= 12'b111111101011;
   47682: result <= 12'b111111101011;
   47683: result <= 12'b111111101011;
   47684: result <= 12'b111111101011;
   47685: result <= 12'b111111101011;
   47686: result <= 12'b111111101011;
   47687: result <= 12'b111111101011;
   47688: result <= 12'b111111101011;
   47689: result <= 12'b111111101011;
   47690: result <= 12'b111111101011;
   47691: result <= 12'b111111101011;
   47692: result <= 12'b111111101011;
   47693: result <= 12'b111111101011;
   47694: result <= 12'b111111101100;
   47695: result <= 12'b111111101100;
   47696: result <= 12'b111111101100;
   47697: result <= 12'b111111101100;
   47698: result <= 12'b111111101100;
   47699: result <= 12'b111111101100;
   47700: result <= 12'b111111101100;
   47701: result <= 12'b111111101100;
   47702: result <= 12'b111111101100;
   47703: result <= 12'b111111101100;
   47704: result <= 12'b111111101100;
   47705: result <= 12'b111111101100;
   47706: result <= 12'b111111101100;
   47707: result <= 12'b111111101100;
   47708: result <= 12'b111111101100;
   47709: result <= 12'b111111101100;
   47710: result <= 12'b111111101100;
   47711: result <= 12'b111111101100;
   47712: result <= 12'b111111101100;
   47713: result <= 12'b111111101100;
   47714: result <= 12'b111111101100;
   47715: result <= 12'b111111101100;
   47716: result <= 12'b111111101100;
   47717: result <= 12'b111111101100;
   47718: result <= 12'b111111101100;
   47719: result <= 12'b111111101100;
   47720: result <= 12'b111111101100;
   47721: result <= 12'b111111101100;
   47722: result <= 12'b111111101100;
   47723: result <= 12'b111111101100;
   47724: result <= 12'b111111101100;
   47725: result <= 12'b111111101100;
   47726: result <= 12'b111111101100;
   47727: result <= 12'b111111101100;
   47728: result <= 12'b111111101100;
   47729: result <= 12'b111111101100;
   47730: result <= 12'b111111101100;
   47731: result <= 12'b111111101101;
   47732: result <= 12'b111111101101;
   47733: result <= 12'b111111101101;
   47734: result <= 12'b111111101101;
   47735: result <= 12'b111111101101;
   47736: result <= 12'b111111101101;
   47737: result <= 12'b111111101101;
   47738: result <= 12'b111111101101;
   47739: result <= 12'b111111101101;
   47740: result <= 12'b111111101101;
   47741: result <= 12'b111111101101;
   47742: result <= 12'b111111101101;
   47743: result <= 12'b111111101101;
   47744: result <= 12'b111111101101;
   47745: result <= 12'b111111101101;
   47746: result <= 12'b111111101101;
   47747: result <= 12'b111111101101;
   47748: result <= 12'b111111101101;
   47749: result <= 12'b111111101101;
   47750: result <= 12'b111111101101;
   47751: result <= 12'b111111101101;
   47752: result <= 12'b111111101101;
   47753: result <= 12'b111111101101;
   47754: result <= 12'b111111101101;
   47755: result <= 12'b111111101101;
   47756: result <= 12'b111111101101;
   47757: result <= 12'b111111101101;
   47758: result <= 12'b111111101101;
   47759: result <= 12'b111111101101;
   47760: result <= 12'b111111101101;
   47761: result <= 12'b111111101101;
   47762: result <= 12'b111111101101;
   47763: result <= 12'b111111101101;
   47764: result <= 12'b111111101101;
   47765: result <= 12'b111111101101;
   47766: result <= 12'b111111101101;
   47767: result <= 12'b111111101101;
   47768: result <= 12'b111111101101;
   47769: result <= 12'b111111101110;
   47770: result <= 12'b111111101110;
   47771: result <= 12'b111111101110;
   47772: result <= 12'b111111101110;
   47773: result <= 12'b111111101110;
   47774: result <= 12'b111111101110;
   47775: result <= 12'b111111101110;
   47776: result <= 12'b111111101110;
   47777: result <= 12'b111111101110;
   47778: result <= 12'b111111101110;
   47779: result <= 12'b111111101110;
   47780: result <= 12'b111111101110;
   47781: result <= 12'b111111101110;
   47782: result <= 12'b111111101110;
   47783: result <= 12'b111111101110;
   47784: result <= 12'b111111101110;
   47785: result <= 12'b111111101110;
   47786: result <= 12'b111111101110;
   47787: result <= 12'b111111101110;
   47788: result <= 12'b111111101110;
   47789: result <= 12'b111111101110;
   47790: result <= 12'b111111101110;
   47791: result <= 12'b111111101110;
   47792: result <= 12'b111111101110;
   47793: result <= 12'b111111101110;
   47794: result <= 12'b111111101110;
   47795: result <= 12'b111111101110;
   47796: result <= 12'b111111101110;
   47797: result <= 12'b111111101110;
   47798: result <= 12'b111111101110;
   47799: result <= 12'b111111101110;
   47800: result <= 12'b111111101110;
   47801: result <= 12'b111111101110;
   47802: result <= 12'b111111101110;
   47803: result <= 12'b111111101110;
   47804: result <= 12'b111111101110;
   47805: result <= 12'b111111101110;
   47806: result <= 12'b111111101110;
   47807: result <= 12'b111111101110;
   47808: result <= 12'b111111101111;
   47809: result <= 12'b111111101111;
   47810: result <= 12'b111111101111;
   47811: result <= 12'b111111101111;
   47812: result <= 12'b111111101111;
   47813: result <= 12'b111111101111;
   47814: result <= 12'b111111101111;
   47815: result <= 12'b111111101111;
   47816: result <= 12'b111111101111;
   47817: result <= 12'b111111101111;
   47818: result <= 12'b111111101111;
   47819: result <= 12'b111111101111;
   47820: result <= 12'b111111101111;
   47821: result <= 12'b111111101111;
   47822: result <= 12'b111111101111;
   47823: result <= 12'b111111101111;
   47824: result <= 12'b111111101111;
   47825: result <= 12'b111111101111;
   47826: result <= 12'b111111101111;
   47827: result <= 12'b111111101111;
   47828: result <= 12'b111111101111;
   47829: result <= 12'b111111101111;
   47830: result <= 12'b111111101111;
   47831: result <= 12'b111111101111;
   47832: result <= 12'b111111101111;
   47833: result <= 12'b111111101111;
   47834: result <= 12'b111111101111;
   47835: result <= 12'b111111101111;
   47836: result <= 12'b111111101111;
   47837: result <= 12'b111111101111;
   47838: result <= 12'b111111101111;
   47839: result <= 12'b111111101111;
   47840: result <= 12'b111111101111;
   47841: result <= 12'b111111101111;
   47842: result <= 12'b111111101111;
   47843: result <= 12'b111111101111;
   47844: result <= 12'b111111101111;
   47845: result <= 12'b111111101111;
   47846: result <= 12'b111111101111;
   47847: result <= 12'b111111101111;
   47848: result <= 12'b111111110000;
   47849: result <= 12'b111111110000;
   47850: result <= 12'b111111110000;
   47851: result <= 12'b111111110000;
   47852: result <= 12'b111111110000;
   47853: result <= 12'b111111110000;
   47854: result <= 12'b111111110000;
   47855: result <= 12'b111111110000;
   47856: result <= 12'b111111110000;
   47857: result <= 12'b111111110000;
   47858: result <= 12'b111111110000;
   47859: result <= 12'b111111110000;
   47860: result <= 12'b111111110000;
   47861: result <= 12'b111111110000;
   47862: result <= 12'b111111110000;
   47863: result <= 12'b111111110000;
   47864: result <= 12'b111111110000;
   47865: result <= 12'b111111110000;
   47866: result <= 12'b111111110000;
   47867: result <= 12'b111111110000;
   47868: result <= 12'b111111110000;
   47869: result <= 12'b111111110000;
   47870: result <= 12'b111111110000;
   47871: result <= 12'b111111110000;
   47872: result <= 12'b111111110000;
   47873: result <= 12'b111111110000;
   47874: result <= 12'b111111110000;
   47875: result <= 12'b111111110000;
   47876: result <= 12'b111111110000;
   47877: result <= 12'b111111110000;
   47878: result <= 12'b111111110000;
   47879: result <= 12'b111111110000;
   47880: result <= 12'b111111110000;
   47881: result <= 12'b111111110000;
   47882: result <= 12'b111111110000;
   47883: result <= 12'b111111110000;
   47884: result <= 12'b111111110000;
   47885: result <= 12'b111111110000;
   47886: result <= 12'b111111110000;
   47887: result <= 12'b111111110000;
   47888: result <= 12'b111111110000;
   47889: result <= 12'b111111110001;
   47890: result <= 12'b111111110001;
   47891: result <= 12'b111111110001;
   47892: result <= 12'b111111110001;
   47893: result <= 12'b111111110001;
   47894: result <= 12'b111111110001;
   47895: result <= 12'b111111110001;
   47896: result <= 12'b111111110001;
   47897: result <= 12'b111111110001;
   47898: result <= 12'b111111110001;
   47899: result <= 12'b111111110001;
   47900: result <= 12'b111111110001;
   47901: result <= 12'b111111110001;
   47902: result <= 12'b111111110001;
   47903: result <= 12'b111111110001;
   47904: result <= 12'b111111110001;
   47905: result <= 12'b111111110001;
   47906: result <= 12'b111111110001;
   47907: result <= 12'b111111110001;
   47908: result <= 12'b111111110001;
   47909: result <= 12'b111111110001;
   47910: result <= 12'b111111110001;
   47911: result <= 12'b111111110001;
   47912: result <= 12'b111111110001;
   47913: result <= 12'b111111110001;
   47914: result <= 12'b111111110001;
   47915: result <= 12'b111111110001;
   47916: result <= 12'b111111110001;
   47917: result <= 12'b111111110001;
   47918: result <= 12'b111111110001;
   47919: result <= 12'b111111110001;
   47920: result <= 12'b111111110001;
   47921: result <= 12'b111111110001;
   47922: result <= 12'b111111110001;
   47923: result <= 12'b111111110001;
   47924: result <= 12'b111111110001;
   47925: result <= 12'b111111110001;
   47926: result <= 12'b111111110001;
   47927: result <= 12'b111111110001;
   47928: result <= 12'b111111110001;
   47929: result <= 12'b111111110001;
   47930: result <= 12'b111111110001;
   47931: result <= 12'b111111110001;
   47932: result <= 12'b111111110010;
   47933: result <= 12'b111111110010;
   47934: result <= 12'b111111110010;
   47935: result <= 12'b111111110010;
   47936: result <= 12'b111111110010;
   47937: result <= 12'b111111110010;
   47938: result <= 12'b111111110010;
   47939: result <= 12'b111111110010;
   47940: result <= 12'b111111110010;
   47941: result <= 12'b111111110010;
   47942: result <= 12'b111111110010;
   47943: result <= 12'b111111110010;
   47944: result <= 12'b111111110010;
   47945: result <= 12'b111111110010;
   47946: result <= 12'b111111110010;
   47947: result <= 12'b111111110010;
   47948: result <= 12'b111111110010;
   47949: result <= 12'b111111110010;
   47950: result <= 12'b111111110010;
   47951: result <= 12'b111111110010;
   47952: result <= 12'b111111110010;
   47953: result <= 12'b111111110010;
   47954: result <= 12'b111111110010;
   47955: result <= 12'b111111110010;
   47956: result <= 12'b111111110010;
   47957: result <= 12'b111111110010;
   47958: result <= 12'b111111110010;
   47959: result <= 12'b111111110010;
   47960: result <= 12'b111111110010;
   47961: result <= 12'b111111110010;
   47962: result <= 12'b111111110010;
   47963: result <= 12'b111111110010;
   47964: result <= 12'b111111110010;
   47965: result <= 12'b111111110010;
   47966: result <= 12'b111111110010;
   47967: result <= 12'b111111110010;
   47968: result <= 12'b111111110010;
   47969: result <= 12'b111111110010;
   47970: result <= 12'b111111110010;
   47971: result <= 12'b111111110010;
   47972: result <= 12'b111111110010;
   47973: result <= 12'b111111110010;
   47974: result <= 12'b111111110010;
   47975: result <= 12'b111111110010;
   47976: result <= 12'b111111110010;
   47977: result <= 12'b111111110011;
   47978: result <= 12'b111111110011;
   47979: result <= 12'b111111110011;
   47980: result <= 12'b111111110011;
   47981: result <= 12'b111111110011;
   47982: result <= 12'b111111110011;
   47983: result <= 12'b111111110011;
   47984: result <= 12'b111111110011;
   47985: result <= 12'b111111110011;
   47986: result <= 12'b111111110011;
   47987: result <= 12'b111111110011;
   47988: result <= 12'b111111110011;
   47989: result <= 12'b111111110011;
   47990: result <= 12'b111111110011;
   47991: result <= 12'b111111110011;
   47992: result <= 12'b111111110011;
   47993: result <= 12'b111111110011;
   47994: result <= 12'b111111110011;
   47995: result <= 12'b111111110011;
   47996: result <= 12'b111111110011;
   47997: result <= 12'b111111110011;
   47998: result <= 12'b111111110011;
   47999: result <= 12'b111111110011;
   48000: result <= 12'b111111110011;
   48001: result <= 12'b111111110011;
   48002: result <= 12'b111111110011;
   48003: result <= 12'b111111110011;
   48004: result <= 12'b111111110011;
   48005: result <= 12'b111111110011;
   48006: result <= 12'b111111110011;
   48007: result <= 12'b111111110011;
   48008: result <= 12'b111111110011;
   48009: result <= 12'b111111110011;
   48010: result <= 12'b111111110011;
   48011: result <= 12'b111111110011;
   48012: result <= 12'b111111110011;
   48013: result <= 12'b111111110011;
   48014: result <= 12'b111111110011;
   48015: result <= 12'b111111110011;
   48016: result <= 12'b111111110011;
   48017: result <= 12'b111111110011;
   48018: result <= 12'b111111110011;
   48019: result <= 12'b111111110011;
   48020: result <= 12'b111111110011;
   48021: result <= 12'b111111110011;
   48022: result <= 12'b111111110011;
   48023: result <= 12'b111111110100;
   48024: result <= 12'b111111110100;
   48025: result <= 12'b111111110100;
   48026: result <= 12'b111111110100;
   48027: result <= 12'b111111110100;
   48028: result <= 12'b111111110100;
   48029: result <= 12'b111111110100;
   48030: result <= 12'b111111110100;
   48031: result <= 12'b111111110100;
   48032: result <= 12'b111111110100;
   48033: result <= 12'b111111110100;
   48034: result <= 12'b111111110100;
   48035: result <= 12'b111111110100;
   48036: result <= 12'b111111110100;
   48037: result <= 12'b111111110100;
   48038: result <= 12'b111111110100;
   48039: result <= 12'b111111110100;
   48040: result <= 12'b111111110100;
   48041: result <= 12'b111111110100;
   48042: result <= 12'b111111110100;
   48043: result <= 12'b111111110100;
   48044: result <= 12'b111111110100;
   48045: result <= 12'b111111110100;
   48046: result <= 12'b111111110100;
   48047: result <= 12'b111111110100;
   48048: result <= 12'b111111110100;
   48049: result <= 12'b111111110100;
   48050: result <= 12'b111111110100;
   48051: result <= 12'b111111110100;
   48052: result <= 12'b111111110100;
   48053: result <= 12'b111111110100;
   48054: result <= 12'b111111110100;
   48055: result <= 12'b111111110100;
   48056: result <= 12'b111111110100;
   48057: result <= 12'b111111110100;
   48058: result <= 12'b111111110100;
   48059: result <= 12'b111111110100;
   48060: result <= 12'b111111110100;
   48061: result <= 12'b111111110100;
   48062: result <= 12'b111111110100;
   48063: result <= 12'b111111110100;
   48064: result <= 12'b111111110100;
   48065: result <= 12'b111111110100;
   48066: result <= 12'b111111110100;
   48067: result <= 12'b111111110100;
   48068: result <= 12'b111111110100;
   48069: result <= 12'b111111110100;
   48070: result <= 12'b111111110100;
   48071: result <= 12'b111111110101;
   48072: result <= 12'b111111110101;
   48073: result <= 12'b111111110101;
   48074: result <= 12'b111111110101;
   48075: result <= 12'b111111110101;
   48076: result <= 12'b111111110101;
   48077: result <= 12'b111111110101;
   48078: result <= 12'b111111110101;
   48079: result <= 12'b111111110101;
   48080: result <= 12'b111111110101;
   48081: result <= 12'b111111110101;
   48082: result <= 12'b111111110101;
   48083: result <= 12'b111111110101;
   48084: result <= 12'b111111110101;
   48085: result <= 12'b111111110101;
   48086: result <= 12'b111111110101;
   48087: result <= 12'b111111110101;
   48088: result <= 12'b111111110101;
   48089: result <= 12'b111111110101;
   48090: result <= 12'b111111110101;
   48091: result <= 12'b111111110101;
   48092: result <= 12'b111111110101;
   48093: result <= 12'b111111110101;
   48094: result <= 12'b111111110101;
   48095: result <= 12'b111111110101;
   48096: result <= 12'b111111110101;
   48097: result <= 12'b111111110101;
   48098: result <= 12'b111111110101;
   48099: result <= 12'b111111110101;
   48100: result <= 12'b111111110101;
   48101: result <= 12'b111111110101;
   48102: result <= 12'b111111110101;
   48103: result <= 12'b111111110101;
   48104: result <= 12'b111111110101;
   48105: result <= 12'b111111110101;
   48106: result <= 12'b111111110101;
   48107: result <= 12'b111111110101;
   48108: result <= 12'b111111110101;
   48109: result <= 12'b111111110101;
   48110: result <= 12'b111111110101;
   48111: result <= 12'b111111110101;
   48112: result <= 12'b111111110101;
   48113: result <= 12'b111111110101;
   48114: result <= 12'b111111110101;
   48115: result <= 12'b111111110101;
   48116: result <= 12'b111111110101;
   48117: result <= 12'b111111110101;
   48118: result <= 12'b111111110101;
   48119: result <= 12'b111111110101;
   48120: result <= 12'b111111110101;
   48121: result <= 12'b111111110110;
   48122: result <= 12'b111111110110;
   48123: result <= 12'b111111110110;
   48124: result <= 12'b111111110110;
   48125: result <= 12'b111111110110;
   48126: result <= 12'b111111110110;
   48127: result <= 12'b111111110110;
   48128: result <= 12'b111111110110;
   48129: result <= 12'b111111110110;
   48130: result <= 12'b111111110110;
   48131: result <= 12'b111111110110;
   48132: result <= 12'b111111110110;
   48133: result <= 12'b111111110110;
   48134: result <= 12'b111111110110;
   48135: result <= 12'b111111110110;
   48136: result <= 12'b111111110110;
   48137: result <= 12'b111111110110;
   48138: result <= 12'b111111110110;
   48139: result <= 12'b111111110110;
   48140: result <= 12'b111111110110;
   48141: result <= 12'b111111110110;
   48142: result <= 12'b111111110110;
   48143: result <= 12'b111111110110;
   48144: result <= 12'b111111110110;
   48145: result <= 12'b111111110110;
   48146: result <= 12'b111111110110;
   48147: result <= 12'b111111110110;
   48148: result <= 12'b111111110110;
   48149: result <= 12'b111111110110;
   48150: result <= 12'b111111110110;
   48151: result <= 12'b111111110110;
   48152: result <= 12'b111111110110;
   48153: result <= 12'b111111110110;
   48154: result <= 12'b111111110110;
   48155: result <= 12'b111111110110;
   48156: result <= 12'b111111110110;
   48157: result <= 12'b111111110110;
   48158: result <= 12'b111111110110;
   48159: result <= 12'b111111110110;
   48160: result <= 12'b111111110110;
   48161: result <= 12'b111111110110;
   48162: result <= 12'b111111110110;
   48163: result <= 12'b111111110110;
   48164: result <= 12'b111111110110;
   48165: result <= 12'b111111110110;
   48166: result <= 12'b111111110110;
   48167: result <= 12'b111111110110;
   48168: result <= 12'b111111110110;
   48169: result <= 12'b111111110110;
   48170: result <= 12'b111111110110;
   48171: result <= 12'b111111110110;
   48172: result <= 12'b111111110110;
   48173: result <= 12'b111111110110;
   48174: result <= 12'b111111110111;
   48175: result <= 12'b111111110111;
   48176: result <= 12'b111111110111;
   48177: result <= 12'b111111110111;
   48178: result <= 12'b111111110111;
   48179: result <= 12'b111111110111;
   48180: result <= 12'b111111110111;
   48181: result <= 12'b111111110111;
   48182: result <= 12'b111111110111;
   48183: result <= 12'b111111110111;
   48184: result <= 12'b111111110111;
   48185: result <= 12'b111111110111;
   48186: result <= 12'b111111110111;
   48187: result <= 12'b111111110111;
   48188: result <= 12'b111111110111;
   48189: result <= 12'b111111110111;
   48190: result <= 12'b111111110111;
   48191: result <= 12'b111111110111;
   48192: result <= 12'b111111110111;
   48193: result <= 12'b111111110111;
   48194: result <= 12'b111111110111;
   48195: result <= 12'b111111110111;
   48196: result <= 12'b111111110111;
   48197: result <= 12'b111111110111;
   48198: result <= 12'b111111110111;
   48199: result <= 12'b111111110111;
   48200: result <= 12'b111111110111;
   48201: result <= 12'b111111110111;
   48202: result <= 12'b111111110111;
   48203: result <= 12'b111111110111;
   48204: result <= 12'b111111110111;
   48205: result <= 12'b111111110111;
   48206: result <= 12'b111111110111;
   48207: result <= 12'b111111110111;
   48208: result <= 12'b111111110111;
   48209: result <= 12'b111111110111;
   48210: result <= 12'b111111110111;
   48211: result <= 12'b111111110111;
   48212: result <= 12'b111111110111;
   48213: result <= 12'b111111110111;
   48214: result <= 12'b111111110111;
   48215: result <= 12'b111111110111;
   48216: result <= 12'b111111110111;
   48217: result <= 12'b111111110111;
   48218: result <= 12'b111111110111;
   48219: result <= 12'b111111110111;
   48220: result <= 12'b111111110111;
   48221: result <= 12'b111111110111;
   48222: result <= 12'b111111110111;
   48223: result <= 12'b111111110111;
   48224: result <= 12'b111111110111;
   48225: result <= 12'b111111110111;
   48226: result <= 12'b111111110111;
   48227: result <= 12'b111111110111;
   48228: result <= 12'b111111110111;
   48229: result <= 12'b111111110111;
   48230: result <= 12'b111111111000;
   48231: result <= 12'b111111111000;
   48232: result <= 12'b111111111000;
   48233: result <= 12'b111111111000;
   48234: result <= 12'b111111111000;
   48235: result <= 12'b111111111000;
   48236: result <= 12'b111111111000;
   48237: result <= 12'b111111111000;
   48238: result <= 12'b111111111000;
   48239: result <= 12'b111111111000;
   48240: result <= 12'b111111111000;
   48241: result <= 12'b111111111000;
   48242: result <= 12'b111111111000;
   48243: result <= 12'b111111111000;
   48244: result <= 12'b111111111000;
   48245: result <= 12'b111111111000;
   48246: result <= 12'b111111111000;
   48247: result <= 12'b111111111000;
   48248: result <= 12'b111111111000;
   48249: result <= 12'b111111111000;
   48250: result <= 12'b111111111000;
   48251: result <= 12'b111111111000;
   48252: result <= 12'b111111111000;
   48253: result <= 12'b111111111000;
   48254: result <= 12'b111111111000;
   48255: result <= 12'b111111111000;
   48256: result <= 12'b111111111000;
   48257: result <= 12'b111111111000;
   48258: result <= 12'b111111111000;
   48259: result <= 12'b111111111000;
   48260: result <= 12'b111111111000;
   48261: result <= 12'b111111111000;
   48262: result <= 12'b111111111000;
   48263: result <= 12'b111111111000;
   48264: result <= 12'b111111111000;
   48265: result <= 12'b111111111000;
   48266: result <= 12'b111111111000;
   48267: result <= 12'b111111111000;
   48268: result <= 12'b111111111000;
   48269: result <= 12'b111111111000;
   48270: result <= 12'b111111111000;
   48271: result <= 12'b111111111000;
   48272: result <= 12'b111111111000;
   48273: result <= 12'b111111111000;
   48274: result <= 12'b111111111000;
   48275: result <= 12'b111111111000;
   48276: result <= 12'b111111111000;
   48277: result <= 12'b111111111000;
   48278: result <= 12'b111111111000;
   48279: result <= 12'b111111111000;
   48280: result <= 12'b111111111000;
   48281: result <= 12'b111111111000;
   48282: result <= 12'b111111111000;
   48283: result <= 12'b111111111000;
   48284: result <= 12'b111111111000;
   48285: result <= 12'b111111111000;
   48286: result <= 12'b111111111000;
   48287: result <= 12'b111111111000;
   48288: result <= 12'b111111111000;
   48289: result <= 12'b111111111000;
   48290: result <= 12'b111111111001;
   48291: result <= 12'b111111111001;
   48292: result <= 12'b111111111001;
   48293: result <= 12'b111111111001;
   48294: result <= 12'b111111111001;
   48295: result <= 12'b111111111001;
   48296: result <= 12'b111111111001;
   48297: result <= 12'b111111111001;
   48298: result <= 12'b111111111001;
   48299: result <= 12'b111111111001;
   48300: result <= 12'b111111111001;
   48301: result <= 12'b111111111001;
   48302: result <= 12'b111111111001;
   48303: result <= 12'b111111111001;
   48304: result <= 12'b111111111001;
   48305: result <= 12'b111111111001;
   48306: result <= 12'b111111111001;
   48307: result <= 12'b111111111001;
   48308: result <= 12'b111111111001;
   48309: result <= 12'b111111111001;
   48310: result <= 12'b111111111001;
   48311: result <= 12'b111111111001;
   48312: result <= 12'b111111111001;
   48313: result <= 12'b111111111001;
   48314: result <= 12'b111111111001;
   48315: result <= 12'b111111111001;
   48316: result <= 12'b111111111001;
   48317: result <= 12'b111111111001;
   48318: result <= 12'b111111111001;
   48319: result <= 12'b111111111001;
   48320: result <= 12'b111111111001;
   48321: result <= 12'b111111111001;
   48322: result <= 12'b111111111001;
   48323: result <= 12'b111111111001;
   48324: result <= 12'b111111111001;
   48325: result <= 12'b111111111001;
   48326: result <= 12'b111111111001;
   48327: result <= 12'b111111111001;
   48328: result <= 12'b111111111001;
   48329: result <= 12'b111111111001;
   48330: result <= 12'b111111111001;
   48331: result <= 12'b111111111001;
   48332: result <= 12'b111111111001;
   48333: result <= 12'b111111111001;
   48334: result <= 12'b111111111001;
   48335: result <= 12'b111111111001;
   48336: result <= 12'b111111111001;
   48337: result <= 12'b111111111001;
   48338: result <= 12'b111111111001;
   48339: result <= 12'b111111111001;
   48340: result <= 12'b111111111001;
   48341: result <= 12'b111111111001;
   48342: result <= 12'b111111111001;
   48343: result <= 12'b111111111001;
   48344: result <= 12'b111111111001;
   48345: result <= 12'b111111111001;
   48346: result <= 12'b111111111001;
   48347: result <= 12'b111111111001;
   48348: result <= 12'b111111111001;
   48349: result <= 12'b111111111001;
   48350: result <= 12'b111111111001;
   48351: result <= 12'b111111111001;
   48352: result <= 12'b111111111001;
   48353: result <= 12'b111111111001;
   48354: result <= 12'b111111111010;
   48355: result <= 12'b111111111010;
   48356: result <= 12'b111111111010;
   48357: result <= 12'b111111111010;
   48358: result <= 12'b111111111010;
   48359: result <= 12'b111111111010;
   48360: result <= 12'b111111111010;
   48361: result <= 12'b111111111010;
   48362: result <= 12'b111111111010;
   48363: result <= 12'b111111111010;
   48364: result <= 12'b111111111010;
   48365: result <= 12'b111111111010;
   48366: result <= 12'b111111111010;
   48367: result <= 12'b111111111010;
   48368: result <= 12'b111111111010;
   48369: result <= 12'b111111111010;
   48370: result <= 12'b111111111010;
   48371: result <= 12'b111111111010;
   48372: result <= 12'b111111111010;
   48373: result <= 12'b111111111010;
   48374: result <= 12'b111111111010;
   48375: result <= 12'b111111111010;
   48376: result <= 12'b111111111010;
   48377: result <= 12'b111111111010;
   48378: result <= 12'b111111111010;
   48379: result <= 12'b111111111010;
   48380: result <= 12'b111111111010;
   48381: result <= 12'b111111111010;
   48382: result <= 12'b111111111010;
   48383: result <= 12'b111111111010;
   48384: result <= 12'b111111111010;
   48385: result <= 12'b111111111010;
   48386: result <= 12'b111111111010;
   48387: result <= 12'b111111111010;
   48388: result <= 12'b111111111010;
   48389: result <= 12'b111111111010;
   48390: result <= 12'b111111111010;
   48391: result <= 12'b111111111010;
   48392: result <= 12'b111111111010;
   48393: result <= 12'b111111111010;
   48394: result <= 12'b111111111010;
   48395: result <= 12'b111111111010;
   48396: result <= 12'b111111111010;
   48397: result <= 12'b111111111010;
   48398: result <= 12'b111111111010;
   48399: result <= 12'b111111111010;
   48400: result <= 12'b111111111010;
   48401: result <= 12'b111111111010;
   48402: result <= 12'b111111111010;
   48403: result <= 12'b111111111010;
   48404: result <= 12'b111111111010;
   48405: result <= 12'b111111111010;
   48406: result <= 12'b111111111010;
   48407: result <= 12'b111111111010;
   48408: result <= 12'b111111111010;
   48409: result <= 12'b111111111010;
   48410: result <= 12'b111111111010;
   48411: result <= 12'b111111111010;
   48412: result <= 12'b111111111010;
   48413: result <= 12'b111111111010;
   48414: result <= 12'b111111111010;
   48415: result <= 12'b111111111010;
   48416: result <= 12'b111111111010;
   48417: result <= 12'b111111111010;
   48418: result <= 12'b111111111010;
   48419: result <= 12'b111111111010;
   48420: result <= 12'b111111111010;
   48421: result <= 12'b111111111010;
   48422: result <= 12'b111111111010;
   48423: result <= 12'b111111111010;
   48424: result <= 12'b111111111011;
   48425: result <= 12'b111111111011;
   48426: result <= 12'b111111111011;
   48427: result <= 12'b111111111011;
   48428: result <= 12'b111111111011;
   48429: result <= 12'b111111111011;
   48430: result <= 12'b111111111011;
   48431: result <= 12'b111111111011;
   48432: result <= 12'b111111111011;
   48433: result <= 12'b111111111011;
   48434: result <= 12'b111111111011;
   48435: result <= 12'b111111111011;
   48436: result <= 12'b111111111011;
   48437: result <= 12'b111111111011;
   48438: result <= 12'b111111111011;
   48439: result <= 12'b111111111011;
   48440: result <= 12'b111111111011;
   48441: result <= 12'b111111111011;
   48442: result <= 12'b111111111011;
   48443: result <= 12'b111111111011;
   48444: result <= 12'b111111111011;
   48445: result <= 12'b111111111011;
   48446: result <= 12'b111111111011;
   48447: result <= 12'b111111111011;
   48448: result <= 12'b111111111011;
   48449: result <= 12'b111111111011;
   48450: result <= 12'b111111111011;
   48451: result <= 12'b111111111011;
   48452: result <= 12'b111111111011;
   48453: result <= 12'b111111111011;
   48454: result <= 12'b111111111011;
   48455: result <= 12'b111111111011;
   48456: result <= 12'b111111111011;
   48457: result <= 12'b111111111011;
   48458: result <= 12'b111111111011;
   48459: result <= 12'b111111111011;
   48460: result <= 12'b111111111011;
   48461: result <= 12'b111111111011;
   48462: result <= 12'b111111111011;
   48463: result <= 12'b111111111011;
   48464: result <= 12'b111111111011;
   48465: result <= 12'b111111111011;
   48466: result <= 12'b111111111011;
   48467: result <= 12'b111111111011;
   48468: result <= 12'b111111111011;
   48469: result <= 12'b111111111011;
   48470: result <= 12'b111111111011;
   48471: result <= 12'b111111111011;
   48472: result <= 12'b111111111011;
   48473: result <= 12'b111111111011;
   48474: result <= 12'b111111111011;
   48475: result <= 12'b111111111011;
   48476: result <= 12'b111111111011;
   48477: result <= 12'b111111111011;
   48478: result <= 12'b111111111011;
   48479: result <= 12'b111111111011;
   48480: result <= 12'b111111111011;
   48481: result <= 12'b111111111011;
   48482: result <= 12'b111111111011;
   48483: result <= 12'b111111111011;
   48484: result <= 12'b111111111011;
   48485: result <= 12'b111111111011;
   48486: result <= 12'b111111111011;
   48487: result <= 12'b111111111011;
   48488: result <= 12'b111111111011;
   48489: result <= 12'b111111111011;
   48490: result <= 12'b111111111011;
   48491: result <= 12'b111111111011;
   48492: result <= 12'b111111111011;
   48493: result <= 12'b111111111011;
   48494: result <= 12'b111111111011;
   48495: result <= 12'b111111111011;
   48496: result <= 12'b111111111011;
   48497: result <= 12'b111111111011;
   48498: result <= 12'b111111111011;
   48499: result <= 12'b111111111011;
   48500: result <= 12'b111111111100;
   48501: result <= 12'b111111111100;
   48502: result <= 12'b111111111100;
   48503: result <= 12'b111111111100;
   48504: result <= 12'b111111111100;
   48505: result <= 12'b111111111100;
   48506: result <= 12'b111111111100;
   48507: result <= 12'b111111111100;
   48508: result <= 12'b111111111100;
   48509: result <= 12'b111111111100;
   48510: result <= 12'b111111111100;
   48511: result <= 12'b111111111100;
   48512: result <= 12'b111111111100;
   48513: result <= 12'b111111111100;
   48514: result <= 12'b111111111100;
   48515: result <= 12'b111111111100;
   48516: result <= 12'b111111111100;
   48517: result <= 12'b111111111100;
   48518: result <= 12'b111111111100;
   48519: result <= 12'b111111111100;
   48520: result <= 12'b111111111100;
   48521: result <= 12'b111111111100;
   48522: result <= 12'b111111111100;
   48523: result <= 12'b111111111100;
   48524: result <= 12'b111111111100;
   48525: result <= 12'b111111111100;
   48526: result <= 12'b111111111100;
   48527: result <= 12'b111111111100;
   48528: result <= 12'b111111111100;
   48529: result <= 12'b111111111100;
   48530: result <= 12'b111111111100;
   48531: result <= 12'b111111111100;
   48532: result <= 12'b111111111100;
   48533: result <= 12'b111111111100;
   48534: result <= 12'b111111111100;
   48535: result <= 12'b111111111100;
   48536: result <= 12'b111111111100;
   48537: result <= 12'b111111111100;
   48538: result <= 12'b111111111100;
   48539: result <= 12'b111111111100;
   48540: result <= 12'b111111111100;
   48541: result <= 12'b111111111100;
   48542: result <= 12'b111111111100;
   48543: result <= 12'b111111111100;
   48544: result <= 12'b111111111100;
   48545: result <= 12'b111111111100;
   48546: result <= 12'b111111111100;
   48547: result <= 12'b111111111100;
   48548: result <= 12'b111111111100;
   48549: result <= 12'b111111111100;
   48550: result <= 12'b111111111100;
   48551: result <= 12'b111111111100;
   48552: result <= 12'b111111111100;
   48553: result <= 12'b111111111100;
   48554: result <= 12'b111111111100;
   48555: result <= 12'b111111111100;
   48556: result <= 12'b111111111100;
   48557: result <= 12'b111111111100;
   48558: result <= 12'b111111111100;
   48559: result <= 12'b111111111100;
   48560: result <= 12'b111111111100;
   48561: result <= 12'b111111111100;
   48562: result <= 12'b111111111100;
   48563: result <= 12'b111111111100;
   48564: result <= 12'b111111111100;
   48565: result <= 12'b111111111100;
   48566: result <= 12'b111111111100;
   48567: result <= 12'b111111111100;
   48568: result <= 12'b111111111100;
   48569: result <= 12'b111111111100;
   48570: result <= 12'b111111111100;
   48571: result <= 12'b111111111100;
   48572: result <= 12'b111111111100;
   48573: result <= 12'b111111111100;
   48574: result <= 12'b111111111100;
   48575: result <= 12'b111111111100;
   48576: result <= 12'b111111111100;
   48577: result <= 12'b111111111100;
   48578: result <= 12'b111111111100;
   48579: result <= 12'b111111111100;
   48580: result <= 12'b111111111100;
   48581: result <= 12'b111111111100;
   48582: result <= 12'b111111111100;
   48583: result <= 12'b111111111100;
   48584: result <= 12'b111111111100;
   48585: result <= 12'b111111111100;
   48586: result <= 12'b111111111100;
   48587: result <= 12'b111111111100;
   48588: result <= 12'b111111111101;
   48589: result <= 12'b111111111101;
   48590: result <= 12'b111111111101;
   48591: result <= 12'b111111111101;
   48592: result <= 12'b111111111101;
   48593: result <= 12'b111111111101;
   48594: result <= 12'b111111111101;
   48595: result <= 12'b111111111101;
   48596: result <= 12'b111111111101;
   48597: result <= 12'b111111111101;
   48598: result <= 12'b111111111101;
   48599: result <= 12'b111111111101;
   48600: result <= 12'b111111111101;
   48601: result <= 12'b111111111101;
   48602: result <= 12'b111111111101;
   48603: result <= 12'b111111111101;
   48604: result <= 12'b111111111101;
   48605: result <= 12'b111111111101;
   48606: result <= 12'b111111111101;
   48607: result <= 12'b111111111101;
   48608: result <= 12'b111111111101;
   48609: result <= 12'b111111111101;
   48610: result <= 12'b111111111101;
   48611: result <= 12'b111111111101;
   48612: result <= 12'b111111111101;
   48613: result <= 12'b111111111101;
   48614: result <= 12'b111111111101;
   48615: result <= 12'b111111111101;
   48616: result <= 12'b111111111101;
   48617: result <= 12'b111111111101;
   48618: result <= 12'b111111111101;
   48619: result <= 12'b111111111101;
   48620: result <= 12'b111111111101;
   48621: result <= 12'b111111111101;
   48622: result <= 12'b111111111101;
   48623: result <= 12'b111111111101;
   48624: result <= 12'b111111111101;
   48625: result <= 12'b111111111101;
   48626: result <= 12'b111111111101;
   48627: result <= 12'b111111111101;
   48628: result <= 12'b111111111101;
   48629: result <= 12'b111111111101;
   48630: result <= 12'b111111111101;
   48631: result <= 12'b111111111101;
   48632: result <= 12'b111111111101;
   48633: result <= 12'b111111111101;
   48634: result <= 12'b111111111101;
   48635: result <= 12'b111111111101;
   48636: result <= 12'b111111111101;
   48637: result <= 12'b111111111101;
   48638: result <= 12'b111111111101;
   48639: result <= 12'b111111111101;
   48640: result <= 12'b111111111101;
   48641: result <= 12'b111111111101;
   48642: result <= 12'b111111111101;
   48643: result <= 12'b111111111101;
   48644: result <= 12'b111111111101;
   48645: result <= 12'b111111111101;
   48646: result <= 12'b111111111101;
   48647: result <= 12'b111111111101;
   48648: result <= 12'b111111111101;
   48649: result <= 12'b111111111101;
   48650: result <= 12'b111111111101;
   48651: result <= 12'b111111111101;
   48652: result <= 12'b111111111101;
   48653: result <= 12'b111111111101;
   48654: result <= 12'b111111111101;
   48655: result <= 12'b111111111101;
   48656: result <= 12'b111111111101;
   48657: result <= 12'b111111111101;
   48658: result <= 12'b111111111101;
   48659: result <= 12'b111111111101;
   48660: result <= 12'b111111111101;
   48661: result <= 12'b111111111101;
   48662: result <= 12'b111111111101;
   48663: result <= 12'b111111111101;
   48664: result <= 12'b111111111101;
   48665: result <= 12'b111111111101;
   48666: result <= 12'b111111111101;
   48667: result <= 12'b111111111101;
   48668: result <= 12'b111111111101;
   48669: result <= 12'b111111111101;
   48670: result <= 12'b111111111101;
   48671: result <= 12'b111111111101;
   48672: result <= 12'b111111111101;
   48673: result <= 12'b111111111101;
   48674: result <= 12'b111111111101;
   48675: result <= 12'b111111111101;
   48676: result <= 12'b111111111101;
   48677: result <= 12'b111111111101;
   48678: result <= 12'b111111111101;
   48679: result <= 12'b111111111101;
   48680: result <= 12'b111111111101;
   48681: result <= 12'b111111111101;
   48682: result <= 12'b111111111101;
   48683: result <= 12'b111111111101;
   48684: result <= 12'b111111111101;
   48685: result <= 12'b111111111101;
   48686: result <= 12'b111111111101;
   48687: result <= 12'b111111111101;
   48688: result <= 12'b111111111101;
   48689: result <= 12'b111111111101;
   48690: result <= 12'b111111111101;
   48691: result <= 12'b111111111101;
   48692: result <= 12'b111111111110;
   48693: result <= 12'b111111111110;
   48694: result <= 12'b111111111110;
   48695: result <= 12'b111111111110;
   48696: result <= 12'b111111111110;
   48697: result <= 12'b111111111110;
   48698: result <= 12'b111111111110;
   48699: result <= 12'b111111111110;
   48700: result <= 12'b111111111110;
   48701: result <= 12'b111111111110;
   48702: result <= 12'b111111111110;
   48703: result <= 12'b111111111110;
   48704: result <= 12'b111111111110;
   48705: result <= 12'b111111111110;
   48706: result <= 12'b111111111110;
   48707: result <= 12'b111111111110;
   48708: result <= 12'b111111111110;
   48709: result <= 12'b111111111110;
   48710: result <= 12'b111111111110;
   48711: result <= 12'b111111111110;
   48712: result <= 12'b111111111110;
   48713: result <= 12'b111111111110;
   48714: result <= 12'b111111111110;
   48715: result <= 12'b111111111110;
   48716: result <= 12'b111111111110;
   48717: result <= 12'b111111111110;
   48718: result <= 12'b111111111110;
   48719: result <= 12'b111111111110;
   48720: result <= 12'b111111111110;
   48721: result <= 12'b111111111110;
   48722: result <= 12'b111111111110;
   48723: result <= 12'b111111111110;
   48724: result <= 12'b111111111110;
   48725: result <= 12'b111111111110;
   48726: result <= 12'b111111111110;
   48727: result <= 12'b111111111110;
   48728: result <= 12'b111111111110;
   48729: result <= 12'b111111111110;
   48730: result <= 12'b111111111110;
   48731: result <= 12'b111111111110;
   48732: result <= 12'b111111111110;
   48733: result <= 12'b111111111110;
   48734: result <= 12'b111111111110;
   48735: result <= 12'b111111111110;
   48736: result <= 12'b111111111110;
   48737: result <= 12'b111111111110;
   48738: result <= 12'b111111111110;
   48739: result <= 12'b111111111110;
   48740: result <= 12'b111111111110;
   48741: result <= 12'b111111111110;
   48742: result <= 12'b111111111110;
   48743: result <= 12'b111111111110;
   48744: result <= 12'b111111111110;
   48745: result <= 12'b111111111110;
   48746: result <= 12'b111111111110;
   48747: result <= 12'b111111111110;
   48748: result <= 12'b111111111110;
   48749: result <= 12'b111111111110;
   48750: result <= 12'b111111111110;
   48751: result <= 12'b111111111110;
   48752: result <= 12'b111111111110;
   48753: result <= 12'b111111111110;
   48754: result <= 12'b111111111110;
   48755: result <= 12'b111111111110;
   48756: result <= 12'b111111111110;
   48757: result <= 12'b111111111110;
   48758: result <= 12'b111111111110;
   48759: result <= 12'b111111111110;
   48760: result <= 12'b111111111110;
   48761: result <= 12'b111111111110;
   48762: result <= 12'b111111111110;
   48763: result <= 12'b111111111110;
   48764: result <= 12'b111111111110;
   48765: result <= 12'b111111111110;
   48766: result <= 12'b111111111110;
   48767: result <= 12'b111111111110;
   48768: result <= 12'b111111111110;
   48769: result <= 12'b111111111110;
   48770: result <= 12'b111111111110;
   48771: result <= 12'b111111111110;
   48772: result <= 12'b111111111110;
   48773: result <= 12'b111111111110;
   48774: result <= 12'b111111111110;
   48775: result <= 12'b111111111110;
   48776: result <= 12'b111111111110;
   48777: result <= 12'b111111111110;
   48778: result <= 12'b111111111110;
   48779: result <= 12'b111111111110;
   48780: result <= 12'b111111111110;
   48781: result <= 12'b111111111110;
   48782: result <= 12'b111111111110;
   48783: result <= 12'b111111111110;
   48784: result <= 12'b111111111110;
   48785: result <= 12'b111111111110;
   48786: result <= 12'b111111111110;
   48787: result <= 12'b111111111110;
   48788: result <= 12'b111111111110;
   48789: result <= 12'b111111111110;
   48790: result <= 12'b111111111110;
   48791: result <= 12'b111111111110;
   48792: result <= 12'b111111111110;
   48793: result <= 12'b111111111110;
   48794: result <= 12'b111111111110;
   48795: result <= 12'b111111111110;
   48796: result <= 12'b111111111110;
   48797: result <= 12'b111111111110;
   48798: result <= 12'b111111111110;
   48799: result <= 12'b111111111110;
   48800: result <= 12'b111111111110;
   48801: result <= 12'b111111111110;
   48802: result <= 12'b111111111110;
   48803: result <= 12'b111111111110;
   48804: result <= 12'b111111111110;
   48805: result <= 12'b111111111110;
   48806: result <= 12'b111111111110;
   48807: result <= 12'b111111111110;
   48808: result <= 12'b111111111110;
   48809: result <= 12'b111111111110;
   48810: result <= 12'b111111111110;
   48811: result <= 12'b111111111110;
   48812: result <= 12'b111111111110;
   48813: result <= 12'b111111111110;
   48814: result <= 12'b111111111110;
   48815: result <= 12'b111111111110;
   48816: result <= 12'b111111111110;
   48817: result <= 12'b111111111110;
   48818: result <= 12'b111111111110;
   48819: result <= 12'b111111111110;
   48820: result <= 12'b111111111110;
   48821: result <= 12'b111111111110;
   48822: result <= 12'b111111111110;
   48823: result <= 12'b111111111110;
   48824: result <= 12'b111111111110;
   48825: result <= 12'b111111111110;
   48826: result <= 12'b111111111110;
   48827: result <= 12'b111111111111;
   48828: result <= 12'b111111111111;
   48829: result <= 12'b111111111111;
   48830: result <= 12'b111111111111;
   48831: result <= 12'b111111111111;
   48832: result <= 12'b111111111111;
   48833: result <= 12'b111111111111;
   48834: result <= 12'b111111111111;
   48835: result <= 12'b111111111111;
   48836: result <= 12'b111111111111;
   48837: result <= 12'b111111111111;
   48838: result <= 12'b111111111111;
   48839: result <= 12'b111111111111;
   48840: result <= 12'b111111111111;
   48841: result <= 12'b111111111111;
   48842: result <= 12'b111111111111;
   48843: result <= 12'b111111111111;
   48844: result <= 12'b111111111111;
   48845: result <= 12'b111111111111;
   48846: result <= 12'b111111111111;
   48847: result <= 12'b111111111111;
   48848: result <= 12'b111111111111;
   48849: result <= 12'b111111111111;
   48850: result <= 12'b111111111111;
   48851: result <= 12'b111111111111;
   48852: result <= 12'b111111111111;
   48853: result <= 12'b111111111111;
   48854: result <= 12'b111111111111;
   48855: result <= 12'b111111111111;
   48856: result <= 12'b111111111111;
   48857: result <= 12'b111111111111;
   48858: result <= 12'b111111111111;
   48859: result <= 12'b111111111111;
   48860: result <= 12'b111111111111;
   48861: result <= 12'b111111111111;
   48862: result <= 12'b111111111111;
   48863: result <= 12'b111111111111;
   48864: result <= 12'b111111111111;
   48865: result <= 12'b111111111111;
   48866: result <= 12'b111111111111;
   48867: result <= 12'b111111111111;
   48868: result <= 12'b111111111111;
   48869: result <= 12'b111111111111;
   48870: result <= 12'b111111111111;
   48871: result <= 12'b111111111111;
   48872: result <= 12'b111111111111;
   48873: result <= 12'b111111111111;
   48874: result <= 12'b111111111111;
   48875: result <= 12'b111111111111;
   48876: result <= 12'b111111111111;
   48877: result <= 12'b111111111111;
   48878: result <= 12'b111111111111;
   48879: result <= 12'b111111111111;
   48880: result <= 12'b111111111111;
   48881: result <= 12'b111111111111;
   48882: result <= 12'b111111111111;
   48883: result <= 12'b111111111111;
   48884: result <= 12'b111111111111;
   48885: result <= 12'b111111111111;
   48886: result <= 12'b111111111111;
   48887: result <= 12'b111111111111;
   48888: result <= 12'b111111111111;
   48889: result <= 12'b111111111111;
   48890: result <= 12'b111111111111;
   48891: result <= 12'b111111111111;
   48892: result <= 12'b111111111111;
   48893: result <= 12'b111111111111;
   48894: result <= 12'b111111111111;
   48895: result <= 12'b111111111111;
   48896: result <= 12'b111111111111;
   48897: result <= 12'b111111111111;
   48898: result <= 12'b111111111111;
   48899: result <= 12'b111111111111;
   48900: result <= 12'b111111111111;
   48901: result <= 12'b111111111111;
   48902: result <= 12'b111111111111;
   48903: result <= 12'b111111111111;
   48904: result <= 12'b111111111111;
   48905: result <= 12'b111111111111;
   48906: result <= 12'b111111111111;
   48907: result <= 12'b111111111111;
   48908: result <= 12'b111111111111;
   48909: result <= 12'b111111111111;
   48910: result <= 12'b111111111111;
   48911: result <= 12'b111111111111;
   48912: result <= 12'b111111111111;
   48913: result <= 12'b111111111111;
   48914: result <= 12'b111111111111;
   48915: result <= 12'b111111111111;
   48916: result <= 12'b111111111111;
   48917: result <= 12'b111111111111;
   48918: result <= 12'b111111111111;
   48919: result <= 12'b111111111111;
   48920: result <= 12'b111111111111;
   48921: result <= 12'b111111111111;
   48922: result <= 12'b111111111111;
   48923: result <= 12'b111111111111;
   48924: result <= 12'b111111111111;
   48925: result <= 12'b111111111111;
   48926: result <= 12'b111111111111;
   48927: result <= 12'b111111111111;
   48928: result <= 12'b111111111111;
   48929: result <= 12'b111111111111;
   48930: result <= 12'b111111111111;
   48931: result <= 12'b111111111111;
   48932: result <= 12'b111111111111;
   48933: result <= 12'b111111111111;
   48934: result <= 12'b111111111111;
   48935: result <= 12'b111111111111;
   48936: result <= 12'b111111111111;
   48937: result <= 12'b111111111111;
   48938: result <= 12'b111111111111;
   48939: result <= 12'b111111111111;
   48940: result <= 12'b111111111111;
   48941: result <= 12'b111111111111;
   48942: result <= 12'b111111111111;
   48943: result <= 12'b111111111111;
   48944: result <= 12'b111111111111;
   48945: result <= 12'b111111111111;
   48946: result <= 12'b111111111111;
   48947: result <= 12'b111111111111;
   48948: result <= 12'b111111111111;
   48949: result <= 12'b111111111111;
   48950: result <= 12'b111111111111;
   48951: result <= 12'b111111111111;
   48952: result <= 12'b111111111111;
   48953: result <= 12'b111111111111;
   48954: result <= 12'b111111111111;
   48955: result <= 12'b111111111111;
   48956: result <= 12'b111111111111;
   48957: result <= 12'b111111111111;
   48958: result <= 12'b111111111111;
   48959: result <= 12'b111111111111;
   48960: result <= 12'b111111111111;
   48961: result <= 12'b111111111111;
   48962: result <= 12'b111111111111;
   48963: result <= 12'b111111111111;
   48964: result <= 12'b111111111111;
   48965: result <= 12'b111111111111;
   48966: result <= 12'b111111111111;
   48967: result <= 12'b111111111111;
   48968: result <= 12'b111111111111;
   48969: result <= 12'b111111111111;
   48970: result <= 12'b111111111111;
   48971: result <= 12'b111111111111;
   48972: result <= 12'b111111111111;
   48973: result <= 12'b111111111111;
   48974: result <= 12'b111111111111;
   48975: result <= 12'b111111111111;
   48976: result <= 12'b111111111111;
   48977: result <= 12'b111111111111;
   48978: result <= 12'b111111111111;
   48979: result <= 12'b111111111111;
   48980: result <= 12'b111111111111;
   48981: result <= 12'b111111111111;
   48982: result <= 12'b111111111111;
   48983: result <= 12'b111111111111;
   48984: result <= 12'b111111111111;
   48985: result <= 12'b111111111111;
   48986: result <= 12'b111111111111;
   48987: result <= 12'b111111111111;
   48988: result <= 12'b111111111111;
   48989: result <= 12'b111111111111;
   48990: result <= 12'b111111111111;
   48991: result <= 12'b111111111111;
   48992: result <= 12'b111111111111;
   48993: result <= 12'b111111111111;
   48994: result <= 12'b111111111111;
   48995: result <= 12'b111111111111;
   48996: result <= 12'b111111111111;
   48997: result <= 12'b111111111111;
   48998: result <= 12'b111111111111;
   48999: result <= 12'b111111111111;
   49000: result <= 12'b111111111111;
   49001: result <= 12'b111111111111;
   49002: result <= 12'b111111111111;
   49003: result <= 12'b111111111111;
   49004: result <= 12'b111111111111;
   49005: result <= 12'b111111111111;
   49006: result <= 12'b111111111111;
   49007: result <= 12'b111111111111;
   49008: result <= 12'b111111111111;
   49009: result <= 12'b111111111111;
   49010: result <= 12'b111111111111;
   49011: result <= 12'b111111111111;
   49012: result <= 12'b111111111111;
   49013: result <= 12'b111111111111;
   49014: result <= 12'b111111111111;
   49015: result <= 12'b111111111111;
   49016: result <= 12'b111111111111;
   49017: result <= 12'b111111111111;
   49018: result <= 12'b111111111111;
   49019: result <= 12'b111111111111;
   49020: result <= 12'b111111111111;
   49021: result <= 12'b111111111111;
   49022: result <= 12'b111111111111;
   49023: result <= 12'b111111111111;
   49024: result <= 12'b111111111111;
   49025: result <= 12'b111111111111;
   49026: result <= 12'b111111111111;
   49027: result <= 12'b111111111111;
   49028: result <= 12'b111111111111;
   49029: result <= 12'b111111111111;
   49030: result <= 12'b111111111111;
   49031: result <= 12'b111111111111;
   49032: result <= 12'b111111111111;
   49033: result <= 12'b111111111111;
   49034: result <= 12'b111111111111;
   49035: result <= 12'b111111111111;
   49036: result <= 12'b111111111111;
   49037: result <= 12'b111111111111;
   49038: result <= 12'b111111111111;
   49039: result <= 12'b111111111111;
   49040: result <= 12'b111111111111;
   49041: result <= 12'b111111111111;
   49042: result <= 12'b111111111111;
   49043: result <= 12'b111111111111;
   49044: result <= 12'b111111111111;
   49045: result <= 12'b111111111111;
   49046: result <= 12'b111111111111;
   49047: result <= 12'b111111111111;
   49048: result <= 12'b111111111111;
   49049: result <= 12'b111111111111;
   49050: result <= 12'b111111111111;
   49051: result <= 12'b111111111111;
   49052: result <= 12'b111111111111;
   49053: result <= 12'b111111111111;
   49054: result <= 12'b111111111111;
   49055: result <= 12'b111111111111;
   49056: result <= 12'b111111111111;
   49057: result <= 12'b111111111111;
   49058: result <= 12'b111111111111;
   49059: result <= 12'b111111111111;
   49060: result <= 12'b111111111111;
   49061: result <= 12'b111111111111;
   49062: result <= 12'b111111111111;
   49063: result <= 12'b111111111111;
   49064: result <= 12'b111111111111;
   49065: result <= 12'b111111111111;
   49066: result <= 12'b111111111111;
   49067: result <= 12'b111111111111;
   49068: result <= 12'b111111111111;
   49069: result <= 12'b111111111111;
   49070: result <= 12'b111111111111;
   49071: result <= 12'b111111111111;
   49072: result <= 12'b111111111111;
   49073: result <= 12'b111111111111;
   49074: result <= 12'b111111111111;
   49075: result <= 12'b111111111111;
   49076: result <= 12'b111111111111;
   49077: result <= 12'b111111111111;
   49078: result <= 12'b111111111111;
   49079: result <= 12'b111111111111;
   49080: result <= 12'b111111111111;
   49081: result <= 12'b111111111111;
   49082: result <= 12'b111111111111;
   49083: result <= 12'b111111111111;
   49084: result <= 12'b111111111111;
   49085: result <= 12'b111111111111;
   49086: result <= 12'b111111111111;
   49087: result <= 12'b111111111111;
   49088: result <= 12'b111111111111;
   49089: result <= 12'b111111111111;
   49090: result <= 12'b111111111111;
   49091: result <= 12'b111111111111;
   49092: result <= 12'b111111111111;
   49093: result <= 12'b111111111111;
   49094: result <= 12'b111111111111;
   49095: result <= 12'b111111111111;
   49096: result <= 12'b111111111111;
   49097: result <= 12'b111111111111;
   49098: result <= 12'b111111111111;
   49099: result <= 12'b111111111111;
   49100: result <= 12'b111111111111;
   49101: result <= 12'b111111111111;
   49102: result <= 12'b111111111111;
   49103: result <= 12'b111111111111;
   49104: result <= 12'b111111111111;
   49105: result <= 12'b111111111111;
   49106: result <= 12'b111111111111;
   49107: result <= 12'b111111111111;
   49108: result <= 12'b111111111111;
   49109: result <= 12'b111111111111;
   49110: result <= 12'b111111111111;
   49111: result <= 12'b111111111111;
   49112: result <= 12'b111111111111;
   49113: result <= 12'b111111111111;
   49114: result <= 12'b111111111111;
   49115: result <= 12'b111111111111;
   49116: result <= 12'b111111111111;
   49117: result <= 12'b111111111111;
   49118: result <= 12'b111111111111;
   49119: result <= 12'b111111111111;
   49120: result <= 12'b111111111111;
   49121: result <= 12'b111111111111;
   49122: result <= 12'b111111111111;
   49123: result <= 12'b111111111111;
   49124: result <= 12'b111111111111;
   49125: result <= 12'b111111111111;
   49126: result <= 12'b111111111111;
   49127: result <= 12'b111111111111;
   49128: result <= 12'b111111111111;
   49129: result <= 12'b111111111111;
   49130: result <= 12'b111111111111;
   49131: result <= 12'b111111111111;
   49132: result <= 12'b111111111111;
   49133: result <= 12'b111111111111;
   49134: result <= 12'b111111111111;
   49135: result <= 12'b111111111111;
   49136: result <= 12'b111111111111;
   49137: result <= 12'b111111111111;
   49138: result <= 12'b111111111111;
   49139: result <= 12'b111111111111;
   49140: result <= 12'b111111111111;
   49141: result <= 12'b111111111111;
   49142: result <= 12'b111111111111;
   49143: result <= 12'b111111111111;
   49144: result <= 12'b111111111111;
   49145: result <= 12'b111111111111;
   49146: result <= 12'b111111111111;
   49147: result <= 12'b111111111111;
   49148: result <= 12'b111111111111;
   49149: result <= 12'b111111111111;
   49150: result <= 12'b111111111111;
   49151: result <= 12'b111111111111;
   49152: result <= 12'b100000000000;
   49153: result <= 12'b111111111111;
   49154: result <= 12'b111111111111;
   49155: result <= 12'b111111111111;
   49156: result <= 12'b111111111111;
   49157: result <= 12'b111111111111;
   49158: result <= 12'b111111111111;
   49159: result <= 12'b111111111111;
   49160: result <= 12'b111111111111;
   49161: result <= 12'b111111111111;
   49162: result <= 12'b111111111111;
   49163: result <= 12'b111111111111;
   49164: result <= 12'b111111111111;
   49165: result <= 12'b111111111111;
   49166: result <= 12'b111111111111;
   49167: result <= 12'b111111111111;
   49168: result <= 12'b111111111111;
   49169: result <= 12'b111111111111;
   49170: result <= 12'b111111111111;
   49171: result <= 12'b111111111111;
   49172: result <= 12'b111111111111;
   49173: result <= 12'b111111111111;
   49174: result <= 12'b111111111111;
   49175: result <= 12'b111111111111;
   49176: result <= 12'b111111111111;
   49177: result <= 12'b111111111111;
   49178: result <= 12'b111111111111;
   49179: result <= 12'b111111111111;
   49180: result <= 12'b111111111111;
   49181: result <= 12'b111111111111;
   49182: result <= 12'b111111111111;
   49183: result <= 12'b111111111111;
   49184: result <= 12'b111111111111;
   49185: result <= 12'b111111111111;
   49186: result <= 12'b111111111111;
   49187: result <= 12'b111111111111;
   49188: result <= 12'b111111111111;
   49189: result <= 12'b111111111111;
   49190: result <= 12'b111111111111;
   49191: result <= 12'b111111111111;
   49192: result <= 12'b111111111111;
   49193: result <= 12'b111111111111;
   49194: result <= 12'b111111111111;
   49195: result <= 12'b111111111111;
   49196: result <= 12'b111111111111;
   49197: result <= 12'b111111111111;
   49198: result <= 12'b111111111111;
   49199: result <= 12'b111111111111;
   49200: result <= 12'b111111111111;
   49201: result <= 12'b111111111111;
   49202: result <= 12'b111111111111;
   49203: result <= 12'b111111111111;
   49204: result <= 12'b111111111111;
   49205: result <= 12'b111111111111;
   49206: result <= 12'b111111111111;
   49207: result <= 12'b111111111111;
   49208: result <= 12'b111111111111;
   49209: result <= 12'b111111111111;
   49210: result <= 12'b111111111111;
   49211: result <= 12'b111111111111;
   49212: result <= 12'b111111111111;
   49213: result <= 12'b111111111111;
   49214: result <= 12'b111111111111;
   49215: result <= 12'b111111111111;
   49216: result <= 12'b111111111111;
   49217: result <= 12'b111111111111;
   49218: result <= 12'b111111111111;
   49219: result <= 12'b111111111111;
   49220: result <= 12'b111111111111;
   49221: result <= 12'b111111111111;
   49222: result <= 12'b111111111111;
   49223: result <= 12'b111111111111;
   49224: result <= 12'b111111111111;
   49225: result <= 12'b111111111111;
   49226: result <= 12'b111111111111;
   49227: result <= 12'b111111111111;
   49228: result <= 12'b111111111111;
   49229: result <= 12'b111111111111;
   49230: result <= 12'b111111111111;
   49231: result <= 12'b111111111111;
   49232: result <= 12'b111111111111;
   49233: result <= 12'b111111111111;
   49234: result <= 12'b111111111111;
   49235: result <= 12'b111111111111;
   49236: result <= 12'b111111111111;
   49237: result <= 12'b111111111111;
   49238: result <= 12'b111111111111;
   49239: result <= 12'b111111111111;
   49240: result <= 12'b111111111111;
   49241: result <= 12'b111111111111;
   49242: result <= 12'b111111111111;
   49243: result <= 12'b111111111111;
   49244: result <= 12'b111111111111;
   49245: result <= 12'b111111111111;
   49246: result <= 12'b111111111111;
   49247: result <= 12'b111111111111;
   49248: result <= 12'b111111111111;
   49249: result <= 12'b111111111111;
   49250: result <= 12'b111111111111;
   49251: result <= 12'b111111111111;
   49252: result <= 12'b111111111111;
   49253: result <= 12'b111111111111;
   49254: result <= 12'b111111111111;
   49255: result <= 12'b111111111111;
   49256: result <= 12'b111111111111;
   49257: result <= 12'b111111111111;
   49258: result <= 12'b111111111111;
   49259: result <= 12'b111111111111;
   49260: result <= 12'b111111111111;
   49261: result <= 12'b111111111111;
   49262: result <= 12'b111111111111;
   49263: result <= 12'b111111111111;
   49264: result <= 12'b111111111111;
   49265: result <= 12'b111111111111;
   49266: result <= 12'b111111111111;
   49267: result <= 12'b111111111111;
   49268: result <= 12'b111111111111;
   49269: result <= 12'b111111111111;
   49270: result <= 12'b111111111111;
   49271: result <= 12'b111111111111;
   49272: result <= 12'b111111111111;
   49273: result <= 12'b111111111111;
   49274: result <= 12'b111111111111;
   49275: result <= 12'b111111111111;
   49276: result <= 12'b111111111111;
   49277: result <= 12'b111111111111;
   49278: result <= 12'b111111111111;
   49279: result <= 12'b111111111111;
   49280: result <= 12'b111111111111;
   49281: result <= 12'b111111111111;
   49282: result <= 12'b111111111111;
   49283: result <= 12'b111111111111;
   49284: result <= 12'b111111111111;
   49285: result <= 12'b111111111111;
   49286: result <= 12'b111111111111;
   49287: result <= 12'b111111111111;
   49288: result <= 12'b111111111111;
   49289: result <= 12'b111111111111;
   49290: result <= 12'b111111111111;
   49291: result <= 12'b111111111111;
   49292: result <= 12'b111111111111;
   49293: result <= 12'b111111111111;
   49294: result <= 12'b111111111111;
   49295: result <= 12'b111111111111;
   49296: result <= 12'b111111111111;
   49297: result <= 12'b111111111111;
   49298: result <= 12'b111111111111;
   49299: result <= 12'b111111111111;
   49300: result <= 12'b111111111111;
   49301: result <= 12'b111111111111;
   49302: result <= 12'b111111111111;
   49303: result <= 12'b111111111111;
   49304: result <= 12'b111111111111;
   49305: result <= 12'b111111111111;
   49306: result <= 12'b111111111111;
   49307: result <= 12'b111111111111;
   49308: result <= 12'b111111111111;
   49309: result <= 12'b111111111111;
   49310: result <= 12'b111111111111;
   49311: result <= 12'b111111111111;
   49312: result <= 12'b111111111111;
   49313: result <= 12'b111111111111;
   49314: result <= 12'b111111111111;
   49315: result <= 12'b111111111111;
   49316: result <= 12'b111111111111;
   49317: result <= 12'b111111111111;
   49318: result <= 12'b111111111111;
   49319: result <= 12'b111111111111;
   49320: result <= 12'b111111111111;
   49321: result <= 12'b111111111111;
   49322: result <= 12'b111111111111;
   49323: result <= 12'b111111111111;
   49324: result <= 12'b111111111111;
   49325: result <= 12'b111111111111;
   49326: result <= 12'b111111111111;
   49327: result <= 12'b111111111111;
   49328: result <= 12'b111111111111;
   49329: result <= 12'b111111111111;
   49330: result <= 12'b111111111111;
   49331: result <= 12'b111111111111;
   49332: result <= 12'b111111111111;
   49333: result <= 12'b111111111111;
   49334: result <= 12'b111111111111;
   49335: result <= 12'b111111111111;
   49336: result <= 12'b111111111111;
   49337: result <= 12'b111111111111;
   49338: result <= 12'b111111111111;
   49339: result <= 12'b111111111111;
   49340: result <= 12'b111111111111;
   49341: result <= 12'b111111111111;
   49342: result <= 12'b111111111111;
   49343: result <= 12'b111111111111;
   49344: result <= 12'b111111111111;
   49345: result <= 12'b111111111111;
   49346: result <= 12'b111111111111;
   49347: result <= 12'b111111111111;
   49348: result <= 12'b111111111111;
   49349: result <= 12'b111111111111;
   49350: result <= 12'b111111111111;
   49351: result <= 12'b111111111111;
   49352: result <= 12'b111111111111;
   49353: result <= 12'b111111111111;
   49354: result <= 12'b111111111111;
   49355: result <= 12'b111111111111;
   49356: result <= 12'b111111111111;
   49357: result <= 12'b111111111111;
   49358: result <= 12'b111111111111;
   49359: result <= 12'b111111111111;
   49360: result <= 12'b111111111111;
   49361: result <= 12'b111111111111;
   49362: result <= 12'b111111111111;
   49363: result <= 12'b111111111111;
   49364: result <= 12'b111111111111;
   49365: result <= 12'b111111111111;
   49366: result <= 12'b111111111111;
   49367: result <= 12'b111111111111;
   49368: result <= 12'b111111111111;
   49369: result <= 12'b111111111111;
   49370: result <= 12'b111111111111;
   49371: result <= 12'b111111111111;
   49372: result <= 12'b111111111111;
   49373: result <= 12'b111111111111;
   49374: result <= 12'b111111111111;
   49375: result <= 12'b111111111111;
   49376: result <= 12'b111111111111;
   49377: result <= 12'b111111111111;
   49378: result <= 12'b111111111111;
   49379: result <= 12'b111111111111;
   49380: result <= 12'b111111111111;
   49381: result <= 12'b111111111111;
   49382: result <= 12'b111111111111;
   49383: result <= 12'b111111111111;
   49384: result <= 12'b111111111111;
   49385: result <= 12'b111111111111;
   49386: result <= 12'b111111111111;
   49387: result <= 12'b111111111111;
   49388: result <= 12'b111111111111;
   49389: result <= 12'b111111111111;
   49390: result <= 12'b111111111111;
   49391: result <= 12'b111111111111;
   49392: result <= 12'b111111111111;
   49393: result <= 12'b111111111111;
   49394: result <= 12'b111111111111;
   49395: result <= 12'b111111111111;
   49396: result <= 12'b111111111111;
   49397: result <= 12'b111111111111;
   49398: result <= 12'b111111111111;
   49399: result <= 12'b111111111111;
   49400: result <= 12'b111111111111;
   49401: result <= 12'b111111111111;
   49402: result <= 12'b111111111111;
   49403: result <= 12'b111111111111;
   49404: result <= 12'b111111111111;
   49405: result <= 12'b111111111111;
   49406: result <= 12'b111111111111;
   49407: result <= 12'b111111111111;
   49408: result <= 12'b111111111111;
   49409: result <= 12'b111111111111;
   49410: result <= 12'b111111111111;
   49411: result <= 12'b111111111111;
   49412: result <= 12'b111111111111;
   49413: result <= 12'b111111111111;
   49414: result <= 12'b111111111111;
   49415: result <= 12'b111111111111;
   49416: result <= 12'b111111111111;
   49417: result <= 12'b111111111111;
   49418: result <= 12'b111111111111;
   49419: result <= 12'b111111111111;
   49420: result <= 12'b111111111111;
   49421: result <= 12'b111111111111;
   49422: result <= 12'b111111111111;
   49423: result <= 12'b111111111111;
   49424: result <= 12'b111111111111;
   49425: result <= 12'b111111111111;
   49426: result <= 12'b111111111111;
   49427: result <= 12'b111111111111;
   49428: result <= 12'b111111111111;
   49429: result <= 12'b111111111111;
   49430: result <= 12'b111111111111;
   49431: result <= 12'b111111111111;
   49432: result <= 12'b111111111111;
   49433: result <= 12'b111111111111;
   49434: result <= 12'b111111111111;
   49435: result <= 12'b111111111111;
   49436: result <= 12'b111111111111;
   49437: result <= 12'b111111111111;
   49438: result <= 12'b111111111111;
   49439: result <= 12'b111111111111;
   49440: result <= 12'b111111111111;
   49441: result <= 12'b111111111111;
   49442: result <= 12'b111111111111;
   49443: result <= 12'b111111111111;
   49444: result <= 12'b111111111111;
   49445: result <= 12'b111111111111;
   49446: result <= 12'b111111111111;
   49447: result <= 12'b111111111111;
   49448: result <= 12'b111111111111;
   49449: result <= 12'b111111111111;
   49450: result <= 12'b111111111111;
   49451: result <= 12'b111111111111;
   49452: result <= 12'b111111111111;
   49453: result <= 12'b111111111111;
   49454: result <= 12'b111111111111;
   49455: result <= 12'b111111111111;
   49456: result <= 12'b111111111111;
   49457: result <= 12'b111111111111;
   49458: result <= 12'b111111111111;
   49459: result <= 12'b111111111111;
   49460: result <= 12'b111111111111;
   49461: result <= 12'b111111111111;
   49462: result <= 12'b111111111111;
   49463: result <= 12'b111111111111;
   49464: result <= 12'b111111111111;
   49465: result <= 12'b111111111111;
   49466: result <= 12'b111111111111;
   49467: result <= 12'b111111111111;
   49468: result <= 12'b111111111111;
   49469: result <= 12'b111111111111;
   49470: result <= 12'b111111111111;
   49471: result <= 12'b111111111111;
   49472: result <= 12'b111111111111;
   49473: result <= 12'b111111111111;
   49474: result <= 12'b111111111111;
   49475: result <= 12'b111111111111;
   49476: result <= 12'b111111111111;
   49477: result <= 12'b111111111111;
   49478: result <= 12'b111111111110;
   49479: result <= 12'b111111111110;
   49480: result <= 12'b111111111110;
   49481: result <= 12'b111111111110;
   49482: result <= 12'b111111111110;
   49483: result <= 12'b111111111110;
   49484: result <= 12'b111111111110;
   49485: result <= 12'b111111111110;
   49486: result <= 12'b111111111110;
   49487: result <= 12'b111111111110;
   49488: result <= 12'b111111111110;
   49489: result <= 12'b111111111110;
   49490: result <= 12'b111111111110;
   49491: result <= 12'b111111111110;
   49492: result <= 12'b111111111110;
   49493: result <= 12'b111111111110;
   49494: result <= 12'b111111111110;
   49495: result <= 12'b111111111110;
   49496: result <= 12'b111111111110;
   49497: result <= 12'b111111111110;
   49498: result <= 12'b111111111110;
   49499: result <= 12'b111111111110;
   49500: result <= 12'b111111111110;
   49501: result <= 12'b111111111110;
   49502: result <= 12'b111111111110;
   49503: result <= 12'b111111111110;
   49504: result <= 12'b111111111110;
   49505: result <= 12'b111111111110;
   49506: result <= 12'b111111111110;
   49507: result <= 12'b111111111110;
   49508: result <= 12'b111111111110;
   49509: result <= 12'b111111111110;
   49510: result <= 12'b111111111110;
   49511: result <= 12'b111111111110;
   49512: result <= 12'b111111111110;
   49513: result <= 12'b111111111110;
   49514: result <= 12'b111111111110;
   49515: result <= 12'b111111111110;
   49516: result <= 12'b111111111110;
   49517: result <= 12'b111111111110;
   49518: result <= 12'b111111111110;
   49519: result <= 12'b111111111110;
   49520: result <= 12'b111111111110;
   49521: result <= 12'b111111111110;
   49522: result <= 12'b111111111110;
   49523: result <= 12'b111111111110;
   49524: result <= 12'b111111111110;
   49525: result <= 12'b111111111110;
   49526: result <= 12'b111111111110;
   49527: result <= 12'b111111111110;
   49528: result <= 12'b111111111110;
   49529: result <= 12'b111111111110;
   49530: result <= 12'b111111111110;
   49531: result <= 12'b111111111110;
   49532: result <= 12'b111111111110;
   49533: result <= 12'b111111111110;
   49534: result <= 12'b111111111110;
   49535: result <= 12'b111111111110;
   49536: result <= 12'b111111111110;
   49537: result <= 12'b111111111110;
   49538: result <= 12'b111111111110;
   49539: result <= 12'b111111111110;
   49540: result <= 12'b111111111110;
   49541: result <= 12'b111111111110;
   49542: result <= 12'b111111111110;
   49543: result <= 12'b111111111110;
   49544: result <= 12'b111111111110;
   49545: result <= 12'b111111111110;
   49546: result <= 12'b111111111110;
   49547: result <= 12'b111111111110;
   49548: result <= 12'b111111111110;
   49549: result <= 12'b111111111110;
   49550: result <= 12'b111111111110;
   49551: result <= 12'b111111111110;
   49552: result <= 12'b111111111110;
   49553: result <= 12'b111111111110;
   49554: result <= 12'b111111111110;
   49555: result <= 12'b111111111110;
   49556: result <= 12'b111111111110;
   49557: result <= 12'b111111111110;
   49558: result <= 12'b111111111110;
   49559: result <= 12'b111111111110;
   49560: result <= 12'b111111111110;
   49561: result <= 12'b111111111110;
   49562: result <= 12'b111111111110;
   49563: result <= 12'b111111111110;
   49564: result <= 12'b111111111110;
   49565: result <= 12'b111111111110;
   49566: result <= 12'b111111111110;
   49567: result <= 12'b111111111110;
   49568: result <= 12'b111111111110;
   49569: result <= 12'b111111111110;
   49570: result <= 12'b111111111110;
   49571: result <= 12'b111111111110;
   49572: result <= 12'b111111111110;
   49573: result <= 12'b111111111110;
   49574: result <= 12'b111111111110;
   49575: result <= 12'b111111111110;
   49576: result <= 12'b111111111110;
   49577: result <= 12'b111111111110;
   49578: result <= 12'b111111111110;
   49579: result <= 12'b111111111110;
   49580: result <= 12'b111111111110;
   49581: result <= 12'b111111111110;
   49582: result <= 12'b111111111110;
   49583: result <= 12'b111111111110;
   49584: result <= 12'b111111111110;
   49585: result <= 12'b111111111110;
   49586: result <= 12'b111111111110;
   49587: result <= 12'b111111111110;
   49588: result <= 12'b111111111110;
   49589: result <= 12'b111111111110;
   49590: result <= 12'b111111111110;
   49591: result <= 12'b111111111110;
   49592: result <= 12'b111111111110;
   49593: result <= 12'b111111111110;
   49594: result <= 12'b111111111110;
   49595: result <= 12'b111111111110;
   49596: result <= 12'b111111111110;
   49597: result <= 12'b111111111110;
   49598: result <= 12'b111111111110;
   49599: result <= 12'b111111111110;
   49600: result <= 12'b111111111110;
   49601: result <= 12'b111111111110;
   49602: result <= 12'b111111111110;
   49603: result <= 12'b111111111110;
   49604: result <= 12'b111111111110;
   49605: result <= 12'b111111111110;
   49606: result <= 12'b111111111110;
   49607: result <= 12'b111111111110;
   49608: result <= 12'b111111111110;
   49609: result <= 12'b111111111110;
   49610: result <= 12'b111111111110;
   49611: result <= 12'b111111111110;
   49612: result <= 12'b111111111110;
   49613: result <= 12'b111111111101;
   49614: result <= 12'b111111111101;
   49615: result <= 12'b111111111101;
   49616: result <= 12'b111111111101;
   49617: result <= 12'b111111111101;
   49618: result <= 12'b111111111101;
   49619: result <= 12'b111111111101;
   49620: result <= 12'b111111111101;
   49621: result <= 12'b111111111101;
   49622: result <= 12'b111111111101;
   49623: result <= 12'b111111111101;
   49624: result <= 12'b111111111101;
   49625: result <= 12'b111111111101;
   49626: result <= 12'b111111111101;
   49627: result <= 12'b111111111101;
   49628: result <= 12'b111111111101;
   49629: result <= 12'b111111111101;
   49630: result <= 12'b111111111101;
   49631: result <= 12'b111111111101;
   49632: result <= 12'b111111111101;
   49633: result <= 12'b111111111101;
   49634: result <= 12'b111111111101;
   49635: result <= 12'b111111111101;
   49636: result <= 12'b111111111101;
   49637: result <= 12'b111111111101;
   49638: result <= 12'b111111111101;
   49639: result <= 12'b111111111101;
   49640: result <= 12'b111111111101;
   49641: result <= 12'b111111111101;
   49642: result <= 12'b111111111101;
   49643: result <= 12'b111111111101;
   49644: result <= 12'b111111111101;
   49645: result <= 12'b111111111101;
   49646: result <= 12'b111111111101;
   49647: result <= 12'b111111111101;
   49648: result <= 12'b111111111101;
   49649: result <= 12'b111111111101;
   49650: result <= 12'b111111111101;
   49651: result <= 12'b111111111101;
   49652: result <= 12'b111111111101;
   49653: result <= 12'b111111111101;
   49654: result <= 12'b111111111101;
   49655: result <= 12'b111111111101;
   49656: result <= 12'b111111111101;
   49657: result <= 12'b111111111101;
   49658: result <= 12'b111111111101;
   49659: result <= 12'b111111111101;
   49660: result <= 12'b111111111101;
   49661: result <= 12'b111111111101;
   49662: result <= 12'b111111111101;
   49663: result <= 12'b111111111101;
   49664: result <= 12'b111111111101;
   49665: result <= 12'b111111111101;
   49666: result <= 12'b111111111101;
   49667: result <= 12'b111111111101;
   49668: result <= 12'b111111111101;
   49669: result <= 12'b111111111101;
   49670: result <= 12'b111111111101;
   49671: result <= 12'b111111111101;
   49672: result <= 12'b111111111101;
   49673: result <= 12'b111111111101;
   49674: result <= 12'b111111111101;
   49675: result <= 12'b111111111101;
   49676: result <= 12'b111111111101;
   49677: result <= 12'b111111111101;
   49678: result <= 12'b111111111101;
   49679: result <= 12'b111111111101;
   49680: result <= 12'b111111111101;
   49681: result <= 12'b111111111101;
   49682: result <= 12'b111111111101;
   49683: result <= 12'b111111111101;
   49684: result <= 12'b111111111101;
   49685: result <= 12'b111111111101;
   49686: result <= 12'b111111111101;
   49687: result <= 12'b111111111101;
   49688: result <= 12'b111111111101;
   49689: result <= 12'b111111111101;
   49690: result <= 12'b111111111101;
   49691: result <= 12'b111111111101;
   49692: result <= 12'b111111111101;
   49693: result <= 12'b111111111101;
   49694: result <= 12'b111111111101;
   49695: result <= 12'b111111111101;
   49696: result <= 12'b111111111101;
   49697: result <= 12'b111111111101;
   49698: result <= 12'b111111111101;
   49699: result <= 12'b111111111101;
   49700: result <= 12'b111111111101;
   49701: result <= 12'b111111111101;
   49702: result <= 12'b111111111101;
   49703: result <= 12'b111111111101;
   49704: result <= 12'b111111111101;
   49705: result <= 12'b111111111101;
   49706: result <= 12'b111111111101;
   49707: result <= 12'b111111111101;
   49708: result <= 12'b111111111101;
   49709: result <= 12'b111111111101;
   49710: result <= 12'b111111111101;
   49711: result <= 12'b111111111101;
   49712: result <= 12'b111111111101;
   49713: result <= 12'b111111111101;
   49714: result <= 12'b111111111101;
   49715: result <= 12'b111111111101;
   49716: result <= 12'b111111111101;
   49717: result <= 12'b111111111100;
   49718: result <= 12'b111111111100;
   49719: result <= 12'b111111111100;
   49720: result <= 12'b111111111100;
   49721: result <= 12'b111111111100;
   49722: result <= 12'b111111111100;
   49723: result <= 12'b111111111100;
   49724: result <= 12'b111111111100;
   49725: result <= 12'b111111111100;
   49726: result <= 12'b111111111100;
   49727: result <= 12'b111111111100;
   49728: result <= 12'b111111111100;
   49729: result <= 12'b111111111100;
   49730: result <= 12'b111111111100;
   49731: result <= 12'b111111111100;
   49732: result <= 12'b111111111100;
   49733: result <= 12'b111111111100;
   49734: result <= 12'b111111111100;
   49735: result <= 12'b111111111100;
   49736: result <= 12'b111111111100;
   49737: result <= 12'b111111111100;
   49738: result <= 12'b111111111100;
   49739: result <= 12'b111111111100;
   49740: result <= 12'b111111111100;
   49741: result <= 12'b111111111100;
   49742: result <= 12'b111111111100;
   49743: result <= 12'b111111111100;
   49744: result <= 12'b111111111100;
   49745: result <= 12'b111111111100;
   49746: result <= 12'b111111111100;
   49747: result <= 12'b111111111100;
   49748: result <= 12'b111111111100;
   49749: result <= 12'b111111111100;
   49750: result <= 12'b111111111100;
   49751: result <= 12'b111111111100;
   49752: result <= 12'b111111111100;
   49753: result <= 12'b111111111100;
   49754: result <= 12'b111111111100;
   49755: result <= 12'b111111111100;
   49756: result <= 12'b111111111100;
   49757: result <= 12'b111111111100;
   49758: result <= 12'b111111111100;
   49759: result <= 12'b111111111100;
   49760: result <= 12'b111111111100;
   49761: result <= 12'b111111111100;
   49762: result <= 12'b111111111100;
   49763: result <= 12'b111111111100;
   49764: result <= 12'b111111111100;
   49765: result <= 12'b111111111100;
   49766: result <= 12'b111111111100;
   49767: result <= 12'b111111111100;
   49768: result <= 12'b111111111100;
   49769: result <= 12'b111111111100;
   49770: result <= 12'b111111111100;
   49771: result <= 12'b111111111100;
   49772: result <= 12'b111111111100;
   49773: result <= 12'b111111111100;
   49774: result <= 12'b111111111100;
   49775: result <= 12'b111111111100;
   49776: result <= 12'b111111111100;
   49777: result <= 12'b111111111100;
   49778: result <= 12'b111111111100;
   49779: result <= 12'b111111111100;
   49780: result <= 12'b111111111100;
   49781: result <= 12'b111111111100;
   49782: result <= 12'b111111111100;
   49783: result <= 12'b111111111100;
   49784: result <= 12'b111111111100;
   49785: result <= 12'b111111111100;
   49786: result <= 12'b111111111100;
   49787: result <= 12'b111111111100;
   49788: result <= 12'b111111111100;
   49789: result <= 12'b111111111100;
   49790: result <= 12'b111111111100;
   49791: result <= 12'b111111111100;
   49792: result <= 12'b111111111100;
   49793: result <= 12'b111111111100;
   49794: result <= 12'b111111111100;
   49795: result <= 12'b111111111100;
   49796: result <= 12'b111111111100;
   49797: result <= 12'b111111111100;
   49798: result <= 12'b111111111100;
   49799: result <= 12'b111111111100;
   49800: result <= 12'b111111111100;
   49801: result <= 12'b111111111100;
   49802: result <= 12'b111111111100;
   49803: result <= 12'b111111111100;
   49804: result <= 12'b111111111100;
   49805: result <= 12'b111111111011;
   49806: result <= 12'b111111111011;
   49807: result <= 12'b111111111011;
   49808: result <= 12'b111111111011;
   49809: result <= 12'b111111111011;
   49810: result <= 12'b111111111011;
   49811: result <= 12'b111111111011;
   49812: result <= 12'b111111111011;
   49813: result <= 12'b111111111011;
   49814: result <= 12'b111111111011;
   49815: result <= 12'b111111111011;
   49816: result <= 12'b111111111011;
   49817: result <= 12'b111111111011;
   49818: result <= 12'b111111111011;
   49819: result <= 12'b111111111011;
   49820: result <= 12'b111111111011;
   49821: result <= 12'b111111111011;
   49822: result <= 12'b111111111011;
   49823: result <= 12'b111111111011;
   49824: result <= 12'b111111111011;
   49825: result <= 12'b111111111011;
   49826: result <= 12'b111111111011;
   49827: result <= 12'b111111111011;
   49828: result <= 12'b111111111011;
   49829: result <= 12'b111111111011;
   49830: result <= 12'b111111111011;
   49831: result <= 12'b111111111011;
   49832: result <= 12'b111111111011;
   49833: result <= 12'b111111111011;
   49834: result <= 12'b111111111011;
   49835: result <= 12'b111111111011;
   49836: result <= 12'b111111111011;
   49837: result <= 12'b111111111011;
   49838: result <= 12'b111111111011;
   49839: result <= 12'b111111111011;
   49840: result <= 12'b111111111011;
   49841: result <= 12'b111111111011;
   49842: result <= 12'b111111111011;
   49843: result <= 12'b111111111011;
   49844: result <= 12'b111111111011;
   49845: result <= 12'b111111111011;
   49846: result <= 12'b111111111011;
   49847: result <= 12'b111111111011;
   49848: result <= 12'b111111111011;
   49849: result <= 12'b111111111011;
   49850: result <= 12'b111111111011;
   49851: result <= 12'b111111111011;
   49852: result <= 12'b111111111011;
   49853: result <= 12'b111111111011;
   49854: result <= 12'b111111111011;
   49855: result <= 12'b111111111011;
   49856: result <= 12'b111111111011;
   49857: result <= 12'b111111111011;
   49858: result <= 12'b111111111011;
   49859: result <= 12'b111111111011;
   49860: result <= 12'b111111111011;
   49861: result <= 12'b111111111011;
   49862: result <= 12'b111111111011;
   49863: result <= 12'b111111111011;
   49864: result <= 12'b111111111011;
   49865: result <= 12'b111111111011;
   49866: result <= 12'b111111111011;
   49867: result <= 12'b111111111011;
   49868: result <= 12'b111111111011;
   49869: result <= 12'b111111111011;
   49870: result <= 12'b111111111011;
   49871: result <= 12'b111111111011;
   49872: result <= 12'b111111111011;
   49873: result <= 12'b111111111011;
   49874: result <= 12'b111111111011;
   49875: result <= 12'b111111111011;
   49876: result <= 12'b111111111011;
   49877: result <= 12'b111111111011;
   49878: result <= 12'b111111111011;
   49879: result <= 12'b111111111011;
   49880: result <= 12'b111111111011;
   49881: result <= 12'b111111111010;
   49882: result <= 12'b111111111010;
   49883: result <= 12'b111111111010;
   49884: result <= 12'b111111111010;
   49885: result <= 12'b111111111010;
   49886: result <= 12'b111111111010;
   49887: result <= 12'b111111111010;
   49888: result <= 12'b111111111010;
   49889: result <= 12'b111111111010;
   49890: result <= 12'b111111111010;
   49891: result <= 12'b111111111010;
   49892: result <= 12'b111111111010;
   49893: result <= 12'b111111111010;
   49894: result <= 12'b111111111010;
   49895: result <= 12'b111111111010;
   49896: result <= 12'b111111111010;
   49897: result <= 12'b111111111010;
   49898: result <= 12'b111111111010;
   49899: result <= 12'b111111111010;
   49900: result <= 12'b111111111010;
   49901: result <= 12'b111111111010;
   49902: result <= 12'b111111111010;
   49903: result <= 12'b111111111010;
   49904: result <= 12'b111111111010;
   49905: result <= 12'b111111111010;
   49906: result <= 12'b111111111010;
   49907: result <= 12'b111111111010;
   49908: result <= 12'b111111111010;
   49909: result <= 12'b111111111010;
   49910: result <= 12'b111111111010;
   49911: result <= 12'b111111111010;
   49912: result <= 12'b111111111010;
   49913: result <= 12'b111111111010;
   49914: result <= 12'b111111111010;
   49915: result <= 12'b111111111010;
   49916: result <= 12'b111111111010;
   49917: result <= 12'b111111111010;
   49918: result <= 12'b111111111010;
   49919: result <= 12'b111111111010;
   49920: result <= 12'b111111111010;
   49921: result <= 12'b111111111010;
   49922: result <= 12'b111111111010;
   49923: result <= 12'b111111111010;
   49924: result <= 12'b111111111010;
   49925: result <= 12'b111111111010;
   49926: result <= 12'b111111111010;
   49927: result <= 12'b111111111010;
   49928: result <= 12'b111111111010;
   49929: result <= 12'b111111111010;
   49930: result <= 12'b111111111010;
   49931: result <= 12'b111111111010;
   49932: result <= 12'b111111111010;
   49933: result <= 12'b111111111010;
   49934: result <= 12'b111111111010;
   49935: result <= 12'b111111111010;
   49936: result <= 12'b111111111010;
   49937: result <= 12'b111111111010;
   49938: result <= 12'b111111111010;
   49939: result <= 12'b111111111010;
   49940: result <= 12'b111111111010;
   49941: result <= 12'b111111111010;
   49942: result <= 12'b111111111010;
   49943: result <= 12'b111111111010;
   49944: result <= 12'b111111111010;
   49945: result <= 12'b111111111010;
   49946: result <= 12'b111111111010;
   49947: result <= 12'b111111111010;
   49948: result <= 12'b111111111010;
   49949: result <= 12'b111111111010;
   49950: result <= 12'b111111111010;
   49951: result <= 12'b111111111001;
   49952: result <= 12'b111111111001;
   49953: result <= 12'b111111111001;
   49954: result <= 12'b111111111001;
   49955: result <= 12'b111111111001;
   49956: result <= 12'b111111111001;
   49957: result <= 12'b111111111001;
   49958: result <= 12'b111111111001;
   49959: result <= 12'b111111111001;
   49960: result <= 12'b111111111001;
   49961: result <= 12'b111111111001;
   49962: result <= 12'b111111111001;
   49963: result <= 12'b111111111001;
   49964: result <= 12'b111111111001;
   49965: result <= 12'b111111111001;
   49966: result <= 12'b111111111001;
   49967: result <= 12'b111111111001;
   49968: result <= 12'b111111111001;
   49969: result <= 12'b111111111001;
   49970: result <= 12'b111111111001;
   49971: result <= 12'b111111111001;
   49972: result <= 12'b111111111001;
   49973: result <= 12'b111111111001;
   49974: result <= 12'b111111111001;
   49975: result <= 12'b111111111001;
   49976: result <= 12'b111111111001;
   49977: result <= 12'b111111111001;
   49978: result <= 12'b111111111001;
   49979: result <= 12'b111111111001;
   49980: result <= 12'b111111111001;
   49981: result <= 12'b111111111001;
   49982: result <= 12'b111111111001;
   49983: result <= 12'b111111111001;
   49984: result <= 12'b111111111001;
   49985: result <= 12'b111111111001;
   49986: result <= 12'b111111111001;
   49987: result <= 12'b111111111001;
   49988: result <= 12'b111111111001;
   49989: result <= 12'b111111111001;
   49990: result <= 12'b111111111001;
   49991: result <= 12'b111111111001;
   49992: result <= 12'b111111111001;
   49993: result <= 12'b111111111001;
   49994: result <= 12'b111111111001;
   49995: result <= 12'b111111111001;
   49996: result <= 12'b111111111001;
   49997: result <= 12'b111111111001;
   49998: result <= 12'b111111111001;
   49999: result <= 12'b111111111001;
   50000: result <= 12'b111111111001;
   50001: result <= 12'b111111111001;
   50002: result <= 12'b111111111001;
   50003: result <= 12'b111111111001;
   50004: result <= 12'b111111111001;
   50005: result <= 12'b111111111001;
   50006: result <= 12'b111111111001;
   50007: result <= 12'b111111111001;
   50008: result <= 12'b111111111001;
   50009: result <= 12'b111111111001;
   50010: result <= 12'b111111111001;
   50011: result <= 12'b111111111001;
   50012: result <= 12'b111111111001;
   50013: result <= 12'b111111111001;
   50014: result <= 12'b111111111001;
   50015: result <= 12'b111111111000;
   50016: result <= 12'b111111111000;
   50017: result <= 12'b111111111000;
   50018: result <= 12'b111111111000;
   50019: result <= 12'b111111111000;
   50020: result <= 12'b111111111000;
   50021: result <= 12'b111111111000;
   50022: result <= 12'b111111111000;
   50023: result <= 12'b111111111000;
   50024: result <= 12'b111111111000;
   50025: result <= 12'b111111111000;
   50026: result <= 12'b111111111000;
   50027: result <= 12'b111111111000;
   50028: result <= 12'b111111111000;
   50029: result <= 12'b111111111000;
   50030: result <= 12'b111111111000;
   50031: result <= 12'b111111111000;
   50032: result <= 12'b111111111000;
   50033: result <= 12'b111111111000;
   50034: result <= 12'b111111111000;
   50035: result <= 12'b111111111000;
   50036: result <= 12'b111111111000;
   50037: result <= 12'b111111111000;
   50038: result <= 12'b111111111000;
   50039: result <= 12'b111111111000;
   50040: result <= 12'b111111111000;
   50041: result <= 12'b111111111000;
   50042: result <= 12'b111111111000;
   50043: result <= 12'b111111111000;
   50044: result <= 12'b111111111000;
   50045: result <= 12'b111111111000;
   50046: result <= 12'b111111111000;
   50047: result <= 12'b111111111000;
   50048: result <= 12'b111111111000;
   50049: result <= 12'b111111111000;
   50050: result <= 12'b111111111000;
   50051: result <= 12'b111111111000;
   50052: result <= 12'b111111111000;
   50053: result <= 12'b111111111000;
   50054: result <= 12'b111111111000;
   50055: result <= 12'b111111111000;
   50056: result <= 12'b111111111000;
   50057: result <= 12'b111111111000;
   50058: result <= 12'b111111111000;
   50059: result <= 12'b111111111000;
   50060: result <= 12'b111111111000;
   50061: result <= 12'b111111111000;
   50062: result <= 12'b111111111000;
   50063: result <= 12'b111111111000;
   50064: result <= 12'b111111111000;
   50065: result <= 12'b111111111000;
   50066: result <= 12'b111111111000;
   50067: result <= 12'b111111111000;
   50068: result <= 12'b111111111000;
   50069: result <= 12'b111111111000;
   50070: result <= 12'b111111111000;
   50071: result <= 12'b111111111000;
   50072: result <= 12'b111111111000;
   50073: result <= 12'b111111111000;
   50074: result <= 12'b111111111000;
   50075: result <= 12'b111111110111;
   50076: result <= 12'b111111110111;
   50077: result <= 12'b111111110111;
   50078: result <= 12'b111111110111;
   50079: result <= 12'b111111110111;
   50080: result <= 12'b111111110111;
   50081: result <= 12'b111111110111;
   50082: result <= 12'b111111110111;
   50083: result <= 12'b111111110111;
   50084: result <= 12'b111111110111;
   50085: result <= 12'b111111110111;
   50086: result <= 12'b111111110111;
   50087: result <= 12'b111111110111;
   50088: result <= 12'b111111110111;
   50089: result <= 12'b111111110111;
   50090: result <= 12'b111111110111;
   50091: result <= 12'b111111110111;
   50092: result <= 12'b111111110111;
   50093: result <= 12'b111111110111;
   50094: result <= 12'b111111110111;
   50095: result <= 12'b111111110111;
   50096: result <= 12'b111111110111;
   50097: result <= 12'b111111110111;
   50098: result <= 12'b111111110111;
   50099: result <= 12'b111111110111;
   50100: result <= 12'b111111110111;
   50101: result <= 12'b111111110111;
   50102: result <= 12'b111111110111;
   50103: result <= 12'b111111110111;
   50104: result <= 12'b111111110111;
   50105: result <= 12'b111111110111;
   50106: result <= 12'b111111110111;
   50107: result <= 12'b111111110111;
   50108: result <= 12'b111111110111;
   50109: result <= 12'b111111110111;
   50110: result <= 12'b111111110111;
   50111: result <= 12'b111111110111;
   50112: result <= 12'b111111110111;
   50113: result <= 12'b111111110111;
   50114: result <= 12'b111111110111;
   50115: result <= 12'b111111110111;
   50116: result <= 12'b111111110111;
   50117: result <= 12'b111111110111;
   50118: result <= 12'b111111110111;
   50119: result <= 12'b111111110111;
   50120: result <= 12'b111111110111;
   50121: result <= 12'b111111110111;
   50122: result <= 12'b111111110111;
   50123: result <= 12'b111111110111;
   50124: result <= 12'b111111110111;
   50125: result <= 12'b111111110111;
   50126: result <= 12'b111111110111;
   50127: result <= 12'b111111110111;
   50128: result <= 12'b111111110111;
   50129: result <= 12'b111111110111;
   50130: result <= 12'b111111110111;
   50131: result <= 12'b111111110110;
   50132: result <= 12'b111111110110;
   50133: result <= 12'b111111110110;
   50134: result <= 12'b111111110110;
   50135: result <= 12'b111111110110;
   50136: result <= 12'b111111110110;
   50137: result <= 12'b111111110110;
   50138: result <= 12'b111111110110;
   50139: result <= 12'b111111110110;
   50140: result <= 12'b111111110110;
   50141: result <= 12'b111111110110;
   50142: result <= 12'b111111110110;
   50143: result <= 12'b111111110110;
   50144: result <= 12'b111111110110;
   50145: result <= 12'b111111110110;
   50146: result <= 12'b111111110110;
   50147: result <= 12'b111111110110;
   50148: result <= 12'b111111110110;
   50149: result <= 12'b111111110110;
   50150: result <= 12'b111111110110;
   50151: result <= 12'b111111110110;
   50152: result <= 12'b111111110110;
   50153: result <= 12'b111111110110;
   50154: result <= 12'b111111110110;
   50155: result <= 12'b111111110110;
   50156: result <= 12'b111111110110;
   50157: result <= 12'b111111110110;
   50158: result <= 12'b111111110110;
   50159: result <= 12'b111111110110;
   50160: result <= 12'b111111110110;
   50161: result <= 12'b111111110110;
   50162: result <= 12'b111111110110;
   50163: result <= 12'b111111110110;
   50164: result <= 12'b111111110110;
   50165: result <= 12'b111111110110;
   50166: result <= 12'b111111110110;
   50167: result <= 12'b111111110110;
   50168: result <= 12'b111111110110;
   50169: result <= 12'b111111110110;
   50170: result <= 12'b111111110110;
   50171: result <= 12'b111111110110;
   50172: result <= 12'b111111110110;
   50173: result <= 12'b111111110110;
   50174: result <= 12'b111111110110;
   50175: result <= 12'b111111110110;
   50176: result <= 12'b111111110110;
   50177: result <= 12'b111111110110;
   50178: result <= 12'b111111110110;
   50179: result <= 12'b111111110110;
   50180: result <= 12'b111111110110;
   50181: result <= 12'b111111110110;
   50182: result <= 12'b111111110110;
   50183: result <= 12'b111111110110;
   50184: result <= 12'b111111110101;
   50185: result <= 12'b111111110101;
   50186: result <= 12'b111111110101;
   50187: result <= 12'b111111110101;
   50188: result <= 12'b111111110101;
   50189: result <= 12'b111111110101;
   50190: result <= 12'b111111110101;
   50191: result <= 12'b111111110101;
   50192: result <= 12'b111111110101;
   50193: result <= 12'b111111110101;
   50194: result <= 12'b111111110101;
   50195: result <= 12'b111111110101;
   50196: result <= 12'b111111110101;
   50197: result <= 12'b111111110101;
   50198: result <= 12'b111111110101;
   50199: result <= 12'b111111110101;
   50200: result <= 12'b111111110101;
   50201: result <= 12'b111111110101;
   50202: result <= 12'b111111110101;
   50203: result <= 12'b111111110101;
   50204: result <= 12'b111111110101;
   50205: result <= 12'b111111110101;
   50206: result <= 12'b111111110101;
   50207: result <= 12'b111111110101;
   50208: result <= 12'b111111110101;
   50209: result <= 12'b111111110101;
   50210: result <= 12'b111111110101;
   50211: result <= 12'b111111110101;
   50212: result <= 12'b111111110101;
   50213: result <= 12'b111111110101;
   50214: result <= 12'b111111110101;
   50215: result <= 12'b111111110101;
   50216: result <= 12'b111111110101;
   50217: result <= 12'b111111110101;
   50218: result <= 12'b111111110101;
   50219: result <= 12'b111111110101;
   50220: result <= 12'b111111110101;
   50221: result <= 12'b111111110101;
   50222: result <= 12'b111111110101;
   50223: result <= 12'b111111110101;
   50224: result <= 12'b111111110101;
   50225: result <= 12'b111111110101;
   50226: result <= 12'b111111110101;
   50227: result <= 12'b111111110101;
   50228: result <= 12'b111111110101;
   50229: result <= 12'b111111110101;
   50230: result <= 12'b111111110101;
   50231: result <= 12'b111111110101;
   50232: result <= 12'b111111110101;
   50233: result <= 12'b111111110101;
   50234: result <= 12'b111111110100;
   50235: result <= 12'b111111110100;
   50236: result <= 12'b111111110100;
   50237: result <= 12'b111111110100;
   50238: result <= 12'b111111110100;
   50239: result <= 12'b111111110100;
   50240: result <= 12'b111111110100;
   50241: result <= 12'b111111110100;
   50242: result <= 12'b111111110100;
   50243: result <= 12'b111111110100;
   50244: result <= 12'b111111110100;
   50245: result <= 12'b111111110100;
   50246: result <= 12'b111111110100;
   50247: result <= 12'b111111110100;
   50248: result <= 12'b111111110100;
   50249: result <= 12'b111111110100;
   50250: result <= 12'b111111110100;
   50251: result <= 12'b111111110100;
   50252: result <= 12'b111111110100;
   50253: result <= 12'b111111110100;
   50254: result <= 12'b111111110100;
   50255: result <= 12'b111111110100;
   50256: result <= 12'b111111110100;
   50257: result <= 12'b111111110100;
   50258: result <= 12'b111111110100;
   50259: result <= 12'b111111110100;
   50260: result <= 12'b111111110100;
   50261: result <= 12'b111111110100;
   50262: result <= 12'b111111110100;
   50263: result <= 12'b111111110100;
   50264: result <= 12'b111111110100;
   50265: result <= 12'b111111110100;
   50266: result <= 12'b111111110100;
   50267: result <= 12'b111111110100;
   50268: result <= 12'b111111110100;
   50269: result <= 12'b111111110100;
   50270: result <= 12'b111111110100;
   50271: result <= 12'b111111110100;
   50272: result <= 12'b111111110100;
   50273: result <= 12'b111111110100;
   50274: result <= 12'b111111110100;
   50275: result <= 12'b111111110100;
   50276: result <= 12'b111111110100;
   50277: result <= 12'b111111110100;
   50278: result <= 12'b111111110100;
   50279: result <= 12'b111111110100;
   50280: result <= 12'b111111110100;
   50281: result <= 12'b111111110100;
   50282: result <= 12'b111111110011;
   50283: result <= 12'b111111110011;
   50284: result <= 12'b111111110011;
   50285: result <= 12'b111111110011;
   50286: result <= 12'b111111110011;
   50287: result <= 12'b111111110011;
   50288: result <= 12'b111111110011;
   50289: result <= 12'b111111110011;
   50290: result <= 12'b111111110011;
   50291: result <= 12'b111111110011;
   50292: result <= 12'b111111110011;
   50293: result <= 12'b111111110011;
   50294: result <= 12'b111111110011;
   50295: result <= 12'b111111110011;
   50296: result <= 12'b111111110011;
   50297: result <= 12'b111111110011;
   50298: result <= 12'b111111110011;
   50299: result <= 12'b111111110011;
   50300: result <= 12'b111111110011;
   50301: result <= 12'b111111110011;
   50302: result <= 12'b111111110011;
   50303: result <= 12'b111111110011;
   50304: result <= 12'b111111110011;
   50305: result <= 12'b111111110011;
   50306: result <= 12'b111111110011;
   50307: result <= 12'b111111110011;
   50308: result <= 12'b111111110011;
   50309: result <= 12'b111111110011;
   50310: result <= 12'b111111110011;
   50311: result <= 12'b111111110011;
   50312: result <= 12'b111111110011;
   50313: result <= 12'b111111110011;
   50314: result <= 12'b111111110011;
   50315: result <= 12'b111111110011;
   50316: result <= 12'b111111110011;
   50317: result <= 12'b111111110011;
   50318: result <= 12'b111111110011;
   50319: result <= 12'b111111110011;
   50320: result <= 12'b111111110011;
   50321: result <= 12'b111111110011;
   50322: result <= 12'b111111110011;
   50323: result <= 12'b111111110011;
   50324: result <= 12'b111111110011;
   50325: result <= 12'b111111110011;
   50326: result <= 12'b111111110011;
   50327: result <= 12'b111111110011;
   50328: result <= 12'b111111110010;
   50329: result <= 12'b111111110010;
   50330: result <= 12'b111111110010;
   50331: result <= 12'b111111110010;
   50332: result <= 12'b111111110010;
   50333: result <= 12'b111111110010;
   50334: result <= 12'b111111110010;
   50335: result <= 12'b111111110010;
   50336: result <= 12'b111111110010;
   50337: result <= 12'b111111110010;
   50338: result <= 12'b111111110010;
   50339: result <= 12'b111111110010;
   50340: result <= 12'b111111110010;
   50341: result <= 12'b111111110010;
   50342: result <= 12'b111111110010;
   50343: result <= 12'b111111110010;
   50344: result <= 12'b111111110010;
   50345: result <= 12'b111111110010;
   50346: result <= 12'b111111110010;
   50347: result <= 12'b111111110010;
   50348: result <= 12'b111111110010;
   50349: result <= 12'b111111110010;
   50350: result <= 12'b111111110010;
   50351: result <= 12'b111111110010;
   50352: result <= 12'b111111110010;
   50353: result <= 12'b111111110010;
   50354: result <= 12'b111111110010;
   50355: result <= 12'b111111110010;
   50356: result <= 12'b111111110010;
   50357: result <= 12'b111111110010;
   50358: result <= 12'b111111110010;
   50359: result <= 12'b111111110010;
   50360: result <= 12'b111111110010;
   50361: result <= 12'b111111110010;
   50362: result <= 12'b111111110010;
   50363: result <= 12'b111111110010;
   50364: result <= 12'b111111110010;
   50365: result <= 12'b111111110010;
   50366: result <= 12'b111111110010;
   50367: result <= 12'b111111110010;
   50368: result <= 12'b111111110010;
   50369: result <= 12'b111111110010;
   50370: result <= 12'b111111110010;
   50371: result <= 12'b111111110010;
   50372: result <= 12'b111111110010;
   50373: result <= 12'b111111110001;
   50374: result <= 12'b111111110001;
   50375: result <= 12'b111111110001;
   50376: result <= 12'b111111110001;
   50377: result <= 12'b111111110001;
   50378: result <= 12'b111111110001;
   50379: result <= 12'b111111110001;
   50380: result <= 12'b111111110001;
   50381: result <= 12'b111111110001;
   50382: result <= 12'b111111110001;
   50383: result <= 12'b111111110001;
   50384: result <= 12'b111111110001;
   50385: result <= 12'b111111110001;
   50386: result <= 12'b111111110001;
   50387: result <= 12'b111111110001;
   50388: result <= 12'b111111110001;
   50389: result <= 12'b111111110001;
   50390: result <= 12'b111111110001;
   50391: result <= 12'b111111110001;
   50392: result <= 12'b111111110001;
   50393: result <= 12'b111111110001;
   50394: result <= 12'b111111110001;
   50395: result <= 12'b111111110001;
   50396: result <= 12'b111111110001;
   50397: result <= 12'b111111110001;
   50398: result <= 12'b111111110001;
   50399: result <= 12'b111111110001;
   50400: result <= 12'b111111110001;
   50401: result <= 12'b111111110001;
   50402: result <= 12'b111111110001;
   50403: result <= 12'b111111110001;
   50404: result <= 12'b111111110001;
   50405: result <= 12'b111111110001;
   50406: result <= 12'b111111110001;
   50407: result <= 12'b111111110001;
   50408: result <= 12'b111111110001;
   50409: result <= 12'b111111110001;
   50410: result <= 12'b111111110001;
   50411: result <= 12'b111111110001;
   50412: result <= 12'b111111110001;
   50413: result <= 12'b111111110001;
   50414: result <= 12'b111111110001;
   50415: result <= 12'b111111110001;
   50416: result <= 12'b111111110000;
   50417: result <= 12'b111111110000;
   50418: result <= 12'b111111110000;
   50419: result <= 12'b111111110000;
   50420: result <= 12'b111111110000;
   50421: result <= 12'b111111110000;
   50422: result <= 12'b111111110000;
   50423: result <= 12'b111111110000;
   50424: result <= 12'b111111110000;
   50425: result <= 12'b111111110000;
   50426: result <= 12'b111111110000;
   50427: result <= 12'b111111110000;
   50428: result <= 12'b111111110000;
   50429: result <= 12'b111111110000;
   50430: result <= 12'b111111110000;
   50431: result <= 12'b111111110000;
   50432: result <= 12'b111111110000;
   50433: result <= 12'b111111110000;
   50434: result <= 12'b111111110000;
   50435: result <= 12'b111111110000;
   50436: result <= 12'b111111110000;
   50437: result <= 12'b111111110000;
   50438: result <= 12'b111111110000;
   50439: result <= 12'b111111110000;
   50440: result <= 12'b111111110000;
   50441: result <= 12'b111111110000;
   50442: result <= 12'b111111110000;
   50443: result <= 12'b111111110000;
   50444: result <= 12'b111111110000;
   50445: result <= 12'b111111110000;
   50446: result <= 12'b111111110000;
   50447: result <= 12'b111111110000;
   50448: result <= 12'b111111110000;
   50449: result <= 12'b111111110000;
   50450: result <= 12'b111111110000;
   50451: result <= 12'b111111110000;
   50452: result <= 12'b111111110000;
   50453: result <= 12'b111111110000;
   50454: result <= 12'b111111110000;
   50455: result <= 12'b111111110000;
   50456: result <= 12'b111111110000;
   50457: result <= 12'b111111101111;
   50458: result <= 12'b111111101111;
   50459: result <= 12'b111111101111;
   50460: result <= 12'b111111101111;
   50461: result <= 12'b111111101111;
   50462: result <= 12'b111111101111;
   50463: result <= 12'b111111101111;
   50464: result <= 12'b111111101111;
   50465: result <= 12'b111111101111;
   50466: result <= 12'b111111101111;
   50467: result <= 12'b111111101111;
   50468: result <= 12'b111111101111;
   50469: result <= 12'b111111101111;
   50470: result <= 12'b111111101111;
   50471: result <= 12'b111111101111;
   50472: result <= 12'b111111101111;
   50473: result <= 12'b111111101111;
   50474: result <= 12'b111111101111;
   50475: result <= 12'b111111101111;
   50476: result <= 12'b111111101111;
   50477: result <= 12'b111111101111;
   50478: result <= 12'b111111101111;
   50479: result <= 12'b111111101111;
   50480: result <= 12'b111111101111;
   50481: result <= 12'b111111101111;
   50482: result <= 12'b111111101111;
   50483: result <= 12'b111111101111;
   50484: result <= 12'b111111101111;
   50485: result <= 12'b111111101111;
   50486: result <= 12'b111111101111;
   50487: result <= 12'b111111101111;
   50488: result <= 12'b111111101111;
   50489: result <= 12'b111111101111;
   50490: result <= 12'b111111101111;
   50491: result <= 12'b111111101111;
   50492: result <= 12'b111111101111;
   50493: result <= 12'b111111101111;
   50494: result <= 12'b111111101111;
   50495: result <= 12'b111111101111;
   50496: result <= 12'b111111101111;
   50497: result <= 12'b111111101110;
   50498: result <= 12'b111111101110;
   50499: result <= 12'b111111101110;
   50500: result <= 12'b111111101110;
   50501: result <= 12'b111111101110;
   50502: result <= 12'b111111101110;
   50503: result <= 12'b111111101110;
   50504: result <= 12'b111111101110;
   50505: result <= 12'b111111101110;
   50506: result <= 12'b111111101110;
   50507: result <= 12'b111111101110;
   50508: result <= 12'b111111101110;
   50509: result <= 12'b111111101110;
   50510: result <= 12'b111111101110;
   50511: result <= 12'b111111101110;
   50512: result <= 12'b111111101110;
   50513: result <= 12'b111111101110;
   50514: result <= 12'b111111101110;
   50515: result <= 12'b111111101110;
   50516: result <= 12'b111111101110;
   50517: result <= 12'b111111101110;
   50518: result <= 12'b111111101110;
   50519: result <= 12'b111111101110;
   50520: result <= 12'b111111101110;
   50521: result <= 12'b111111101110;
   50522: result <= 12'b111111101110;
   50523: result <= 12'b111111101110;
   50524: result <= 12'b111111101110;
   50525: result <= 12'b111111101110;
   50526: result <= 12'b111111101110;
   50527: result <= 12'b111111101110;
   50528: result <= 12'b111111101110;
   50529: result <= 12'b111111101110;
   50530: result <= 12'b111111101110;
   50531: result <= 12'b111111101110;
   50532: result <= 12'b111111101110;
   50533: result <= 12'b111111101110;
   50534: result <= 12'b111111101110;
   50535: result <= 12'b111111101110;
   50536: result <= 12'b111111101101;
   50537: result <= 12'b111111101101;
   50538: result <= 12'b111111101101;
   50539: result <= 12'b111111101101;
   50540: result <= 12'b111111101101;
   50541: result <= 12'b111111101101;
   50542: result <= 12'b111111101101;
   50543: result <= 12'b111111101101;
   50544: result <= 12'b111111101101;
   50545: result <= 12'b111111101101;
   50546: result <= 12'b111111101101;
   50547: result <= 12'b111111101101;
   50548: result <= 12'b111111101101;
   50549: result <= 12'b111111101101;
   50550: result <= 12'b111111101101;
   50551: result <= 12'b111111101101;
   50552: result <= 12'b111111101101;
   50553: result <= 12'b111111101101;
   50554: result <= 12'b111111101101;
   50555: result <= 12'b111111101101;
   50556: result <= 12'b111111101101;
   50557: result <= 12'b111111101101;
   50558: result <= 12'b111111101101;
   50559: result <= 12'b111111101101;
   50560: result <= 12'b111111101101;
   50561: result <= 12'b111111101101;
   50562: result <= 12'b111111101101;
   50563: result <= 12'b111111101101;
   50564: result <= 12'b111111101101;
   50565: result <= 12'b111111101101;
   50566: result <= 12'b111111101101;
   50567: result <= 12'b111111101101;
   50568: result <= 12'b111111101101;
   50569: result <= 12'b111111101101;
   50570: result <= 12'b111111101101;
   50571: result <= 12'b111111101101;
   50572: result <= 12'b111111101101;
   50573: result <= 12'b111111101101;
   50574: result <= 12'b111111101100;
   50575: result <= 12'b111111101100;
   50576: result <= 12'b111111101100;
   50577: result <= 12'b111111101100;
   50578: result <= 12'b111111101100;
   50579: result <= 12'b111111101100;
   50580: result <= 12'b111111101100;
   50581: result <= 12'b111111101100;
   50582: result <= 12'b111111101100;
   50583: result <= 12'b111111101100;
   50584: result <= 12'b111111101100;
   50585: result <= 12'b111111101100;
   50586: result <= 12'b111111101100;
   50587: result <= 12'b111111101100;
   50588: result <= 12'b111111101100;
   50589: result <= 12'b111111101100;
   50590: result <= 12'b111111101100;
   50591: result <= 12'b111111101100;
   50592: result <= 12'b111111101100;
   50593: result <= 12'b111111101100;
   50594: result <= 12'b111111101100;
   50595: result <= 12'b111111101100;
   50596: result <= 12'b111111101100;
   50597: result <= 12'b111111101100;
   50598: result <= 12'b111111101100;
   50599: result <= 12'b111111101100;
   50600: result <= 12'b111111101100;
   50601: result <= 12'b111111101100;
   50602: result <= 12'b111111101100;
   50603: result <= 12'b111111101100;
   50604: result <= 12'b111111101100;
   50605: result <= 12'b111111101100;
   50606: result <= 12'b111111101100;
   50607: result <= 12'b111111101100;
   50608: result <= 12'b111111101100;
   50609: result <= 12'b111111101100;
   50610: result <= 12'b111111101100;
   50611: result <= 12'b111111101011;
   50612: result <= 12'b111111101011;
   50613: result <= 12'b111111101011;
   50614: result <= 12'b111111101011;
   50615: result <= 12'b111111101011;
   50616: result <= 12'b111111101011;
   50617: result <= 12'b111111101011;
   50618: result <= 12'b111111101011;
   50619: result <= 12'b111111101011;
   50620: result <= 12'b111111101011;
   50621: result <= 12'b111111101011;
   50622: result <= 12'b111111101011;
   50623: result <= 12'b111111101011;
   50624: result <= 12'b111111101011;
   50625: result <= 12'b111111101011;
   50626: result <= 12'b111111101011;
   50627: result <= 12'b111111101011;
   50628: result <= 12'b111111101011;
   50629: result <= 12'b111111101011;
   50630: result <= 12'b111111101011;
   50631: result <= 12'b111111101011;
   50632: result <= 12'b111111101011;
   50633: result <= 12'b111111101011;
   50634: result <= 12'b111111101011;
   50635: result <= 12'b111111101011;
   50636: result <= 12'b111111101011;
   50637: result <= 12'b111111101011;
   50638: result <= 12'b111111101011;
   50639: result <= 12'b111111101011;
   50640: result <= 12'b111111101011;
   50641: result <= 12'b111111101011;
   50642: result <= 12'b111111101011;
   50643: result <= 12'b111111101011;
   50644: result <= 12'b111111101011;
   50645: result <= 12'b111111101011;
   50646: result <= 12'b111111101011;
   50647: result <= 12'b111111101010;
   50648: result <= 12'b111111101010;
   50649: result <= 12'b111111101010;
   50650: result <= 12'b111111101010;
   50651: result <= 12'b111111101010;
   50652: result <= 12'b111111101010;
   50653: result <= 12'b111111101010;
   50654: result <= 12'b111111101010;
   50655: result <= 12'b111111101010;
   50656: result <= 12'b111111101010;
   50657: result <= 12'b111111101010;
   50658: result <= 12'b111111101010;
   50659: result <= 12'b111111101010;
   50660: result <= 12'b111111101010;
   50661: result <= 12'b111111101010;
   50662: result <= 12'b111111101010;
   50663: result <= 12'b111111101010;
   50664: result <= 12'b111111101010;
   50665: result <= 12'b111111101010;
   50666: result <= 12'b111111101010;
   50667: result <= 12'b111111101010;
   50668: result <= 12'b111111101010;
   50669: result <= 12'b111111101010;
   50670: result <= 12'b111111101010;
   50671: result <= 12'b111111101010;
   50672: result <= 12'b111111101010;
   50673: result <= 12'b111111101010;
   50674: result <= 12'b111111101010;
   50675: result <= 12'b111111101010;
   50676: result <= 12'b111111101010;
   50677: result <= 12'b111111101010;
   50678: result <= 12'b111111101010;
   50679: result <= 12'b111111101010;
   50680: result <= 12'b111111101010;
   50681: result <= 12'b111111101010;
   50682: result <= 12'b111111101010;
   50683: result <= 12'b111111101001;
   50684: result <= 12'b111111101001;
   50685: result <= 12'b111111101001;
   50686: result <= 12'b111111101001;
   50687: result <= 12'b111111101001;
   50688: result <= 12'b111111101001;
   50689: result <= 12'b111111101001;
   50690: result <= 12'b111111101001;
   50691: result <= 12'b111111101001;
   50692: result <= 12'b111111101001;
   50693: result <= 12'b111111101001;
   50694: result <= 12'b111111101001;
   50695: result <= 12'b111111101001;
   50696: result <= 12'b111111101001;
   50697: result <= 12'b111111101001;
   50698: result <= 12'b111111101001;
   50699: result <= 12'b111111101001;
   50700: result <= 12'b111111101001;
   50701: result <= 12'b111111101001;
   50702: result <= 12'b111111101001;
   50703: result <= 12'b111111101001;
   50704: result <= 12'b111111101001;
   50705: result <= 12'b111111101001;
   50706: result <= 12'b111111101001;
   50707: result <= 12'b111111101001;
   50708: result <= 12'b111111101001;
   50709: result <= 12'b111111101001;
   50710: result <= 12'b111111101001;
   50711: result <= 12'b111111101001;
   50712: result <= 12'b111111101001;
   50713: result <= 12'b111111101001;
   50714: result <= 12'b111111101001;
   50715: result <= 12'b111111101001;
   50716: result <= 12'b111111101001;
   50717: result <= 12'b111111101000;
   50718: result <= 12'b111111101000;
   50719: result <= 12'b111111101000;
   50720: result <= 12'b111111101000;
   50721: result <= 12'b111111101000;
   50722: result <= 12'b111111101000;
   50723: result <= 12'b111111101000;
   50724: result <= 12'b111111101000;
   50725: result <= 12'b111111101000;
   50726: result <= 12'b111111101000;
   50727: result <= 12'b111111101000;
   50728: result <= 12'b111111101000;
   50729: result <= 12'b111111101000;
   50730: result <= 12'b111111101000;
   50731: result <= 12'b111111101000;
   50732: result <= 12'b111111101000;
   50733: result <= 12'b111111101000;
   50734: result <= 12'b111111101000;
   50735: result <= 12'b111111101000;
   50736: result <= 12'b111111101000;
   50737: result <= 12'b111111101000;
   50738: result <= 12'b111111101000;
   50739: result <= 12'b111111101000;
   50740: result <= 12'b111111101000;
   50741: result <= 12'b111111101000;
   50742: result <= 12'b111111101000;
   50743: result <= 12'b111111101000;
   50744: result <= 12'b111111101000;
   50745: result <= 12'b111111101000;
   50746: result <= 12'b111111101000;
   50747: result <= 12'b111111101000;
   50748: result <= 12'b111111101000;
   50749: result <= 12'b111111101000;
   50750: result <= 12'b111111101000;
   50751: result <= 12'b111111100111;
   50752: result <= 12'b111111100111;
   50753: result <= 12'b111111100111;
   50754: result <= 12'b111111100111;
   50755: result <= 12'b111111100111;
   50756: result <= 12'b111111100111;
   50757: result <= 12'b111111100111;
   50758: result <= 12'b111111100111;
   50759: result <= 12'b111111100111;
   50760: result <= 12'b111111100111;
   50761: result <= 12'b111111100111;
   50762: result <= 12'b111111100111;
   50763: result <= 12'b111111100111;
   50764: result <= 12'b111111100111;
   50765: result <= 12'b111111100111;
   50766: result <= 12'b111111100111;
   50767: result <= 12'b111111100111;
   50768: result <= 12'b111111100111;
   50769: result <= 12'b111111100111;
   50770: result <= 12'b111111100111;
   50771: result <= 12'b111111100111;
   50772: result <= 12'b111111100111;
   50773: result <= 12'b111111100111;
   50774: result <= 12'b111111100111;
   50775: result <= 12'b111111100111;
   50776: result <= 12'b111111100111;
   50777: result <= 12'b111111100111;
   50778: result <= 12'b111111100111;
   50779: result <= 12'b111111100111;
   50780: result <= 12'b111111100111;
   50781: result <= 12'b111111100111;
   50782: result <= 12'b111111100111;
   50783: result <= 12'b111111100111;
   50784: result <= 12'b111111100110;
   50785: result <= 12'b111111100110;
   50786: result <= 12'b111111100110;
   50787: result <= 12'b111111100110;
   50788: result <= 12'b111111100110;
   50789: result <= 12'b111111100110;
   50790: result <= 12'b111111100110;
   50791: result <= 12'b111111100110;
   50792: result <= 12'b111111100110;
   50793: result <= 12'b111111100110;
   50794: result <= 12'b111111100110;
   50795: result <= 12'b111111100110;
   50796: result <= 12'b111111100110;
   50797: result <= 12'b111111100110;
   50798: result <= 12'b111111100110;
   50799: result <= 12'b111111100110;
   50800: result <= 12'b111111100110;
   50801: result <= 12'b111111100110;
   50802: result <= 12'b111111100110;
   50803: result <= 12'b111111100110;
   50804: result <= 12'b111111100110;
   50805: result <= 12'b111111100110;
   50806: result <= 12'b111111100110;
   50807: result <= 12'b111111100110;
   50808: result <= 12'b111111100110;
   50809: result <= 12'b111111100110;
   50810: result <= 12'b111111100110;
   50811: result <= 12'b111111100110;
   50812: result <= 12'b111111100110;
   50813: result <= 12'b111111100110;
   50814: result <= 12'b111111100110;
   50815: result <= 12'b111111100110;
   50816: result <= 12'b111111100101;
   50817: result <= 12'b111111100101;
   50818: result <= 12'b111111100101;
   50819: result <= 12'b111111100101;
   50820: result <= 12'b111111100101;
   50821: result <= 12'b111111100101;
   50822: result <= 12'b111111100101;
   50823: result <= 12'b111111100101;
   50824: result <= 12'b111111100101;
   50825: result <= 12'b111111100101;
   50826: result <= 12'b111111100101;
   50827: result <= 12'b111111100101;
   50828: result <= 12'b111111100101;
   50829: result <= 12'b111111100101;
   50830: result <= 12'b111111100101;
   50831: result <= 12'b111111100101;
   50832: result <= 12'b111111100101;
   50833: result <= 12'b111111100101;
   50834: result <= 12'b111111100101;
   50835: result <= 12'b111111100101;
   50836: result <= 12'b111111100101;
   50837: result <= 12'b111111100101;
   50838: result <= 12'b111111100101;
   50839: result <= 12'b111111100101;
   50840: result <= 12'b111111100101;
   50841: result <= 12'b111111100101;
   50842: result <= 12'b111111100101;
   50843: result <= 12'b111111100101;
   50844: result <= 12'b111111100101;
   50845: result <= 12'b111111100101;
   50846: result <= 12'b111111100101;
   50847: result <= 12'b111111100101;
   50848: result <= 12'b111111100100;
   50849: result <= 12'b111111100100;
   50850: result <= 12'b111111100100;
   50851: result <= 12'b111111100100;
   50852: result <= 12'b111111100100;
   50853: result <= 12'b111111100100;
   50854: result <= 12'b111111100100;
   50855: result <= 12'b111111100100;
   50856: result <= 12'b111111100100;
   50857: result <= 12'b111111100100;
   50858: result <= 12'b111111100100;
   50859: result <= 12'b111111100100;
   50860: result <= 12'b111111100100;
   50861: result <= 12'b111111100100;
   50862: result <= 12'b111111100100;
   50863: result <= 12'b111111100100;
   50864: result <= 12'b111111100100;
   50865: result <= 12'b111111100100;
   50866: result <= 12'b111111100100;
   50867: result <= 12'b111111100100;
   50868: result <= 12'b111111100100;
   50869: result <= 12'b111111100100;
   50870: result <= 12'b111111100100;
   50871: result <= 12'b111111100100;
   50872: result <= 12'b111111100100;
   50873: result <= 12'b111111100100;
   50874: result <= 12'b111111100100;
   50875: result <= 12'b111111100100;
   50876: result <= 12'b111111100100;
   50877: result <= 12'b111111100100;
   50878: result <= 12'b111111100100;
   50879: result <= 12'b111111100011;
   50880: result <= 12'b111111100011;
   50881: result <= 12'b111111100011;
   50882: result <= 12'b111111100011;
   50883: result <= 12'b111111100011;
   50884: result <= 12'b111111100011;
   50885: result <= 12'b111111100011;
   50886: result <= 12'b111111100011;
   50887: result <= 12'b111111100011;
   50888: result <= 12'b111111100011;
   50889: result <= 12'b111111100011;
   50890: result <= 12'b111111100011;
   50891: result <= 12'b111111100011;
   50892: result <= 12'b111111100011;
   50893: result <= 12'b111111100011;
   50894: result <= 12'b111111100011;
   50895: result <= 12'b111111100011;
   50896: result <= 12'b111111100011;
   50897: result <= 12'b111111100011;
   50898: result <= 12'b111111100011;
   50899: result <= 12'b111111100011;
   50900: result <= 12'b111111100011;
   50901: result <= 12'b111111100011;
   50902: result <= 12'b111111100011;
   50903: result <= 12'b111111100011;
   50904: result <= 12'b111111100011;
   50905: result <= 12'b111111100011;
   50906: result <= 12'b111111100011;
   50907: result <= 12'b111111100011;
   50908: result <= 12'b111111100011;
   50909: result <= 12'b111111100011;
   50910: result <= 12'b111111100010;
   50911: result <= 12'b111111100010;
   50912: result <= 12'b111111100010;
   50913: result <= 12'b111111100010;
   50914: result <= 12'b111111100010;
   50915: result <= 12'b111111100010;
   50916: result <= 12'b111111100010;
   50917: result <= 12'b111111100010;
   50918: result <= 12'b111111100010;
   50919: result <= 12'b111111100010;
   50920: result <= 12'b111111100010;
   50921: result <= 12'b111111100010;
   50922: result <= 12'b111111100010;
   50923: result <= 12'b111111100010;
   50924: result <= 12'b111111100010;
   50925: result <= 12'b111111100010;
   50926: result <= 12'b111111100010;
   50927: result <= 12'b111111100010;
   50928: result <= 12'b111111100010;
   50929: result <= 12'b111111100010;
   50930: result <= 12'b111111100010;
   50931: result <= 12'b111111100010;
   50932: result <= 12'b111111100010;
   50933: result <= 12'b111111100010;
   50934: result <= 12'b111111100010;
   50935: result <= 12'b111111100010;
   50936: result <= 12'b111111100010;
   50937: result <= 12'b111111100010;
   50938: result <= 12'b111111100010;
   50939: result <= 12'b111111100010;
   50940: result <= 12'b111111100001;
   50941: result <= 12'b111111100001;
   50942: result <= 12'b111111100001;
   50943: result <= 12'b111111100001;
   50944: result <= 12'b111111100001;
   50945: result <= 12'b111111100001;
   50946: result <= 12'b111111100001;
   50947: result <= 12'b111111100001;
   50948: result <= 12'b111111100001;
   50949: result <= 12'b111111100001;
   50950: result <= 12'b111111100001;
   50951: result <= 12'b111111100001;
   50952: result <= 12'b111111100001;
   50953: result <= 12'b111111100001;
   50954: result <= 12'b111111100001;
   50955: result <= 12'b111111100001;
   50956: result <= 12'b111111100001;
   50957: result <= 12'b111111100001;
   50958: result <= 12'b111111100001;
   50959: result <= 12'b111111100001;
   50960: result <= 12'b111111100001;
   50961: result <= 12'b111111100001;
   50962: result <= 12'b111111100001;
   50963: result <= 12'b111111100001;
   50964: result <= 12'b111111100001;
   50965: result <= 12'b111111100001;
   50966: result <= 12'b111111100001;
   50967: result <= 12'b111111100001;
   50968: result <= 12'b111111100001;
   50969: result <= 12'b111111100001;
   50970: result <= 12'b111111100000;
   50971: result <= 12'b111111100000;
   50972: result <= 12'b111111100000;
   50973: result <= 12'b111111100000;
   50974: result <= 12'b111111100000;
   50975: result <= 12'b111111100000;
   50976: result <= 12'b111111100000;
   50977: result <= 12'b111111100000;
   50978: result <= 12'b111111100000;
   50979: result <= 12'b111111100000;
   50980: result <= 12'b111111100000;
   50981: result <= 12'b111111100000;
   50982: result <= 12'b111111100000;
   50983: result <= 12'b111111100000;
   50984: result <= 12'b111111100000;
   50985: result <= 12'b111111100000;
   50986: result <= 12'b111111100000;
   50987: result <= 12'b111111100000;
   50988: result <= 12'b111111100000;
   50989: result <= 12'b111111100000;
   50990: result <= 12'b111111100000;
   50991: result <= 12'b111111100000;
   50992: result <= 12'b111111100000;
   50993: result <= 12'b111111100000;
   50994: result <= 12'b111111100000;
   50995: result <= 12'b111111100000;
   50996: result <= 12'b111111100000;
   50997: result <= 12'b111111100000;
   50998: result <= 12'b111111100000;
   50999: result <= 12'b111111011111;
   51000: result <= 12'b111111011111;
   51001: result <= 12'b111111011111;
   51002: result <= 12'b111111011111;
   51003: result <= 12'b111111011111;
   51004: result <= 12'b111111011111;
   51005: result <= 12'b111111011111;
   51006: result <= 12'b111111011111;
   51007: result <= 12'b111111011111;
   51008: result <= 12'b111111011111;
   51009: result <= 12'b111111011111;
   51010: result <= 12'b111111011111;
   51011: result <= 12'b111111011111;
   51012: result <= 12'b111111011111;
   51013: result <= 12'b111111011111;
   51014: result <= 12'b111111011111;
   51015: result <= 12'b111111011111;
   51016: result <= 12'b111111011111;
   51017: result <= 12'b111111011111;
   51018: result <= 12'b111111011111;
   51019: result <= 12'b111111011111;
   51020: result <= 12'b111111011111;
   51021: result <= 12'b111111011111;
   51022: result <= 12'b111111011111;
   51023: result <= 12'b111111011111;
   51024: result <= 12'b111111011111;
   51025: result <= 12'b111111011111;
   51026: result <= 12'b111111011111;
   51027: result <= 12'b111111011110;
   51028: result <= 12'b111111011110;
   51029: result <= 12'b111111011110;
   51030: result <= 12'b111111011110;
   51031: result <= 12'b111111011110;
   51032: result <= 12'b111111011110;
   51033: result <= 12'b111111011110;
   51034: result <= 12'b111111011110;
   51035: result <= 12'b111111011110;
   51036: result <= 12'b111111011110;
   51037: result <= 12'b111111011110;
   51038: result <= 12'b111111011110;
   51039: result <= 12'b111111011110;
   51040: result <= 12'b111111011110;
   51041: result <= 12'b111111011110;
   51042: result <= 12'b111111011110;
   51043: result <= 12'b111111011110;
   51044: result <= 12'b111111011110;
   51045: result <= 12'b111111011110;
   51046: result <= 12'b111111011110;
   51047: result <= 12'b111111011110;
   51048: result <= 12'b111111011110;
   51049: result <= 12'b111111011110;
   51050: result <= 12'b111111011110;
   51051: result <= 12'b111111011110;
   51052: result <= 12'b111111011110;
   51053: result <= 12'b111111011110;
   51054: result <= 12'b111111011110;
   51055: result <= 12'b111111011110;
   51056: result <= 12'b111111011101;
   51057: result <= 12'b111111011101;
   51058: result <= 12'b111111011101;
   51059: result <= 12'b111111011101;
   51060: result <= 12'b111111011101;
   51061: result <= 12'b111111011101;
   51062: result <= 12'b111111011101;
   51063: result <= 12'b111111011101;
   51064: result <= 12'b111111011101;
   51065: result <= 12'b111111011101;
   51066: result <= 12'b111111011101;
   51067: result <= 12'b111111011101;
   51068: result <= 12'b111111011101;
   51069: result <= 12'b111111011101;
   51070: result <= 12'b111111011101;
   51071: result <= 12'b111111011101;
   51072: result <= 12'b111111011101;
   51073: result <= 12'b111111011101;
   51074: result <= 12'b111111011101;
   51075: result <= 12'b111111011101;
   51076: result <= 12'b111111011101;
   51077: result <= 12'b111111011101;
   51078: result <= 12'b111111011101;
   51079: result <= 12'b111111011101;
   51080: result <= 12'b111111011101;
   51081: result <= 12'b111111011101;
   51082: result <= 12'b111111011101;
   51083: result <= 12'b111111011101;
   51084: result <= 12'b111111011100;
   51085: result <= 12'b111111011100;
   51086: result <= 12'b111111011100;
   51087: result <= 12'b111111011100;
   51088: result <= 12'b111111011100;
   51089: result <= 12'b111111011100;
   51090: result <= 12'b111111011100;
   51091: result <= 12'b111111011100;
   51092: result <= 12'b111111011100;
   51093: result <= 12'b111111011100;
   51094: result <= 12'b111111011100;
   51095: result <= 12'b111111011100;
   51096: result <= 12'b111111011100;
   51097: result <= 12'b111111011100;
   51098: result <= 12'b111111011100;
   51099: result <= 12'b111111011100;
   51100: result <= 12'b111111011100;
   51101: result <= 12'b111111011100;
   51102: result <= 12'b111111011100;
   51103: result <= 12'b111111011100;
   51104: result <= 12'b111111011100;
   51105: result <= 12'b111111011100;
   51106: result <= 12'b111111011100;
   51107: result <= 12'b111111011100;
   51108: result <= 12'b111111011100;
   51109: result <= 12'b111111011100;
   51110: result <= 12'b111111011100;
   51111: result <= 12'b111111011011;
   51112: result <= 12'b111111011011;
   51113: result <= 12'b111111011011;
   51114: result <= 12'b111111011011;
   51115: result <= 12'b111111011011;
   51116: result <= 12'b111111011011;
   51117: result <= 12'b111111011011;
   51118: result <= 12'b111111011011;
   51119: result <= 12'b111111011011;
   51120: result <= 12'b111111011011;
   51121: result <= 12'b111111011011;
   51122: result <= 12'b111111011011;
   51123: result <= 12'b111111011011;
   51124: result <= 12'b111111011011;
   51125: result <= 12'b111111011011;
   51126: result <= 12'b111111011011;
   51127: result <= 12'b111111011011;
   51128: result <= 12'b111111011011;
   51129: result <= 12'b111111011011;
   51130: result <= 12'b111111011011;
   51131: result <= 12'b111111011011;
   51132: result <= 12'b111111011011;
   51133: result <= 12'b111111011011;
   51134: result <= 12'b111111011011;
   51135: result <= 12'b111111011011;
   51136: result <= 12'b111111011011;
   51137: result <= 12'b111111011011;
   51138: result <= 12'b111111011010;
   51139: result <= 12'b111111011010;
   51140: result <= 12'b111111011010;
   51141: result <= 12'b111111011010;
   51142: result <= 12'b111111011010;
   51143: result <= 12'b111111011010;
   51144: result <= 12'b111111011010;
   51145: result <= 12'b111111011010;
   51146: result <= 12'b111111011010;
   51147: result <= 12'b111111011010;
   51148: result <= 12'b111111011010;
   51149: result <= 12'b111111011010;
   51150: result <= 12'b111111011010;
   51151: result <= 12'b111111011010;
   51152: result <= 12'b111111011010;
   51153: result <= 12'b111111011010;
   51154: result <= 12'b111111011010;
   51155: result <= 12'b111111011010;
   51156: result <= 12'b111111011010;
   51157: result <= 12'b111111011010;
   51158: result <= 12'b111111011010;
   51159: result <= 12'b111111011010;
   51160: result <= 12'b111111011010;
   51161: result <= 12'b111111011010;
   51162: result <= 12'b111111011010;
   51163: result <= 12'b111111011010;
   51164: result <= 12'b111111011010;
   51165: result <= 12'b111111011001;
   51166: result <= 12'b111111011001;
   51167: result <= 12'b111111011001;
   51168: result <= 12'b111111011001;
   51169: result <= 12'b111111011001;
   51170: result <= 12'b111111011001;
   51171: result <= 12'b111111011001;
   51172: result <= 12'b111111011001;
   51173: result <= 12'b111111011001;
   51174: result <= 12'b111111011001;
   51175: result <= 12'b111111011001;
   51176: result <= 12'b111111011001;
   51177: result <= 12'b111111011001;
   51178: result <= 12'b111111011001;
   51179: result <= 12'b111111011001;
   51180: result <= 12'b111111011001;
   51181: result <= 12'b111111011001;
   51182: result <= 12'b111111011001;
   51183: result <= 12'b111111011001;
   51184: result <= 12'b111111011001;
   51185: result <= 12'b111111011001;
   51186: result <= 12'b111111011001;
   51187: result <= 12'b111111011001;
   51188: result <= 12'b111111011001;
   51189: result <= 12'b111111011001;
   51190: result <= 12'b111111011001;
   51191: result <= 12'b111111011000;
   51192: result <= 12'b111111011000;
   51193: result <= 12'b111111011000;
   51194: result <= 12'b111111011000;
   51195: result <= 12'b111111011000;
   51196: result <= 12'b111111011000;
   51197: result <= 12'b111111011000;
   51198: result <= 12'b111111011000;
   51199: result <= 12'b111111011000;
   51200: result <= 12'b111111011000;
   51201: result <= 12'b111111011000;
   51202: result <= 12'b111111011000;
   51203: result <= 12'b111111011000;
   51204: result <= 12'b111111011000;
   51205: result <= 12'b111111011000;
   51206: result <= 12'b111111011000;
   51207: result <= 12'b111111011000;
   51208: result <= 12'b111111011000;
   51209: result <= 12'b111111011000;
   51210: result <= 12'b111111011000;
   51211: result <= 12'b111111011000;
   51212: result <= 12'b111111011000;
   51213: result <= 12'b111111011000;
   51214: result <= 12'b111111011000;
   51215: result <= 12'b111111011000;
   51216: result <= 12'b111111011000;
   51217: result <= 12'b111111010111;
   51218: result <= 12'b111111010111;
   51219: result <= 12'b111111010111;
   51220: result <= 12'b111111010111;
   51221: result <= 12'b111111010111;
   51222: result <= 12'b111111010111;
   51223: result <= 12'b111111010111;
   51224: result <= 12'b111111010111;
   51225: result <= 12'b111111010111;
   51226: result <= 12'b111111010111;
   51227: result <= 12'b111111010111;
   51228: result <= 12'b111111010111;
   51229: result <= 12'b111111010111;
   51230: result <= 12'b111111010111;
   51231: result <= 12'b111111010111;
   51232: result <= 12'b111111010111;
   51233: result <= 12'b111111010111;
   51234: result <= 12'b111111010111;
   51235: result <= 12'b111111010111;
   51236: result <= 12'b111111010111;
   51237: result <= 12'b111111010111;
   51238: result <= 12'b111111010111;
   51239: result <= 12'b111111010111;
   51240: result <= 12'b111111010111;
   51241: result <= 12'b111111010111;
   51242: result <= 12'b111111010111;
   51243: result <= 12'b111111010110;
   51244: result <= 12'b111111010110;
   51245: result <= 12'b111111010110;
   51246: result <= 12'b111111010110;
   51247: result <= 12'b111111010110;
   51248: result <= 12'b111111010110;
   51249: result <= 12'b111111010110;
   51250: result <= 12'b111111010110;
   51251: result <= 12'b111111010110;
   51252: result <= 12'b111111010110;
   51253: result <= 12'b111111010110;
   51254: result <= 12'b111111010110;
   51255: result <= 12'b111111010110;
   51256: result <= 12'b111111010110;
   51257: result <= 12'b111111010110;
   51258: result <= 12'b111111010110;
   51259: result <= 12'b111111010110;
   51260: result <= 12'b111111010110;
   51261: result <= 12'b111111010110;
   51262: result <= 12'b111111010110;
   51263: result <= 12'b111111010110;
   51264: result <= 12'b111111010110;
   51265: result <= 12'b111111010110;
   51266: result <= 12'b111111010110;
   51267: result <= 12'b111111010110;
   51268: result <= 12'b111111010110;
   51269: result <= 12'b111111010101;
   51270: result <= 12'b111111010101;
   51271: result <= 12'b111111010101;
   51272: result <= 12'b111111010101;
   51273: result <= 12'b111111010101;
   51274: result <= 12'b111111010101;
   51275: result <= 12'b111111010101;
   51276: result <= 12'b111111010101;
   51277: result <= 12'b111111010101;
   51278: result <= 12'b111111010101;
   51279: result <= 12'b111111010101;
   51280: result <= 12'b111111010101;
   51281: result <= 12'b111111010101;
   51282: result <= 12'b111111010101;
   51283: result <= 12'b111111010101;
   51284: result <= 12'b111111010101;
   51285: result <= 12'b111111010101;
   51286: result <= 12'b111111010101;
   51287: result <= 12'b111111010101;
   51288: result <= 12'b111111010101;
   51289: result <= 12'b111111010101;
   51290: result <= 12'b111111010101;
   51291: result <= 12'b111111010101;
   51292: result <= 12'b111111010101;
   51293: result <= 12'b111111010101;
   51294: result <= 12'b111111010100;
   51295: result <= 12'b111111010100;
   51296: result <= 12'b111111010100;
   51297: result <= 12'b111111010100;
   51298: result <= 12'b111111010100;
   51299: result <= 12'b111111010100;
   51300: result <= 12'b111111010100;
   51301: result <= 12'b111111010100;
   51302: result <= 12'b111111010100;
   51303: result <= 12'b111111010100;
   51304: result <= 12'b111111010100;
   51305: result <= 12'b111111010100;
   51306: result <= 12'b111111010100;
   51307: result <= 12'b111111010100;
   51308: result <= 12'b111111010100;
   51309: result <= 12'b111111010100;
   51310: result <= 12'b111111010100;
   51311: result <= 12'b111111010100;
   51312: result <= 12'b111111010100;
   51313: result <= 12'b111111010100;
   51314: result <= 12'b111111010100;
   51315: result <= 12'b111111010100;
   51316: result <= 12'b111111010100;
   51317: result <= 12'b111111010100;
   51318: result <= 12'b111111010011;
   51319: result <= 12'b111111010011;
   51320: result <= 12'b111111010011;
   51321: result <= 12'b111111010011;
   51322: result <= 12'b111111010011;
   51323: result <= 12'b111111010011;
   51324: result <= 12'b111111010011;
   51325: result <= 12'b111111010011;
   51326: result <= 12'b111111010011;
   51327: result <= 12'b111111010011;
   51328: result <= 12'b111111010011;
   51329: result <= 12'b111111010011;
   51330: result <= 12'b111111010011;
   51331: result <= 12'b111111010011;
   51332: result <= 12'b111111010011;
   51333: result <= 12'b111111010011;
   51334: result <= 12'b111111010011;
   51335: result <= 12'b111111010011;
   51336: result <= 12'b111111010011;
   51337: result <= 12'b111111010011;
   51338: result <= 12'b111111010011;
   51339: result <= 12'b111111010011;
   51340: result <= 12'b111111010011;
   51341: result <= 12'b111111010011;
   51342: result <= 12'b111111010011;
   51343: result <= 12'b111111010010;
   51344: result <= 12'b111111010010;
   51345: result <= 12'b111111010010;
   51346: result <= 12'b111111010010;
   51347: result <= 12'b111111010010;
   51348: result <= 12'b111111010010;
   51349: result <= 12'b111111010010;
   51350: result <= 12'b111111010010;
   51351: result <= 12'b111111010010;
   51352: result <= 12'b111111010010;
   51353: result <= 12'b111111010010;
   51354: result <= 12'b111111010010;
   51355: result <= 12'b111111010010;
   51356: result <= 12'b111111010010;
   51357: result <= 12'b111111010010;
   51358: result <= 12'b111111010010;
   51359: result <= 12'b111111010010;
   51360: result <= 12'b111111010010;
   51361: result <= 12'b111111010010;
   51362: result <= 12'b111111010010;
   51363: result <= 12'b111111010010;
   51364: result <= 12'b111111010010;
   51365: result <= 12'b111111010010;
   51366: result <= 12'b111111010010;
   51367: result <= 12'b111111010001;
   51368: result <= 12'b111111010001;
   51369: result <= 12'b111111010001;
   51370: result <= 12'b111111010001;
   51371: result <= 12'b111111010001;
   51372: result <= 12'b111111010001;
   51373: result <= 12'b111111010001;
   51374: result <= 12'b111111010001;
   51375: result <= 12'b111111010001;
   51376: result <= 12'b111111010001;
   51377: result <= 12'b111111010001;
   51378: result <= 12'b111111010001;
   51379: result <= 12'b111111010001;
   51380: result <= 12'b111111010001;
   51381: result <= 12'b111111010001;
   51382: result <= 12'b111111010001;
   51383: result <= 12'b111111010001;
   51384: result <= 12'b111111010001;
   51385: result <= 12'b111111010001;
   51386: result <= 12'b111111010001;
   51387: result <= 12'b111111010001;
   51388: result <= 12'b111111010001;
   51389: result <= 12'b111111010001;
   51390: result <= 12'b111111010001;
   51391: result <= 12'b111111010000;
   51392: result <= 12'b111111010000;
   51393: result <= 12'b111111010000;
   51394: result <= 12'b111111010000;
   51395: result <= 12'b111111010000;
   51396: result <= 12'b111111010000;
   51397: result <= 12'b111111010000;
   51398: result <= 12'b111111010000;
   51399: result <= 12'b111111010000;
   51400: result <= 12'b111111010000;
   51401: result <= 12'b111111010000;
   51402: result <= 12'b111111010000;
   51403: result <= 12'b111111010000;
   51404: result <= 12'b111111010000;
   51405: result <= 12'b111111010000;
   51406: result <= 12'b111111010000;
   51407: result <= 12'b111111010000;
   51408: result <= 12'b111111010000;
   51409: result <= 12'b111111010000;
   51410: result <= 12'b111111010000;
   51411: result <= 12'b111111010000;
   51412: result <= 12'b111111010000;
   51413: result <= 12'b111111010000;
   51414: result <= 12'b111111010000;
   51415: result <= 12'b111111001111;
   51416: result <= 12'b111111001111;
   51417: result <= 12'b111111001111;
   51418: result <= 12'b111111001111;
   51419: result <= 12'b111111001111;
   51420: result <= 12'b111111001111;
   51421: result <= 12'b111111001111;
   51422: result <= 12'b111111001111;
   51423: result <= 12'b111111001111;
   51424: result <= 12'b111111001111;
   51425: result <= 12'b111111001111;
   51426: result <= 12'b111111001111;
   51427: result <= 12'b111111001111;
   51428: result <= 12'b111111001111;
   51429: result <= 12'b111111001111;
   51430: result <= 12'b111111001111;
   51431: result <= 12'b111111001111;
   51432: result <= 12'b111111001111;
   51433: result <= 12'b111111001111;
   51434: result <= 12'b111111001111;
   51435: result <= 12'b111111001111;
   51436: result <= 12'b111111001111;
   51437: result <= 12'b111111001111;
   51438: result <= 12'b111111001111;
   51439: result <= 12'b111111001110;
   51440: result <= 12'b111111001110;
   51441: result <= 12'b111111001110;
   51442: result <= 12'b111111001110;
   51443: result <= 12'b111111001110;
   51444: result <= 12'b111111001110;
   51445: result <= 12'b111111001110;
   51446: result <= 12'b111111001110;
   51447: result <= 12'b111111001110;
   51448: result <= 12'b111111001110;
   51449: result <= 12'b111111001110;
   51450: result <= 12'b111111001110;
   51451: result <= 12'b111111001110;
   51452: result <= 12'b111111001110;
   51453: result <= 12'b111111001110;
   51454: result <= 12'b111111001110;
   51455: result <= 12'b111111001110;
   51456: result <= 12'b111111001110;
   51457: result <= 12'b111111001110;
   51458: result <= 12'b111111001110;
   51459: result <= 12'b111111001110;
   51460: result <= 12'b111111001110;
   51461: result <= 12'b111111001110;
   51462: result <= 12'b111111001101;
   51463: result <= 12'b111111001101;
   51464: result <= 12'b111111001101;
   51465: result <= 12'b111111001101;
   51466: result <= 12'b111111001101;
   51467: result <= 12'b111111001101;
   51468: result <= 12'b111111001101;
   51469: result <= 12'b111111001101;
   51470: result <= 12'b111111001101;
   51471: result <= 12'b111111001101;
   51472: result <= 12'b111111001101;
   51473: result <= 12'b111111001101;
   51474: result <= 12'b111111001101;
   51475: result <= 12'b111111001101;
   51476: result <= 12'b111111001101;
   51477: result <= 12'b111111001101;
   51478: result <= 12'b111111001101;
   51479: result <= 12'b111111001101;
   51480: result <= 12'b111111001101;
   51481: result <= 12'b111111001101;
   51482: result <= 12'b111111001101;
   51483: result <= 12'b111111001101;
   51484: result <= 12'b111111001101;
   51485: result <= 12'b111111001100;
   51486: result <= 12'b111111001100;
   51487: result <= 12'b111111001100;
   51488: result <= 12'b111111001100;
   51489: result <= 12'b111111001100;
   51490: result <= 12'b111111001100;
   51491: result <= 12'b111111001100;
   51492: result <= 12'b111111001100;
   51493: result <= 12'b111111001100;
   51494: result <= 12'b111111001100;
   51495: result <= 12'b111111001100;
   51496: result <= 12'b111111001100;
   51497: result <= 12'b111111001100;
   51498: result <= 12'b111111001100;
   51499: result <= 12'b111111001100;
   51500: result <= 12'b111111001100;
   51501: result <= 12'b111111001100;
   51502: result <= 12'b111111001100;
   51503: result <= 12'b111111001100;
   51504: result <= 12'b111111001100;
   51505: result <= 12'b111111001100;
   51506: result <= 12'b111111001100;
   51507: result <= 12'b111111001100;
   51508: result <= 12'b111111001011;
   51509: result <= 12'b111111001011;
   51510: result <= 12'b111111001011;
   51511: result <= 12'b111111001011;
   51512: result <= 12'b111111001011;
   51513: result <= 12'b111111001011;
   51514: result <= 12'b111111001011;
   51515: result <= 12'b111111001011;
   51516: result <= 12'b111111001011;
   51517: result <= 12'b111111001011;
   51518: result <= 12'b111111001011;
   51519: result <= 12'b111111001011;
   51520: result <= 12'b111111001011;
   51521: result <= 12'b111111001011;
   51522: result <= 12'b111111001011;
   51523: result <= 12'b111111001011;
   51524: result <= 12'b111111001011;
   51525: result <= 12'b111111001011;
   51526: result <= 12'b111111001011;
   51527: result <= 12'b111111001011;
   51528: result <= 12'b111111001011;
   51529: result <= 12'b111111001011;
   51530: result <= 12'b111111001011;
   51531: result <= 12'b111111001010;
   51532: result <= 12'b111111001010;
   51533: result <= 12'b111111001010;
   51534: result <= 12'b111111001010;
   51535: result <= 12'b111111001010;
   51536: result <= 12'b111111001010;
   51537: result <= 12'b111111001010;
   51538: result <= 12'b111111001010;
   51539: result <= 12'b111111001010;
   51540: result <= 12'b111111001010;
   51541: result <= 12'b111111001010;
   51542: result <= 12'b111111001010;
   51543: result <= 12'b111111001010;
   51544: result <= 12'b111111001010;
   51545: result <= 12'b111111001010;
   51546: result <= 12'b111111001010;
   51547: result <= 12'b111111001010;
   51548: result <= 12'b111111001010;
   51549: result <= 12'b111111001010;
   51550: result <= 12'b111111001010;
   51551: result <= 12'b111111001010;
   51552: result <= 12'b111111001010;
   51553: result <= 12'b111111001001;
   51554: result <= 12'b111111001001;
   51555: result <= 12'b111111001001;
   51556: result <= 12'b111111001001;
   51557: result <= 12'b111111001001;
   51558: result <= 12'b111111001001;
   51559: result <= 12'b111111001001;
   51560: result <= 12'b111111001001;
   51561: result <= 12'b111111001001;
   51562: result <= 12'b111111001001;
   51563: result <= 12'b111111001001;
   51564: result <= 12'b111111001001;
   51565: result <= 12'b111111001001;
   51566: result <= 12'b111111001001;
   51567: result <= 12'b111111001001;
   51568: result <= 12'b111111001001;
   51569: result <= 12'b111111001001;
   51570: result <= 12'b111111001001;
   51571: result <= 12'b111111001001;
   51572: result <= 12'b111111001001;
   51573: result <= 12'b111111001001;
   51574: result <= 12'b111111001001;
   51575: result <= 12'b111111001000;
   51576: result <= 12'b111111001000;
   51577: result <= 12'b111111001000;
   51578: result <= 12'b111111001000;
   51579: result <= 12'b111111001000;
   51580: result <= 12'b111111001000;
   51581: result <= 12'b111111001000;
   51582: result <= 12'b111111001000;
   51583: result <= 12'b111111001000;
   51584: result <= 12'b111111001000;
   51585: result <= 12'b111111001000;
   51586: result <= 12'b111111001000;
   51587: result <= 12'b111111001000;
   51588: result <= 12'b111111001000;
   51589: result <= 12'b111111001000;
   51590: result <= 12'b111111001000;
   51591: result <= 12'b111111001000;
   51592: result <= 12'b111111001000;
   51593: result <= 12'b111111001000;
   51594: result <= 12'b111111001000;
   51595: result <= 12'b111111001000;
   51596: result <= 12'b111111001000;
   51597: result <= 12'b111111000111;
   51598: result <= 12'b111111000111;
   51599: result <= 12'b111111000111;
   51600: result <= 12'b111111000111;
   51601: result <= 12'b111111000111;
   51602: result <= 12'b111111000111;
   51603: result <= 12'b111111000111;
   51604: result <= 12'b111111000111;
   51605: result <= 12'b111111000111;
   51606: result <= 12'b111111000111;
   51607: result <= 12'b111111000111;
   51608: result <= 12'b111111000111;
   51609: result <= 12'b111111000111;
   51610: result <= 12'b111111000111;
   51611: result <= 12'b111111000111;
   51612: result <= 12'b111111000111;
   51613: result <= 12'b111111000111;
   51614: result <= 12'b111111000111;
   51615: result <= 12'b111111000111;
   51616: result <= 12'b111111000111;
   51617: result <= 12'b111111000111;
   51618: result <= 12'b111111000111;
   51619: result <= 12'b111111000110;
   51620: result <= 12'b111111000110;
   51621: result <= 12'b111111000110;
   51622: result <= 12'b111111000110;
   51623: result <= 12'b111111000110;
   51624: result <= 12'b111111000110;
   51625: result <= 12'b111111000110;
   51626: result <= 12'b111111000110;
   51627: result <= 12'b111111000110;
   51628: result <= 12'b111111000110;
   51629: result <= 12'b111111000110;
   51630: result <= 12'b111111000110;
   51631: result <= 12'b111111000110;
   51632: result <= 12'b111111000110;
   51633: result <= 12'b111111000110;
   51634: result <= 12'b111111000110;
   51635: result <= 12'b111111000110;
   51636: result <= 12'b111111000110;
   51637: result <= 12'b111111000110;
   51638: result <= 12'b111111000110;
   51639: result <= 12'b111111000110;
   51640: result <= 12'b111111000110;
   51641: result <= 12'b111111000101;
   51642: result <= 12'b111111000101;
   51643: result <= 12'b111111000101;
   51644: result <= 12'b111111000101;
   51645: result <= 12'b111111000101;
   51646: result <= 12'b111111000101;
   51647: result <= 12'b111111000101;
   51648: result <= 12'b111111000101;
   51649: result <= 12'b111111000101;
   51650: result <= 12'b111111000101;
   51651: result <= 12'b111111000101;
   51652: result <= 12'b111111000101;
   51653: result <= 12'b111111000101;
   51654: result <= 12'b111111000101;
   51655: result <= 12'b111111000101;
   51656: result <= 12'b111111000101;
   51657: result <= 12'b111111000101;
   51658: result <= 12'b111111000101;
   51659: result <= 12'b111111000101;
   51660: result <= 12'b111111000101;
   51661: result <= 12'b111111000101;
   51662: result <= 12'b111111000100;
   51663: result <= 12'b111111000100;
   51664: result <= 12'b111111000100;
   51665: result <= 12'b111111000100;
   51666: result <= 12'b111111000100;
   51667: result <= 12'b111111000100;
   51668: result <= 12'b111111000100;
   51669: result <= 12'b111111000100;
   51670: result <= 12'b111111000100;
   51671: result <= 12'b111111000100;
   51672: result <= 12'b111111000100;
   51673: result <= 12'b111111000100;
   51674: result <= 12'b111111000100;
   51675: result <= 12'b111111000100;
   51676: result <= 12'b111111000100;
   51677: result <= 12'b111111000100;
   51678: result <= 12'b111111000100;
   51679: result <= 12'b111111000100;
   51680: result <= 12'b111111000100;
   51681: result <= 12'b111111000100;
   51682: result <= 12'b111111000100;
   51683: result <= 12'b111111000011;
   51684: result <= 12'b111111000011;
   51685: result <= 12'b111111000011;
   51686: result <= 12'b111111000011;
   51687: result <= 12'b111111000011;
   51688: result <= 12'b111111000011;
   51689: result <= 12'b111111000011;
   51690: result <= 12'b111111000011;
   51691: result <= 12'b111111000011;
   51692: result <= 12'b111111000011;
   51693: result <= 12'b111111000011;
   51694: result <= 12'b111111000011;
   51695: result <= 12'b111111000011;
   51696: result <= 12'b111111000011;
   51697: result <= 12'b111111000011;
   51698: result <= 12'b111111000011;
   51699: result <= 12'b111111000011;
   51700: result <= 12'b111111000011;
   51701: result <= 12'b111111000011;
   51702: result <= 12'b111111000011;
   51703: result <= 12'b111111000011;
   51704: result <= 12'b111111000011;
   51705: result <= 12'b111111000010;
   51706: result <= 12'b111111000010;
   51707: result <= 12'b111111000010;
   51708: result <= 12'b111111000010;
   51709: result <= 12'b111111000010;
   51710: result <= 12'b111111000010;
   51711: result <= 12'b111111000010;
   51712: result <= 12'b111111000010;
   51713: result <= 12'b111111000010;
   51714: result <= 12'b111111000010;
   51715: result <= 12'b111111000010;
   51716: result <= 12'b111111000010;
   51717: result <= 12'b111111000010;
   51718: result <= 12'b111111000010;
   51719: result <= 12'b111111000010;
   51720: result <= 12'b111111000010;
   51721: result <= 12'b111111000010;
   51722: result <= 12'b111111000010;
   51723: result <= 12'b111111000010;
   51724: result <= 12'b111111000010;
   51725: result <= 12'b111111000010;
   51726: result <= 12'b111111000001;
   51727: result <= 12'b111111000001;
   51728: result <= 12'b111111000001;
   51729: result <= 12'b111111000001;
   51730: result <= 12'b111111000001;
   51731: result <= 12'b111111000001;
   51732: result <= 12'b111111000001;
   51733: result <= 12'b111111000001;
   51734: result <= 12'b111111000001;
   51735: result <= 12'b111111000001;
   51736: result <= 12'b111111000001;
   51737: result <= 12'b111111000001;
   51738: result <= 12'b111111000001;
   51739: result <= 12'b111111000001;
   51740: result <= 12'b111111000001;
   51741: result <= 12'b111111000001;
   51742: result <= 12'b111111000001;
   51743: result <= 12'b111111000001;
   51744: result <= 12'b111111000001;
   51745: result <= 12'b111111000001;
   51746: result <= 12'b111111000000;
   51747: result <= 12'b111111000000;
   51748: result <= 12'b111111000000;
   51749: result <= 12'b111111000000;
   51750: result <= 12'b111111000000;
   51751: result <= 12'b111111000000;
   51752: result <= 12'b111111000000;
   51753: result <= 12'b111111000000;
   51754: result <= 12'b111111000000;
   51755: result <= 12'b111111000000;
   51756: result <= 12'b111111000000;
   51757: result <= 12'b111111000000;
   51758: result <= 12'b111111000000;
   51759: result <= 12'b111111000000;
   51760: result <= 12'b111111000000;
   51761: result <= 12'b111111000000;
   51762: result <= 12'b111111000000;
   51763: result <= 12'b111111000000;
   51764: result <= 12'b111111000000;
   51765: result <= 12'b111111000000;
   51766: result <= 12'b111111000000;
   51767: result <= 12'b111110111111;
   51768: result <= 12'b111110111111;
   51769: result <= 12'b111110111111;
   51770: result <= 12'b111110111111;
   51771: result <= 12'b111110111111;
   51772: result <= 12'b111110111111;
   51773: result <= 12'b111110111111;
   51774: result <= 12'b111110111111;
   51775: result <= 12'b111110111111;
   51776: result <= 12'b111110111111;
   51777: result <= 12'b111110111111;
   51778: result <= 12'b111110111111;
   51779: result <= 12'b111110111111;
   51780: result <= 12'b111110111111;
   51781: result <= 12'b111110111111;
   51782: result <= 12'b111110111111;
   51783: result <= 12'b111110111111;
   51784: result <= 12'b111110111111;
   51785: result <= 12'b111110111111;
   51786: result <= 12'b111110111111;
   51787: result <= 12'b111110111110;
   51788: result <= 12'b111110111110;
   51789: result <= 12'b111110111110;
   51790: result <= 12'b111110111110;
   51791: result <= 12'b111110111110;
   51792: result <= 12'b111110111110;
   51793: result <= 12'b111110111110;
   51794: result <= 12'b111110111110;
   51795: result <= 12'b111110111110;
   51796: result <= 12'b111110111110;
   51797: result <= 12'b111110111110;
   51798: result <= 12'b111110111110;
   51799: result <= 12'b111110111110;
   51800: result <= 12'b111110111110;
   51801: result <= 12'b111110111110;
   51802: result <= 12'b111110111110;
   51803: result <= 12'b111110111110;
   51804: result <= 12'b111110111110;
   51805: result <= 12'b111110111110;
   51806: result <= 12'b111110111110;
   51807: result <= 12'b111110111110;
   51808: result <= 12'b111110111101;
   51809: result <= 12'b111110111101;
   51810: result <= 12'b111110111101;
   51811: result <= 12'b111110111101;
   51812: result <= 12'b111110111101;
   51813: result <= 12'b111110111101;
   51814: result <= 12'b111110111101;
   51815: result <= 12'b111110111101;
   51816: result <= 12'b111110111101;
   51817: result <= 12'b111110111101;
   51818: result <= 12'b111110111101;
   51819: result <= 12'b111110111101;
   51820: result <= 12'b111110111101;
   51821: result <= 12'b111110111101;
   51822: result <= 12'b111110111101;
   51823: result <= 12'b111110111101;
   51824: result <= 12'b111110111101;
   51825: result <= 12'b111110111101;
   51826: result <= 12'b111110111101;
   51827: result <= 12'b111110111101;
   51828: result <= 12'b111110111100;
   51829: result <= 12'b111110111100;
   51830: result <= 12'b111110111100;
   51831: result <= 12'b111110111100;
   51832: result <= 12'b111110111100;
   51833: result <= 12'b111110111100;
   51834: result <= 12'b111110111100;
   51835: result <= 12'b111110111100;
   51836: result <= 12'b111110111100;
   51837: result <= 12'b111110111100;
   51838: result <= 12'b111110111100;
   51839: result <= 12'b111110111100;
   51840: result <= 12'b111110111100;
   51841: result <= 12'b111110111100;
   51842: result <= 12'b111110111100;
   51843: result <= 12'b111110111100;
   51844: result <= 12'b111110111100;
   51845: result <= 12'b111110111100;
   51846: result <= 12'b111110111100;
   51847: result <= 12'b111110111100;
   51848: result <= 12'b111110111011;
   51849: result <= 12'b111110111011;
   51850: result <= 12'b111110111011;
   51851: result <= 12'b111110111011;
   51852: result <= 12'b111110111011;
   51853: result <= 12'b111110111011;
   51854: result <= 12'b111110111011;
   51855: result <= 12'b111110111011;
   51856: result <= 12'b111110111011;
   51857: result <= 12'b111110111011;
   51858: result <= 12'b111110111011;
   51859: result <= 12'b111110111011;
   51860: result <= 12'b111110111011;
   51861: result <= 12'b111110111011;
   51862: result <= 12'b111110111011;
   51863: result <= 12'b111110111011;
   51864: result <= 12'b111110111011;
   51865: result <= 12'b111110111011;
   51866: result <= 12'b111110111011;
   51867: result <= 12'b111110111011;
   51868: result <= 12'b111110111010;
   51869: result <= 12'b111110111010;
   51870: result <= 12'b111110111010;
   51871: result <= 12'b111110111010;
   51872: result <= 12'b111110111010;
   51873: result <= 12'b111110111010;
   51874: result <= 12'b111110111010;
   51875: result <= 12'b111110111010;
   51876: result <= 12'b111110111010;
   51877: result <= 12'b111110111010;
   51878: result <= 12'b111110111010;
   51879: result <= 12'b111110111010;
   51880: result <= 12'b111110111010;
   51881: result <= 12'b111110111010;
   51882: result <= 12'b111110111010;
   51883: result <= 12'b111110111010;
   51884: result <= 12'b111110111010;
   51885: result <= 12'b111110111010;
   51886: result <= 12'b111110111010;
   51887: result <= 12'b111110111001;
   51888: result <= 12'b111110111001;
   51889: result <= 12'b111110111001;
   51890: result <= 12'b111110111001;
   51891: result <= 12'b111110111001;
   51892: result <= 12'b111110111001;
   51893: result <= 12'b111110111001;
   51894: result <= 12'b111110111001;
   51895: result <= 12'b111110111001;
   51896: result <= 12'b111110111001;
   51897: result <= 12'b111110111001;
   51898: result <= 12'b111110111001;
   51899: result <= 12'b111110111001;
   51900: result <= 12'b111110111001;
   51901: result <= 12'b111110111001;
   51902: result <= 12'b111110111001;
   51903: result <= 12'b111110111001;
   51904: result <= 12'b111110111001;
   51905: result <= 12'b111110111001;
   51906: result <= 12'b111110111001;
   51907: result <= 12'b111110111000;
   51908: result <= 12'b111110111000;
   51909: result <= 12'b111110111000;
   51910: result <= 12'b111110111000;
   51911: result <= 12'b111110111000;
   51912: result <= 12'b111110111000;
   51913: result <= 12'b111110111000;
   51914: result <= 12'b111110111000;
   51915: result <= 12'b111110111000;
   51916: result <= 12'b111110111000;
   51917: result <= 12'b111110111000;
   51918: result <= 12'b111110111000;
   51919: result <= 12'b111110111000;
   51920: result <= 12'b111110111000;
   51921: result <= 12'b111110111000;
   51922: result <= 12'b111110111000;
   51923: result <= 12'b111110111000;
   51924: result <= 12'b111110111000;
   51925: result <= 12'b111110111000;
   51926: result <= 12'b111110110111;
   51927: result <= 12'b111110110111;
   51928: result <= 12'b111110110111;
   51929: result <= 12'b111110110111;
   51930: result <= 12'b111110110111;
   51931: result <= 12'b111110110111;
   51932: result <= 12'b111110110111;
   51933: result <= 12'b111110110111;
   51934: result <= 12'b111110110111;
   51935: result <= 12'b111110110111;
   51936: result <= 12'b111110110111;
   51937: result <= 12'b111110110111;
   51938: result <= 12'b111110110111;
   51939: result <= 12'b111110110111;
   51940: result <= 12'b111110110111;
   51941: result <= 12'b111110110111;
   51942: result <= 12'b111110110111;
   51943: result <= 12'b111110110111;
   51944: result <= 12'b111110110111;
   51945: result <= 12'b111110110111;
   51946: result <= 12'b111110110110;
   51947: result <= 12'b111110110110;
   51948: result <= 12'b111110110110;
   51949: result <= 12'b111110110110;
   51950: result <= 12'b111110110110;
   51951: result <= 12'b111110110110;
   51952: result <= 12'b111110110110;
   51953: result <= 12'b111110110110;
   51954: result <= 12'b111110110110;
   51955: result <= 12'b111110110110;
   51956: result <= 12'b111110110110;
   51957: result <= 12'b111110110110;
   51958: result <= 12'b111110110110;
   51959: result <= 12'b111110110110;
   51960: result <= 12'b111110110110;
   51961: result <= 12'b111110110110;
   51962: result <= 12'b111110110110;
   51963: result <= 12'b111110110110;
   51964: result <= 12'b111110110110;
   51965: result <= 12'b111110110101;
   51966: result <= 12'b111110110101;
   51967: result <= 12'b111110110101;
   51968: result <= 12'b111110110101;
   51969: result <= 12'b111110110101;
   51970: result <= 12'b111110110101;
   51971: result <= 12'b111110110101;
   51972: result <= 12'b111110110101;
   51973: result <= 12'b111110110101;
   51974: result <= 12'b111110110101;
   51975: result <= 12'b111110110101;
   51976: result <= 12'b111110110101;
   51977: result <= 12'b111110110101;
   51978: result <= 12'b111110110101;
   51979: result <= 12'b111110110101;
   51980: result <= 12'b111110110101;
   51981: result <= 12'b111110110101;
   51982: result <= 12'b111110110101;
   51983: result <= 12'b111110110101;
   51984: result <= 12'b111110110100;
   51985: result <= 12'b111110110100;
   51986: result <= 12'b111110110100;
   51987: result <= 12'b111110110100;
   51988: result <= 12'b111110110100;
   51989: result <= 12'b111110110100;
   51990: result <= 12'b111110110100;
   51991: result <= 12'b111110110100;
   51992: result <= 12'b111110110100;
   51993: result <= 12'b111110110100;
   51994: result <= 12'b111110110100;
   51995: result <= 12'b111110110100;
   51996: result <= 12'b111110110100;
   51997: result <= 12'b111110110100;
   51998: result <= 12'b111110110100;
   51999: result <= 12'b111110110100;
   52000: result <= 12'b111110110100;
   52001: result <= 12'b111110110100;
   52002: result <= 12'b111110110100;
   52003: result <= 12'b111110110011;
   52004: result <= 12'b111110110011;
   52005: result <= 12'b111110110011;
   52006: result <= 12'b111110110011;
   52007: result <= 12'b111110110011;
   52008: result <= 12'b111110110011;
   52009: result <= 12'b111110110011;
   52010: result <= 12'b111110110011;
   52011: result <= 12'b111110110011;
   52012: result <= 12'b111110110011;
   52013: result <= 12'b111110110011;
   52014: result <= 12'b111110110011;
   52015: result <= 12'b111110110011;
   52016: result <= 12'b111110110011;
   52017: result <= 12'b111110110011;
   52018: result <= 12'b111110110011;
   52019: result <= 12'b111110110011;
   52020: result <= 12'b111110110011;
   52021: result <= 12'b111110110011;
   52022: result <= 12'b111110110010;
   52023: result <= 12'b111110110010;
   52024: result <= 12'b111110110010;
   52025: result <= 12'b111110110010;
   52026: result <= 12'b111110110010;
   52027: result <= 12'b111110110010;
   52028: result <= 12'b111110110010;
   52029: result <= 12'b111110110010;
   52030: result <= 12'b111110110010;
   52031: result <= 12'b111110110010;
   52032: result <= 12'b111110110010;
   52033: result <= 12'b111110110010;
   52034: result <= 12'b111110110010;
   52035: result <= 12'b111110110010;
   52036: result <= 12'b111110110010;
   52037: result <= 12'b111110110010;
   52038: result <= 12'b111110110010;
   52039: result <= 12'b111110110010;
   52040: result <= 12'b111110110001;
   52041: result <= 12'b111110110001;
   52042: result <= 12'b111110110001;
   52043: result <= 12'b111110110001;
   52044: result <= 12'b111110110001;
   52045: result <= 12'b111110110001;
   52046: result <= 12'b111110110001;
   52047: result <= 12'b111110110001;
   52048: result <= 12'b111110110001;
   52049: result <= 12'b111110110001;
   52050: result <= 12'b111110110001;
   52051: result <= 12'b111110110001;
   52052: result <= 12'b111110110001;
   52053: result <= 12'b111110110001;
   52054: result <= 12'b111110110001;
   52055: result <= 12'b111110110001;
   52056: result <= 12'b111110110001;
   52057: result <= 12'b111110110001;
   52058: result <= 12'b111110110001;
   52059: result <= 12'b111110110000;
   52060: result <= 12'b111110110000;
   52061: result <= 12'b111110110000;
   52062: result <= 12'b111110110000;
   52063: result <= 12'b111110110000;
   52064: result <= 12'b111110110000;
   52065: result <= 12'b111110110000;
   52066: result <= 12'b111110110000;
   52067: result <= 12'b111110110000;
   52068: result <= 12'b111110110000;
   52069: result <= 12'b111110110000;
   52070: result <= 12'b111110110000;
   52071: result <= 12'b111110110000;
   52072: result <= 12'b111110110000;
   52073: result <= 12'b111110110000;
   52074: result <= 12'b111110110000;
   52075: result <= 12'b111110110000;
   52076: result <= 12'b111110110000;
   52077: result <= 12'b111110101111;
   52078: result <= 12'b111110101111;
   52079: result <= 12'b111110101111;
   52080: result <= 12'b111110101111;
   52081: result <= 12'b111110101111;
   52082: result <= 12'b111110101111;
   52083: result <= 12'b111110101111;
   52084: result <= 12'b111110101111;
   52085: result <= 12'b111110101111;
   52086: result <= 12'b111110101111;
   52087: result <= 12'b111110101111;
   52088: result <= 12'b111110101111;
   52089: result <= 12'b111110101111;
   52090: result <= 12'b111110101111;
   52091: result <= 12'b111110101111;
   52092: result <= 12'b111110101111;
   52093: result <= 12'b111110101111;
   52094: result <= 12'b111110101111;
   52095: result <= 12'b111110101111;
   52096: result <= 12'b111110101110;
   52097: result <= 12'b111110101110;
   52098: result <= 12'b111110101110;
   52099: result <= 12'b111110101110;
   52100: result <= 12'b111110101110;
   52101: result <= 12'b111110101110;
   52102: result <= 12'b111110101110;
   52103: result <= 12'b111110101110;
   52104: result <= 12'b111110101110;
   52105: result <= 12'b111110101110;
   52106: result <= 12'b111110101110;
   52107: result <= 12'b111110101110;
   52108: result <= 12'b111110101110;
   52109: result <= 12'b111110101110;
   52110: result <= 12'b111110101110;
   52111: result <= 12'b111110101110;
   52112: result <= 12'b111110101110;
   52113: result <= 12'b111110101110;
   52114: result <= 12'b111110101101;
   52115: result <= 12'b111110101101;
   52116: result <= 12'b111110101101;
   52117: result <= 12'b111110101101;
   52118: result <= 12'b111110101101;
   52119: result <= 12'b111110101101;
   52120: result <= 12'b111110101101;
   52121: result <= 12'b111110101101;
   52122: result <= 12'b111110101101;
   52123: result <= 12'b111110101101;
   52124: result <= 12'b111110101101;
   52125: result <= 12'b111110101101;
   52126: result <= 12'b111110101101;
   52127: result <= 12'b111110101101;
   52128: result <= 12'b111110101101;
   52129: result <= 12'b111110101101;
   52130: result <= 12'b111110101101;
   52131: result <= 12'b111110101101;
   52132: result <= 12'b111110101100;
   52133: result <= 12'b111110101100;
   52134: result <= 12'b111110101100;
   52135: result <= 12'b111110101100;
   52136: result <= 12'b111110101100;
   52137: result <= 12'b111110101100;
   52138: result <= 12'b111110101100;
   52139: result <= 12'b111110101100;
   52140: result <= 12'b111110101100;
   52141: result <= 12'b111110101100;
   52142: result <= 12'b111110101100;
   52143: result <= 12'b111110101100;
   52144: result <= 12'b111110101100;
   52145: result <= 12'b111110101100;
   52146: result <= 12'b111110101100;
   52147: result <= 12'b111110101100;
   52148: result <= 12'b111110101100;
   52149: result <= 12'b111110101100;
   52150: result <= 12'b111110101011;
   52151: result <= 12'b111110101011;
   52152: result <= 12'b111110101011;
   52153: result <= 12'b111110101011;
   52154: result <= 12'b111110101011;
   52155: result <= 12'b111110101011;
   52156: result <= 12'b111110101011;
   52157: result <= 12'b111110101011;
   52158: result <= 12'b111110101011;
   52159: result <= 12'b111110101011;
   52160: result <= 12'b111110101011;
   52161: result <= 12'b111110101011;
   52162: result <= 12'b111110101011;
   52163: result <= 12'b111110101011;
   52164: result <= 12'b111110101011;
   52165: result <= 12'b111110101011;
   52166: result <= 12'b111110101011;
   52167: result <= 12'b111110101011;
   52168: result <= 12'b111110101010;
   52169: result <= 12'b111110101010;
   52170: result <= 12'b111110101010;
   52171: result <= 12'b111110101010;
   52172: result <= 12'b111110101010;
   52173: result <= 12'b111110101010;
   52174: result <= 12'b111110101010;
   52175: result <= 12'b111110101010;
   52176: result <= 12'b111110101010;
   52177: result <= 12'b111110101010;
   52178: result <= 12'b111110101010;
   52179: result <= 12'b111110101010;
   52180: result <= 12'b111110101010;
   52181: result <= 12'b111110101010;
   52182: result <= 12'b111110101010;
   52183: result <= 12'b111110101010;
   52184: result <= 12'b111110101010;
   52185: result <= 12'b111110101010;
   52186: result <= 12'b111110101001;
   52187: result <= 12'b111110101001;
   52188: result <= 12'b111110101001;
   52189: result <= 12'b111110101001;
   52190: result <= 12'b111110101001;
   52191: result <= 12'b111110101001;
   52192: result <= 12'b111110101001;
   52193: result <= 12'b111110101001;
   52194: result <= 12'b111110101001;
   52195: result <= 12'b111110101001;
   52196: result <= 12'b111110101001;
   52197: result <= 12'b111110101001;
   52198: result <= 12'b111110101001;
   52199: result <= 12'b111110101001;
   52200: result <= 12'b111110101001;
   52201: result <= 12'b111110101001;
   52202: result <= 12'b111110101001;
   52203: result <= 12'b111110101001;
   52204: result <= 12'b111110101000;
   52205: result <= 12'b111110101000;
   52206: result <= 12'b111110101000;
   52207: result <= 12'b111110101000;
   52208: result <= 12'b111110101000;
   52209: result <= 12'b111110101000;
   52210: result <= 12'b111110101000;
   52211: result <= 12'b111110101000;
   52212: result <= 12'b111110101000;
   52213: result <= 12'b111110101000;
   52214: result <= 12'b111110101000;
   52215: result <= 12'b111110101000;
   52216: result <= 12'b111110101000;
   52217: result <= 12'b111110101000;
   52218: result <= 12'b111110101000;
   52219: result <= 12'b111110101000;
   52220: result <= 12'b111110101000;
   52221: result <= 12'b111110100111;
   52222: result <= 12'b111110100111;
   52223: result <= 12'b111110100111;
   52224: result <= 12'b111110100111;
   52225: result <= 12'b111110100111;
   52226: result <= 12'b111110100111;
   52227: result <= 12'b111110100111;
   52228: result <= 12'b111110100111;
   52229: result <= 12'b111110100111;
   52230: result <= 12'b111110100111;
   52231: result <= 12'b111110100111;
   52232: result <= 12'b111110100111;
   52233: result <= 12'b111110100111;
   52234: result <= 12'b111110100111;
   52235: result <= 12'b111110100111;
   52236: result <= 12'b111110100111;
   52237: result <= 12'b111110100111;
   52238: result <= 12'b111110100111;
   52239: result <= 12'b111110100110;
   52240: result <= 12'b111110100110;
   52241: result <= 12'b111110100110;
   52242: result <= 12'b111110100110;
   52243: result <= 12'b111110100110;
   52244: result <= 12'b111110100110;
   52245: result <= 12'b111110100110;
   52246: result <= 12'b111110100110;
   52247: result <= 12'b111110100110;
   52248: result <= 12'b111110100110;
   52249: result <= 12'b111110100110;
   52250: result <= 12'b111110100110;
   52251: result <= 12'b111110100110;
   52252: result <= 12'b111110100110;
   52253: result <= 12'b111110100110;
   52254: result <= 12'b111110100110;
   52255: result <= 12'b111110100110;
   52256: result <= 12'b111110100101;
   52257: result <= 12'b111110100101;
   52258: result <= 12'b111110100101;
   52259: result <= 12'b111110100101;
   52260: result <= 12'b111110100101;
   52261: result <= 12'b111110100101;
   52262: result <= 12'b111110100101;
   52263: result <= 12'b111110100101;
   52264: result <= 12'b111110100101;
   52265: result <= 12'b111110100101;
   52266: result <= 12'b111110100101;
   52267: result <= 12'b111110100101;
   52268: result <= 12'b111110100101;
   52269: result <= 12'b111110100101;
   52270: result <= 12'b111110100101;
   52271: result <= 12'b111110100101;
   52272: result <= 12'b111110100101;
   52273: result <= 12'b111110100100;
   52274: result <= 12'b111110100100;
   52275: result <= 12'b111110100100;
   52276: result <= 12'b111110100100;
   52277: result <= 12'b111110100100;
   52278: result <= 12'b111110100100;
   52279: result <= 12'b111110100100;
   52280: result <= 12'b111110100100;
   52281: result <= 12'b111110100100;
   52282: result <= 12'b111110100100;
   52283: result <= 12'b111110100100;
   52284: result <= 12'b111110100100;
   52285: result <= 12'b111110100100;
   52286: result <= 12'b111110100100;
   52287: result <= 12'b111110100100;
   52288: result <= 12'b111110100100;
   52289: result <= 12'b111110100100;
   52290: result <= 12'b111110100100;
   52291: result <= 12'b111110100011;
   52292: result <= 12'b111110100011;
   52293: result <= 12'b111110100011;
   52294: result <= 12'b111110100011;
   52295: result <= 12'b111110100011;
   52296: result <= 12'b111110100011;
   52297: result <= 12'b111110100011;
   52298: result <= 12'b111110100011;
   52299: result <= 12'b111110100011;
   52300: result <= 12'b111110100011;
   52301: result <= 12'b111110100011;
   52302: result <= 12'b111110100011;
   52303: result <= 12'b111110100011;
   52304: result <= 12'b111110100011;
   52305: result <= 12'b111110100011;
   52306: result <= 12'b111110100011;
   52307: result <= 12'b111110100011;
   52308: result <= 12'b111110100010;
   52309: result <= 12'b111110100010;
   52310: result <= 12'b111110100010;
   52311: result <= 12'b111110100010;
   52312: result <= 12'b111110100010;
   52313: result <= 12'b111110100010;
   52314: result <= 12'b111110100010;
   52315: result <= 12'b111110100010;
   52316: result <= 12'b111110100010;
   52317: result <= 12'b111110100010;
   52318: result <= 12'b111110100010;
   52319: result <= 12'b111110100010;
   52320: result <= 12'b111110100010;
   52321: result <= 12'b111110100010;
   52322: result <= 12'b111110100010;
   52323: result <= 12'b111110100010;
   52324: result <= 12'b111110100010;
   52325: result <= 12'b111110100001;
   52326: result <= 12'b111110100001;
   52327: result <= 12'b111110100001;
   52328: result <= 12'b111110100001;
   52329: result <= 12'b111110100001;
   52330: result <= 12'b111110100001;
   52331: result <= 12'b111110100001;
   52332: result <= 12'b111110100001;
   52333: result <= 12'b111110100001;
   52334: result <= 12'b111110100001;
   52335: result <= 12'b111110100001;
   52336: result <= 12'b111110100001;
   52337: result <= 12'b111110100001;
   52338: result <= 12'b111110100001;
   52339: result <= 12'b111110100001;
   52340: result <= 12'b111110100001;
   52341: result <= 12'b111110100001;
   52342: result <= 12'b111110100000;
   52343: result <= 12'b111110100000;
   52344: result <= 12'b111110100000;
   52345: result <= 12'b111110100000;
   52346: result <= 12'b111110100000;
   52347: result <= 12'b111110100000;
   52348: result <= 12'b111110100000;
   52349: result <= 12'b111110100000;
   52350: result <= 12'b111110100000;
   52351: result <= 12'b111110100000;
   52352: result <= 12'b111110100000;
   52353: result <= 12'b111110100000;
   52354: result <= 12'b111110100000;
   52355: result <= 12'b111110100000;
   52356: result <= 12'b111110100000;
   52357: result <= 12'b111110100000;
   52358: result <= 12'b111110100000;
   52359: result <= 12'b111110011111;
   52360: result <= 12'b111110011111;
   52361: result <= 12'b111110011111;
   52362: result <= 12'b111110011111;
   52363: result <= 12'b111110011111;
   52364: result <= 12'b111110011111;
   52365: result <= 12'b111110011111;
   52366: result <= 12'b111110011111;
   52367: result <= 12'b111110011111;
   52368: result <= 12'b111110011111;
   52369: result <= 12'b111110011111;
   52370: result <= 12'b111110011111;
   52371: result <= 12'b111110011111;
   52372: result <= 12'b111110011111;
   52373: result <= 12'b111110011111;
   52374: result <= 12'b111110011111;
   52375: result <= 12'b111110011111;
   52376: result <= 12'b111110011110;
   52377: result <= 12'b111110011110;
   52378: result <= 12'b111110011110;
   52379: result <= 12'b111110011110;
   52380: result <= 12'b111110011110;
   52381: result <= 12'b111110011110;
   52382: result <= 12'b111110011110;
   52383: result <= 12'b111110011110;
   52384: result <= 12'b111110011110;
   52385: result <= 12'b111110011110;
   52386: result <= 12'b111110011110;
   52387: result <= 12'b111110011110;
   52388: result <= 12'b111110011110;
   52389: result <= 12'b111110011110;
   52390: result <= 12'b111110011110;
   52391: result <= 12'b111110011110;
   52392: result <= 12'b111110011101;
   52393: result <= 12'b111110011101;
   52394: result <= 12'b111110011101;
   52395: result <= 12'b111110011101;
   52396: result <= 12'b111110011101;
   52397: result <= 12'b111110011101;
   52398: result <= 12'b111110011101;
   52399: result <= 12'b111110011101;
   52400: result <= 12'b111110011101;
   52401: result <= 12'b111110011101;
   52402: result <= 12'b111110011101;
   52403: result <= 12'b111110011101;
   52404: result <= 12'b111110011101;
   52405: result <= 12'b111110011101;
   52406: result <= 12'b111110011101;
   52407: result <= 12'b111110011101;
   52408: result <= 12'b111110011101;
   52409: result <= 12'b111110011100;
   52410: result <= 12'b111110011100;
   52411: result <= 12'b111110011100;
   52412: result <= 12'b111110011100;
   52413: result <= 12'b111110011100;
   52414: result <= 12'b111110011100;
   52415: result <= 12'b111110011100;
   52416: result <= 12'b111110011100;
   52417: result <= 12'b111110011100;
   52418: result <= 12'b111110011100;
   52419: result <= 12'b111110011100;
   52420: result <= 12'b111110011100;
   52421: result <= 12'b111110011100;
   52422: result <= 12'b111110011100;
   52423: result <= 12'b111110011100;
   52424: result <= 12'b111110011100;
   52425: result <= 12'b111110011011;
   52426: result <= 12'b111110011011;
   52427: result <= 12'b111110011011;
   52428: result <= 12'b111110011011;
   52429: result <= 12'b111110011011;
   52430: result <= 12'b111110011011;
   52431: result <= 12'b111110011011;
   52432: result <= 12'b111110011011;
   52433: result <= 12'b111110011011;
   52434: result <= 12'b111110011011;
   52435: result <= 12'b111110011011;
   52436: result <= 12'b111110011011;
   52437: result <= 12'b111110011011;
   52438: result <= 12'b111110011011;
   52439: result <= 12'b111110011011;
   52440: result <= 12'b111110011011;
   52441: result <= 12'b111110011011;
   52442: result <= 12'b111110011010;
   52443: result <= 12'b111110011010;
   52444: result <= 12'b111110011010;
   52445: result <= 12'b111110011010;
   52446: result <= 12'b111110011010;
   52447: result <= 12'b111110011010;
   52448: result <= 12'b111110011010;
   52449: result <= 12'b111110011010;
   52450: result <= 12'b111110011010;
   52451: result <= 12'b111110011010;
   52452: result <= 12'b111110011010;
   52453: result <= 12'b111110011010;
   52454: result <= 12'b111110011010;
   52455: result <= 12'b111110011010;
   52456: result <= 12'b111110011010;
   52457: result <= 12'b111110011010;
   52458: result <= 12'b111110011001;
   52459: result <= 12'b111110011001;
   52460: result <= 12'b111110011001;
   52461: result <= 12'b111110011001;
   52462: result <= 12'b111110011001;
   52463: result <= 12'b111110011001;
   52464: result <= 12'b111110011001;
   52465: result <= 12'b111110011001;
   52466: result <= 12'b111110011001;
   52467: result <= 12'b111110011001;
   52468: result <= 12'b111110011001;
   52469: result <= 12'b111110011001;
   52470: result <= 12'b111110011001;
   52471: result <= 12'b111110011001;
   52472: result <= 12'b111110011001;
   52473: result <= 12'b111110011001;
   52474: result <= 12'b111110011001;
   52475: result <= 12'b111110011000;
   52476: result <= 12'b111110011000;
   52477: result <= 12'b111110011000;
   52478: result <= 12'b111110011000;
   52479: result <= 12'b111110011000;
   52480: result <= 12'b111110011000;
   52481: result <= 12'b111110011000;
   52482: result <= 12'b111110011000;
   52483: result <= 12'b111110011000;
   52484: result <= 12'b111110011000;
   52485: result <= 12'b111110011000;
   52486: result <= 12'b111110011000;
   52487: result <= 12'b111110011000;
   52488: result <= 12'b111110011000;
   52489: result <= 12'b111110011000;
   52490: result <= 12'b111110011000;
   52491: result <= 12'b111110010111;
   52492: result <= 12'b111110010111;
   52493: result <= 12'b111110010111;
   52494: result <= 12'b111110010111;
   52495: result <= 12'b111110010111;
   52496: result <= 12'b111110010111;
   52497: result <= 12'b111110010111;
   52498: result <= 12'b111110010111;
   52499: result <= 12'b111110010111;
   52500: result <= 12'b111110010111;
   52501: result <= 12'b111110010111;
   52502: result <= 12'b111110010111;
   52503: result <= 12'b111110010111;
   52504: result <= 12'b111110010111;
   52505: result <= 12'b111110010111;
   52506: result <= 12'b111110010111;
   52507: result <= 12'b111110010110;
   52508: result <= 12'b111110010110;
   52509: result <= 12'b111110010110;
   52510: result <= 12'b111110010110;
   52511: result <= 12'b111110010110;
   52512: result <= 12'b111110010110;
   52513: result <= 12'b111110010110;
   52514: result <= 12'b111110010110;
   52515: result <= 12'b111110010110;
   52516: result <= 12'b111110010110;
   52517: result <= 12'b111110010110;
   52518: result <= 12'b111110010110;
   52519: result <= 12'b111110010110;
   52520: result <= 12'b111110010110;
   52521: result <= 12'b111110010110;
   52522: result <= 12'b111110010110;
   52523: result <= 12'b111110010101;
   52524: result <= 12'b111110010101;
   52525: result <= 12'b111110010101;
   52526: result <= 12'b111110010101;
   52527: result <= 12'b111110010101;
   52528: result <= 12'b111110010101;
   52529: result <= 12'b111110010101;
   52530: result <= 12'b111110010101;
   52531: result <= 12'b111110010101;
   52532: result <= 12'b111110010101;
   52533: result <= 12'b111110010101;
   52534: result <= 12'b111110010101;
   52535: result <= 12'b111110010101;
   52536: result <= 12'b111110010101;
   52537: result <= 12'b111110010101;
   52538: result <= 12'b111110010101;
   52539: result <= 12'b111110010100;
   52540: result <= 12'b111110010100;
   52541: result <= 12'b111110010100;
   52542: result <= 12'b111110010100;
   52543: result <= 12'b111110010100;
   52544: result <= 12'b111110010100;
   52545: result <= 12'b111110010100;
   52546: result <= 12'b111110010100;
   52547: result <= 12'b111110010100;
   52548: result <= 12'b111110010100;
   52549: result <= 12'b111110010100;
   52550: result <= 12'b111110010100;
   52551: result <= 12'b111110010100;
   52552: result <= 12'b111110010100;
   52553: result <= 12'b111110010100;
   52554: result <= 12'b111110010100;
   52555: result <= 12'b111110010011;
   52556: result <= 12'b111110010011;
   52557: result <= 12'b111110010011;
   52558: result <= 12'b111110010011;
   52559: result <= 12'b111110010011;
   52560: result <= 12'b111110010011;
   52561: result <= 12'b111110010011;
   52562: result <= 12'b111110010011;
   52563: result <= 12'b111110010011;
   52564: result <= 12'b111110010011;
   52565: result <= 12'b111110010011;
   52566: result <= 12'b111110010011;
   52567: result <= 12'b111110010011;
   52568: result <= 12'b111110010011;
   52569: result <= 12'b111110010011;
   52570: result <= 12'b111110010011;
   52571: result <= 12'b111110010010;
   52572: result <= 12'b111110010010;
   52573: result <= 12'b111110010010;
   52574: result <= 12'b111110010010;
   52575: result <= 12'b111110010010;
   52576: result <= 12'b111110010010;
   52577: result <= 12'b111110010010;
   52578: result <= 12'b111110010010;
   52579: result <= 12'b111110010010;
   52580: result <= 12'b111110010010;
   52581: result <= 12'b111110010010;
   52582: result <= 12'b111110010010;
   52583: result <= 12'b111110010010;
   52584: result <= 12'b111110010010;
   52585: result <= 12'b111110010010;
   52586: result <= 12'b111110010010;
   52587: result <= 12'b111110010001;
   52588: result <= 12'b111110010001;
   52589: result <= 12'b111110010001;
   52590: result <= 12'b111110010001;
   52591: result <= 12'b111110010001;
   52592: result <= 12'b111110010001;
   52593: result <= 12'b111110010001;
   52594: result <= 12'b111110010001;
   52595: result <= 12'b111110010001;
   52596: result <= 12'b111110010001;
   52597: result <= 12'b111110010001;
   52598: result <= 12'b111110010001;
   52599: result <= 12'b111110010001;
   52600: result <= 12'b111110010001;
   52601: result <= 12'b111110010001;
   52602: result <= 12'b111110010000;
   52603: result <= 12'b111110010000;
   52604: result <= 12'b111110010000;
   52605: result <= 12'b111110010000;
   52606: result <= 12'b111110010000;
   52607: result <= 12'b111110010000;
   52608: result <= 12'b111110010000;
   52609: result <= 12'b111110010000;
   52610: result <= 12'b111110010000;
   52611: result <= 12'b111110010000;
   52612: result <= 12'b111110010000;
   52613: result <= 12'b111110010000;
   52614: result <= 12'b111110010000;
   52615: result <= 12'b111110010000;
   52616: result <= 12'b111110010000;
   52617: result <= 12'b111110010000;
   52618: result <= 12'b111110001111;
   52619: result <= 12'b111110001111;
   52620: result <= 12'b111110001111;
   52621: result <= 12'b111110001111;
   52622: result <= 12'b111110001111;
   52623: result <= 12'b111110001111;
   52624: result <= 12'b111110001111;
   52625: result <= 12'b111110001111;
   52626: result <= 12'b111110001111;
   52627: result <= 12'b111110001111;
   52628: result <= 12'b111110001111;
   52629: result <= 12'b111110001111;
   52630: result <= 12'b111110001111;
   52631: result <= 12'b111110001111;
   52632: result <= 12'b111110001111;
   52633: result <= 12'b111110001111;
   52634: result <= 12'b111110001110;
   52635: result <= 12'b111110001110;
   52636: result <= 12'b111110001110;
   52637: result <= 12'b111110001110;
   52638: result <= 12'b111110001110;
   52639: result <= 12'b111110001110;
   52640: result <= 12'b111110001110;
   52641: result <= 12'b111110001110;
   52642: result <= 12'b111110001110;
   52643: result <= 12'b111110001110;
   52644: result <= 12'b111110001110;
   52645: result <= 12'b111110001110;
   52646: result <= 12'b111110001110;
   52647: result <= 12'b111110001110;
   52648: result <= 12'b111110001110;
   52649: result <= 12'b111110001101;
   52650: result <= 12'b111110001101;
   52651: result <= 12'b111110001101;
   52652: result <= 12'b111110001101;
   52653: result <= 12'b111110001101;
   52654: result <= 12'b111110001101;
   52655: result <= 12'b111110001101;
   52656: result <= 12'b111110001101;
   52657: result <= 12'b111110001101;
   52658: result <= 12'b111110001101;
   52659: result <= 12'b111110001101;
   52660: result <= 12'b111110001101;
   52661: result <= 12'b111110001101;
   52662: result <= 12'b111110001101;
   52663: result <= 12'b111110001101;
   52664: result <= 12'b111110001100;
   52665: result <= 12'b111110001100;
   52666: result <= 12'b111110001100;
   52667: result <= 12'b111110001100;
   52668: result <= 12'b111110001100;
   52669: result <= 12'b111110001100;
   52670: result <= 12'b111110001100;
   52671: result <= 12'b111110001100;
   52672: result <= 12'b111110001100;
   52673: result <= 12'b111110001100;
   52674: result <= 12'b111110001100;
   52675: result <= 12'b111110001100;
   52676: result <= 12'b111110001100;
   52677: result <= 12'b111110001100;
   52678: result <= 12'b111110001100;
   52679: result <= 12'b111110001100;
   52680: result <= 12'b111110001011;
   52681: result <= 12'b111110001011;
   52682: result <= 12'b111110001011;
   52683: result <= 12'b111110001011;
   52684: result <= 12'b111110001011;
   52685: result <= 12'b111110001011;
   52686: result <= 12'b111110001011;
   52687: result <= 12'b111110001011;
   52688: result <= 12'b111110001011;
   52689: result <= 12'b111110001011;
   52690: result <= 12'b111110001011;
   52691: result <= 12'b111110001011;
   52692: result <= 12'b111110001011;
   52693: result <= 12'b111110001011;
   52694: result <= 12'b111110001011;
   52695: result <= 12'b111110001010;
   52696: result <= 12'b111110001010;
   52697: result <= 12'b111110001010;
   52698: result <= 12'b111110001010;
   52699: result <= 12'b111110001010;
   52700: result <= 12'b111110001010;
   52701: result <= 12'b111110001010;
   52702: result <= 12'b111110001010;
   52703: result <= 12'b111110001010;
   52704: result <= 12'b111110001010;
   52705: result <= 12'b111110001010;
   52706: result <= 12'b111110001010;
   52707: result <= 12'b111110001010;
   52708: result <= 12'b111110001010;
   52709: result <= 12'b111110001010;
   52710: result <= 12'b111110001001;
   52711: result <= 12'b111110001001;
   52712: result <= 12'b111110001001;
   52713: result <= 12'b111110001001;
   52714: result <= 12'b111110001001;
   52715: result <= 12'b111110001001;
   52716: result <= 12'b111110001001;
   52717: result <= 12'b111110001001;
   52718: result <= 12'b111110001001;
   52719: result <= 12'b111110001001;
   52720: result <= 12'b111110001001;
   52721: result <= 12'b111110001001;
   52722: result <= 12'b111110001001;
   52723: result <= 12'b111110001001;
   52724: result <= 12'b111110001001;
   52725: result <= 12'b111110001001;
   52726: result <= 12'b111110001000;
   52727: result <= 12'b111110001000;
   52728: result <= 12'b111110001000;
   52729: result <= 12'b111110001000;
   52730: result <= 12'b111110001000;
   52731: result <= 12'b111110001000;
   52732: result <= 12'b111110001000;
   52733: result <= 12'b111110001000;
   52734: result <= 12'b111110001000;
   52735: result <= 12'b111110001000;
   52736: result <= 12'b111110001000;
   52737: result <= 12'b111110001000;
   52738: result <= 12'b111110001000;
   52739: result <= 12'b111110001000;
   52740: result <= 12'b111110001000;
   52741: result <= 12'b111110000111;
   52742: result <= 12'b111110000111;
   52743: result <= 12'b111110000111;
   52744: result <= 12'b111110000111;
   52745: result <= 12'b111110000111;
   52746: result <= 12'b111110000111;
   52747: result <= 12'b111110000111;
   52748: result <= 12'b111110000111;
   52749: result <= 12'b111110000111;
   52750: result <= 12'b111110000111;
   52751: result <= 12'b111110000111;
   52752: result <= 12'b111110000111;
   52753: result <= 12'b111110000111;
   52754: result <= 12'b111110000111;
   52755: result <= 12'b111110000111;
   52756: result <= 12'b111110000110;
   52757: result <= 12'b111110000110;
   52758: result <= 12'b111110000110;
   52759: result <= 12'b111110000110;
   52760: result <= 12'b111110000110;
   52761: result <= 12'b111110000110;
   52762: result <= 12'b111110000110;
   52763: result <= 12'b111110000110;
   52764: result <= 12'b111110000110;
   52765: result <= 12'b111110000110;
   52766: result <= 12'b111110000110;
   52767: result <= 12'b111110000110;
   52768: result <= 12'b111110000110;
   52769: result <= 12'b111110000110;
   52770: result <= 12'b111110000110;
   52771: result <= 12'b111110000101;
   52772: result <= 12'b111110000101;
   52773: result <= 12'b111110000101;
   52774: result <= 12'b111110000101;
   52775: result <= 12'b111110000101;
   52776: result <= 12'b111110000101;
   52777: result <= 12'b111110000101;
   52778: result <= 12'b111110000101;
   52779: result <= 12'b111110000101;
   52780: result <= 12'b111110000101;
   52781: result <= 12'b111110000101;
   52782: result <= 12'b111110000101;
   52783: result <= 12'b111110000101;
   52784: result <= 12'b111110000101;
   52785: result <= 12'b111110000101;
   52786: result <= 12'b111110000100;
   52787: result <= 12'b111110000100;
   52788: result <= 12'b111110000100;
   52789: result <= 12'b111110000100;
   52790: result <= 12'b111110000100;
   52791: result <= 12'b111110000100;
   52792: result <= 12'b111110000100;
   52793: result <= 12'b111110000100;
   52794: result <= 12'b111110000100;
   52795: result <= 12'b111110000100;
   52796: result <= 12'b111110000100;
   52797: result <= 12'b111110000100;
   52798: result <= 12'b111110000100;
   52799: result <= 12'b111110000100;
   52800: result <= 12'b111110000100;
   52801: result <= 12'b111110000011;
   52802: result <= 12'b111110000011;
   52803: result <= 12'b111110000011;
   52804: result <= 12'b111110000011;
   52805: result <= 12'b111110000011;
   52806: result <= 12'b111110000011;
   52807: result <= 12'b111110000011;
   52808: result <= 12'b111110000011;
   52809: result <= 12'b111110000011;
   52810: result <= 12'b111110000011;
   52811: result <= 12'b111110000011;
   52812: result <= 12'b111110000011;
   52813: result <= 12'b111110000011;
   52814: result <= 12'b111110000011;
   52815: result <= 12'b111110000011;
   52816: result <= 12'b111110000010;
   52817: result <= 12'b111110000010;
   52818: result <= 12'b111110000010;
   52819: result <= 12'b111110000010;
   52820: result <= 12'b111110000010;
   52821: result <= 12'b111110000010;
   52822: result <= 12'b111110000010;
   52823: result <= 12'b111110000010;
   52824: result <= 12'b111110000010;
   52825: result <= 12'b111110000010;
   52826: result <= 12'b111110000010;
   52827: result <= 12'b111110000010;
   52828: result <= 12'b111110000010;
   52829: result <= 12'b111110000010;
   52830: result <= 12'b111110000001;
   52831: result <= 12'b111110000001;
   52832: result <= 12'b111110000001;
   52833: result <= 12'b111110000001;
   52834: result <= 12'b111110000001;
   52835: result <= 12'b111110000001;
   52836: result <= 12'b111110000001;
   52837: result <= 12'b111110000001;
   52838: result <= 12'b111110000001;
   52839: result <= 12'b111110000001;
   52840: result <= 12'b111110000001;
   52841: result <= 12'b111110000001;
   52842: result <= 12'b111110000001;
   52843: result <= 12'b111110000001;
   52844: result <= 12'b111110000001;
   52845: result <= 12'b111110000000;
   52846: result <= 12'b111110000000;
   52847: result <= 12'b111110000000;
   52848: result <= 12'b111110000000;
   52849: result <= 12'b111110000000;
   52850: result <= 12'b111110000000;
   52851: result <= 12'b111110000000;
   52852: result <= 12'b111110000000;
   52853: result <= 12'b111110000000;
   52854: result <= 12'b111110000000;
   52855: result <= 12'b111110000000;
   52856: result <= 12'b111110000000;
   52857: result <= 12'b111110000000;
   52858: result <= 12'b111110000000;
   52859: result <= 12'b111110000000;
   52860: result <= 12'b111101111111;
   52861: result <= 12'b111101111111;
   52862: result <= 12'b111101111111;
   52863: result <= 12'b111101111111;
   52864: result <= 12'b111101111111;
   52865: result <= 12'b111101111111;
   52866: result <= 12'b111101111111;
   52867: result <= 12'b111101111111;
   52868: result <= 12'b111101111111;
   52869: result <= 12'b111101111111;
   52870: result <= 12'b111101111111;
   52871: result <= 12'b111101111111;
   52872: result <= 12'b111101111111;
   52873: result <= 12'b111101111111;
   52874: result <= 12'b111101111110;
   52875: result <= 12'b111101111110;
   52876: result <= 12'b111101111110;
   52877: result <= 12'b111101111110;
   52878: result <= 12'b111101111110;
   52879: result <= 12'b111101111110;
   52880: result <= 12'b111101111110;
   52881: result <= 12'b111101111110;
   52882: result <= 12'b111101111110;
   52883: result <= 12'b111101111110;
   52884: result <= 12'b111101111110;
   52885: result <= 12'b111101111110;
   52886: result <= 12'b111101111110;
   52887: result <= 12'b111101111110;
   52888: result <= 12'b111101111110;
   52889: result <= 12'b111101111101;
   52890: result <= 12'b111101111101;
   52891: result <= 12'b111101111101;
   52892: result <= 12'b111101111101;
   52893: result <= 12'b111101111101;
   52894: result <= 12'b111101111101;
   52895: result <= 12'b111101111101;
   52896: result <= 12'b111101111101;
   52897: result <= 12'b111101111101;
   52898: result <= 12'b111101111101;
   52899: result <= 12'b111101111101;
   52900: result <= 12'b111101111101;
   52901: result <= 12'b111101111101;
   52902: result <= 12'b111101111101;
   52903: result <= 12'b111101111100;
   52904: result <= 12'b111101111100;
   52905: result <= 12'b111101111100;
   52906: result <= 12'b111101111100;
   52907: result <= 12'b111101111100;
   52908: result <= 12'b111101111100;
   52909: result <= 12'b111101111100;
   52910: result <= 12'b111101111100;
   52911: result <= 12'b111101111100;
   52912: result <= 12'b111101111100;
   52913: result <= 12'b111101111100;
   52914: result <= 12'b111101111100;
   52915: result <= 12'b111101111100;
   52916: result <= 12'b111101111100;
   52917: result <= 12'b111101111100;
   52918: result <= 12'b111101111011;
   52919: result <= 12'b111101111011;
   52920: result <= 12'b111101111011;
   52921: result <= 12'b111101111011;
   52922: result <= 12'b111101111011;
   52923: result <= 12'b111101111011;
   52924: result <= 12'b111101111011;
   52925: result <= 12'b111101111011;
   52926: result <= 12'b111101111011;
   52927: result <= 12'b111101111011;
   52928: result <= 12'b111101111011;
   52929: result <= 12'b111101111011;
   52930: result <= 12'b111101111011;
   52931: result <= 12'b111101111011;
   52932: result <= 12'b111101111010;
   52933: result <= 12'b111101111010;
   52934: result <= 12'b111101111010;
   52935: result <= 12'b111101111010;
   52936: result <= 12'b111101111010;
   52937: result <= 12'b111101111010;
   52938: result <= 12'b111101111010;
   52939: result <= 12'b111101111010;
   52940: result <= 12'b111101111010;
   52941: result <= 12'b111101111010;
   52942: result <= 12'b111101111010;
   52943: result <= 12'b111101111010;
   52944: result <= 12'b111101111010;
   52945: result <= 12'b111101111010;
   52946: result <= 12'b111101111010;
   52947: result <= 12'b111101111001;
   52948: result <= 12'b111101111001;
   52949: result <= 12'b111101111001;
   52950: result <= 12'b111101111001;
   52951: result <= 12'b111101111001;
   52952: result <= 12'b111101111001;
   52953: result <= 12'b111101111001;
   52954: result <= 12'b111101111001;
   52955: result <= 12'b111101111001;
   52956: result <= 12'b111101111001;
   52957: result <= 12'b111101111001;
   52958: result <= 12'b111101111001;
   52959: result <= 12'b111101111001;
   52960: result <= 12'b111101111001;
   52961: result <= 12'b111101111000;
   52962: result <= 12'b111101111000;
   52963: result <= 12'b111101111000;
   52964: result <= 12'b111101111000;
   52965: result <= 12'b111101111000;
   52966: result <= 12'b111101111000;
   52967: result <= 12'b111101111000;
   52968: result <= 12'b111101111000;
   52969: result <= 12'b111101111000;
   52970: result <= 12'b111101111000;
   52971: result <= 12'b111101111000;
   52972: result <= 12'b111101111000;
   52973: result <= 12'b111101111000;
   52974: result <= 12'b111101111000;
   52975: result <= 12'b111101110111;
   52976: result <= 12'b111101110111;
   52977: result <= 12'b111101110111;
   52978: result <= 12'b111101110111;
   52979: result <= 12'b111101110111;
   52980: result <= 12'b111101110111;
   52981: result <= 12'b111101110111;
   52982: result <= 12'b111101110111;
   52983: result <= 12'b111101110111;
   52984: result <= 12'b111101110111;
   52985: result <= 12'b111101110111;
   52986: result <= 12'b111101110111;
   52987: result <= 12'b111101110111;
   52988: result <= 12'b111101110111;
   52989: result <= 12'b111101110110;
   52990: result <= 12'b111101110110;
   52991: result <= 12'b111101110110;
   52992: result <= 12'b111101110110;
   52993: result <= 12'b111101110110;
   52994: result <= 12'b111101110110;
   52995: result <= 12'b111101110110;
   52996: result <= 12'b111101110110;
   52997: result <= 12'b111101110110;
   52998: result <= 12'b111101110110;
   52999: result <= 12'b111101110110;
   53000: result <= 12'b111101110110;
   53001: result <= 12'b111101110110;
   53002: result <= 12'b111101110110;
   53003: result <= 12'b111101110101;
   53004: result <= 12'b111101110101;
   53005: result <= 12'b111101110101;
   53006: result <= 12'b111101110101;
   53007: result <= 12'b111101110101;
   53008: result <= 12'b111101110101;
   53009: result <= 12'b111101110101;
   53010: result <= 12'b111101110101;
   53011: result <= 12'b111101110101;
   53012: result <= 12'b111101110101;
   53013: result <= 12'b111101110101;
   53014: result <= 12'b111101110101;
   53015: result <= 12'b111101110101;
   53016: result <= 12'b111101110101;
   53017: result <= 12'b111101110100;
   53018: result <= 12'b111101110100;
   53019: result <= 12'b111101110100;
   53020: result <= 12'b111101110100;
   53021: result <= 12'b111101110100;
   53022: result <= 12'b111101110100;
   53023: result <= 12'b111101110100;
   53024: result <= 12'b111101110100;
   53025: result <= 12'b111101110100;
   53026: result <= 12'b111101110100;
   53027: result <= 12'b111101110100;
   53028: result <= 12'b111101110100;
   53029: result <= 12'b111101110100;
   53030: result <= 12'b111101110100;
   53031: result <= 12'b111101110011;
   53032: result <= 12'b111101110011;
   53033: result <= 12'b111101110011;
   53034: result <= 12'b111101110011;
   53035: result <= 12'b111101110011;
   53036: result <= 12'b111101110011;
   53037: result <= 12'b111101110011;
   53038: result <= 12'b111101110011;
   53039: result <= 12'b111101110011;
   53040: result <= 12'b111101110011;
   53041: result <= 12'b111101110011;
   53042: result <= 12'b111101110011;
   53043: result <= 12'b111101110011;
   53044: result <= 12'b111101110011;
   53045: result <= 12'b111101110010;
   53046: result <= 12'b111101110010;
   53047: result <= 12'b111101110010;
   53048: result <= 12'b111101110010;
   53049: result <= 12'b111101110010;
   53050: result <= 12'b111101110010;
   53051: result <= 12'b111101110010;
   53052: result <= 12'b111101110010;
   53053: result <= 12'b111101110010;
   53054: result <= 12'b111101110010;
   53055: result <= 12'b111101110010;
   53056: result <= 12'b111101110010;
   53057: result <= 12'b111101110010;
   53058: result <= 12'b111101110010;
   53059: result <= 12'b111101110001;
   53060: result <= 12'b111101110001;
   53061: result <= 12'b111101110001;
   53062: result <= 12'b111101110001;
   53063: result <= 12'b111101110001;
   53064: result <= 12'b111101110001;
   53065: result <= 12'b111101110001;
   53066: result <= 12'b111101110001;
   53067: result <= 12'b111101110001;
   53068: result <= 12'b111101110001;
   53069: result <= 12'b111101110001;
   53070: result <= 12'b111101110001;
   53071: result <= 12'b111101110001;
   53072: result <= 12'b111101110001;
   53073: result <= 12'b111101110000;
   53074: result <= 12'b111101110000;
   53075: result <= 12'b111101110000;
   53076: result <= 12'b111101110000;
   53077: result <= 12'b111101110000;
   53078: result <= 12'b111101110000;
   53079: result <= 12'b111101110000;
   53080: result <= 12'b111101110000;
   53081: result <= 12'b111101110000;
   53082: result <= 12'b111101110000;
   53083: result <= 12'b111101110000;
   53084: result <= 12'b111101110000;
   53085: result <= 12'b111101110000;
   53086: result <= 12'b111101110000;
   53087: result <= 12'b111101101111;
   53088: result <= 12'b111101101111;
   53089: result <= 12'b111101101111;
   53090: result <= 12'b111101101111;
   53091: result <= 12'b111101101111;
   53092: result <= 12'b111101101111;
   53093: result <= 12'b111101101111;
   53094: result <= 12'b111101101111;
   53095: result <= 12'b111101101111;
   53096: result <= 12'b111101101111;
   53097: result <= 12'b111101101111;
   53098: result <= 12'b111101101111;
   53099: result <= 12'b111101101111;
   53100: result <= 12'b111101101111;
   53101: result <= 12'b111101101110;
   53102: result <= 12'b111101101110;
   53103: result <= 12'b111101101110;
   53104: result <= 12'b111101101110;
   53105: result <= 12'b111101101110;
   53106: result <= 12'b111101101110;
   53107: result <= 12'b111101101110;
   53108: result <= 12'b111101101110;
   53109: result <= 12'b111101101110;
   53110: result <= 12'b111101101110;
   53111: result <= 12'b111101101110;
   53112: result <= 12'b111101101110;
   53113: result <= 12'b111101101110;
   53114: result <= 12'b111101101110;
   53115: result <= 12'b111101101101;
   53116: result <= 12'b111101101101;
   53117: result <= 12'b111101101101;
   53118: result <= 12'b111101101101;
   53119: result <= 12'b111101101101;
   53120: result <= 12'b111101101101;
   53121: result <= 12'b111101101101;
   53122: result <= 12'b111101101101;
   53123: result <= 12'b111101101101;
   53124: result <= 12'b111101101101;
   53125: result <= 12'b111101101101;
   53126: result <= 12'b111101101101;
   53127: result <= 12'b111101101101;
   53128: result <= 12'b111101101100;
   53129: result <= 12'b111101101100;
   53130: result <= 12'b111101101100;
   53131: result <= 12'b111101101100;
   53132: result <= 12'b111101101100;
   53133: result <= 12'b111101101100;
   53134: result <= 12'b111101101100;
   53135: result <= 12'b111101101100;
   53136: result <= 12'b111101101100;
   53137: result <= 12'b111101101100;
   53138: result <= 12'b111101101100;
   53139: result <= 12'b111101101100;
   53140: result <= 12'b111101101100;
   53141: result <= 12'b111101101100;
   53142: result <= 12'b111101101011;
   53143: result <= 12'b111101101011;
   53144: result <= 12'b111101101011;
   53145: result <= 12'b111101101011;
   53146: result <= 12'b111101101011;
   53147: result <= 12'b111101101011;
   53148: result <= 12'b111101101011;
   53149: result <= 12'b111101101011;
   53150: result <= 12'b111101101011;
   53151: result <= 12'b111101101011;
   53152: result <= 12'b111101101011;
   53153: result <= 12'b111101101011;
   53154: result <= 12'b111101101011;
   53155: result <= 12'b111101101011;
   53156: result <= 12'b111101101010;
   53157: result <= 12'b111101101010;
   53158: result <= 12'b111101101010;
   53159: result <= 12'b111101101010;
   53160: result <= 12'b111101101010;
   53161: result <= 12'b111101101010;
   53162: result <= 12'b111101101010;
   53163: result <= 12'b111101101010;
   53164: result <= 12'b111101101010;
   53165: result <= 12'b111101101010;
   53166: result <= 12'b111101101010;
   53167: result <= 12'b111101101010;
   53168: result <= 12'b111101101010;
   53169: result <= 12'b111101101001;
   53170: result <= 12'b111101101001;
   53171: result <= 12'b111101101001;
   53172: result <= 12'b111101101001;
   53173: result <= 12'b111101101001;
   53174: result <= 12'b111101101001;
   53175: result <= 12'b111101101001;
   53176: result <= 12'b111101101001;
   53177: result <= 12'b111101101001;
   53178: result <= 12'b111101101001;
   53179: result <= 12'b111101101001;
   53180: result <= 12'b111101101001;
   53181: result <= 12'b111101101001;
   53182: result <= 12'b111101101001;
   53183: result <= 12'b111101101000;
   53184: result <= 12'b111101101000;
   53185: result <= 12'b111101101000;
   53186: result <= 12'b111101101000;
   53187: result <= 12'b111101101000;
   53188: result <= 12'b111101101000;
   53189: result <= 12'b111101101000;
   53190: result <= 12'b111101101000;
   53191: result <= 12'b111101101000;
   53192: result <= 12'b111101101000;
   53193: result <= 12'b111101101000;
   53194: result <= 12'b111101101000;
   53195: result <= 12'b111101101000;
   53196: result <= 12'b111101100111;
   53197: result <= 12'b111101100111;
   53198: result <= 12'b111101100111;
   53199: result <= 12'b111101100111;
   53200: result <= 12'b111101100111;
   53201: result <= 12'b111101100111;
   53202: result <= 12'b111101100111;
   53203: result <= 12'b111101100111;
   53204: result <= 12'b111101100111;
   53205: result <= 12'b111101100111;
   53206: result <= 12'b111101100111;
   53207: result <= 12'b111101100111;
   53208: result <= 12'b111101100111;
   53209: result <= 12'b111101100111;
   53210: result <= 12'b111101100110;
   53211: result <= 12'b111101100110;
   53212: result <= 12'b111101100110;
   53213: result <= 12'b111101100110;
   53214: result <= 12'b111101100110;
   53215: result <= 12'b111101100110;
   53216: result <= 12'b111101100110;
   53217: result <= 12'b111101100110;
   53218: result <= 12'b111101100110;
   53219: result <= 12'b111101100110;
   53220: result <= 12'b111101100110;
   53221: result <= 12'b111101100110;
   53222: result <= 12'b111101100110;
   53223: result <= 12'b111101100101;
   53224: result <= 12'b111101100101;
   53225: result <= 12'b111101100101;
   53226: result <= 12'b111101100101;
   53227: result <= 12'b111101100101;
   53228: result <= 12'b111101100101;
   53229: result <= 12'b111101100101;
   53230: result <= 12'b111101100101;
   53231: result <= 12'b111101100101;
   53232: result <= 12'b111101100101;
   53233: result <= 12'b111101100101;
   53234: result <= 12'b111101100101;
   53235: result <= 12'b111101100101;
   53236: result <= 12'b111101100101;
   53237: result <= 12'b111101100100;
   53238: result <= 12'b111101100100;
   53239: result <= 12'b111101100100;
   53240: result <= 12'b111101100100;
   53241: result <= 12'b111101100100;
   53242: result <= 12'b111101100100;
   53243: result <= 12'b111101100100;
   53244: result <= 12'b111101100100;
   53245: result <= 12'b111101100100;
   53246: result <= 12'b111101100100;
   53247: result <= 12'b111101100100;
   53248: result <= 12'b111101100100;
   53249: result <= 12'b111101100100;
   53250: result <= 12'b111101100011;
   53251: result <= 12'b111101100011;
   53252: result <= 12'b111101100011;
   53253: result <= 12'b111101100011;
   53254: result <= 12'b111101100011;
   53255: result <= 12'b111101100011;
   53256: result <= 12'b111101100011;
   53257: result <= 12'b111101100011;
   53258: result <= 12'b111101100011;
   53259: result <= 12'b111101100011;
   53260: result <= 12'b111101100011;
   53261: result <= 12'b111101100011;
   53262: result <= 12'b111101100011;
   53263: result <= 12'b111101100010;
   53264: result <= 12'b111101100010;
   53265: result <= 12'b111101100010;
   53266: result <= 12'b111101100010;
   53267: result <= 12'b111101100010;
   53268: result <= 12'b111101100010;
   53269: result <= 12'b111101100010;
   53270: result <= 12'b111101100010;
   53271: result <= 12'b111101100010;
   53272: result <= 12'b111101100010;
   53273: result <= 12'b111101100010;
   53274: result <= 12'b111101100010;
   53275: result <= 12'b111101100010;
   53276: result <= 12'b111101100001;
   53277: result <= 12'b111101100001;
   53278: result <= 12'b111101100001;
   53279: result <= 12'b111101100001;
   53280: result <= 12'b111101100001;
   53281: result <= 12'b111101100001;
   53282: result <= 12'b111101100001;
   53283: result <= 12'b111101100001;
   53284: result <= 12'b111101100001;
   53285: result <= 12'b111101100001;
   53286: result <= 12'b111101100001;
   53287: result <= 12'b111101100001;
   53288: result <= 12'b111101100001;
   53289: result <= 12'b111101100001;
   53290: result <= 12'b111101100000;
   53291: result <= 12'b111101100000;
   53292: result <= 12'b111101100000;
   53293: result <= 12'b111101100000;
   53294: result <= 12'b111101100000;
   53295: result <= 12'b111101100000;
   53296: result <= 12'b111101100000;
   53297: result <= 12'b111101100000;
   53298: result <= 12'b111101100000;
   53299: result <= 12'b111101100000;
   53300: result <= 12'b111101100000;
   53301: result <= 12'b111101100000;
   53302: result <= 12'b111101100000;
   53303: result <= 12'b111101011111;
   53304: result <= 12'b111101011111;
   53305: result <= 12'b111101011111;
   53306: result <= 12'b111101011111;
   53307: result <= 12'b111101011111;
   53308: result <= 12'b111101011111;
   53309: result <= 12'b111101011111;
   53310: result <= 12'b111101011111;
   53311: result <= 12'b111101011111;
   53312: result <= 12'b111101011111;
   53313: result <= 12'b111101011111;
   53314: result <= 12'b111101011111;
   53315: result <= 12'b111101011111;
   53316: result <= 12'b111101011110;
   53317: result <= 12'b111101011110;
   53318: result <= 12'b111101011110;
   53319: result <= 12'b111101011110;
   53320: result <= 12'b111101011110;
   53321: result <= 12'b111101011110;
   53322: result <= 12'b111101011110;
   53323: result <= 12'b111101011110;
   53324: result <= 12'b111101011110;
   53325: result <= 12'b111101011110;
   53326: result <= 12'b111101011110;
   53327: result <= 12'b111101011110;
   53328: result <= 12'b111101011110;
   53329: result <= 12'b111101011101;
   53330: result <= 12'b111101011101;
   53331: result <= 12'b111101011101;
   53332: result <= 12'b111101011101;
   53333: result <= 12'b111101011101;
   53334: result <= 12'b111101011101;
   53335: result <= 12'b111101011101;
   53336: result <= 12'b111101011101;
   53337: result <= 12'b111101011101;
   53338: result <= 12'b111101011101;
   53339: result <= 12'b111101011101;
   53340: result <= 12'b111101011101;
   53341: result <= 12'b111101011101;
   53342: result <= 12'b111101011100;
   53343: result <= 12'b111101011100;
   53344: result <= 12'b111101011100;
   53345: result <= 12'b111101011100;
   53346: result <= 12'b111101011100;
   53347: result <= 12'b111101011100;
   53348: result <= 12'b111101011100;
   53349: result <= 12'b111101011100;
   53350: result <= 12'b111101011100;
   53351: result <= 12'b111101011100;
   53352: result <= 12'b111101011100;
   53353: result <= 12'b111101011100;
   53354: result <= 12'b111101011100;
   53355: result <= 12'b111101011011;
   53356: result <= 12'b111101011011;
   53357: result <= 12'b111101011011;
   53358: result <= 12'b111101011011;
   53359: result <= 12'b111101011011;
   53360: result <= 12'b111101011011;
   53361: result <= 12'b111101011011;
   53362: result <= 12'b111101011011;
   53363: result <= 12'b111101011011;
   53364: result <= 12'b111101011011;
   53365: result <= 12'b111101011011;
   53366: result <= 12'b111101011011;
   53367: result <= 12'b111101011011;
   53368: result <= 12'b111101011010;
   53369: result <= 12'b111101011010;
   53370: result <= 12'b111101011010;
   53371: result <= 12'b111101011010;
   53372: result <= 12'b111101011010;
   53373: result <= 12'b111101011010;
   53374: result <= 12'b111101011010;
   53375: result <= 12'b111101011010;
   53376: result <= 12'b111101011010;
   53377: result <= 12'b111101011010;
   53378: result <= 12'b111101011010;
   53379: result <= 12'b111101011010;
   53380: result <= 12'b111101011010;
   53381: result <= 12'b111101011001;
   53382: result <= 12'b111101011001;
   53383: result <= 12'b111101011001;
   53384: result <= 12'b111101011001;
   53385: result <= 12'b111101011001;
   53386: result <= 12'b111101011001;
   53387: result <= 12'b111101011001;
   53388: result <= 12'b111101011001;
   53389: result <= 12'b111101011001;
   53390: result <= 12'b111101011001;
   53391: result <= 12'b111101011001;
   53392: result <= 12'b111101011001;
   53393: result <= 12'b111101011001;
   53394: result <= 12'b111101011000;
   53395: result <= 12'b111101011000;
   53396: result <= 12'b111101011000;
   53397: result <= 12'b111101011000;
   53398: result <= 12'b111101011000;
   53399: result <= 12'b111101011000;
   53400: result <= 12'b111101011000;
   53401: result <= 12'b111101011000;
   53402: result <= 12'b111101011000;
   53403: result <= 12'b111101011000;
   53404: result <= 12'b111101011000;
   53405: result <= 12'b111101011000;
   53406: result <= 12'b111101011000;
   53407: result <= 12'b111101010111;
   53408: result <= 12'b111101010111;
   53409: result <= 12'b111101010111;
   53410: result <= 12'b111101010111;
   53411: result <= 12'b111101010111;
   53412: result <= 12'b111101010111;
   53413: result <= 12'b111101010111;
   53414: result <= 12'b111101010111;
   53415: result <= 12'b111101010111;
   53416: result <= 12'b111101010111;
   53417: result <= 12'b111101010111;
   53418: result <= 12'b111101010111;
   53419: result <= 12'b111101010111;
   53420: result <= 12'b111101010110;
   53421: result <= 12'b111101010110;
   53422: result <= 12'b111101010110;
   53423: result <= 12'b111101010110;
   53424: result <= 12'b111101010110;
   53425: result <= 12'b111101010110;
   53426: result <= 12'b111101010110;
   53427: result <= 12'b111101010110;
   53428: result <= 12'b111101010110;
   53429: result <= 12'b111101010110;
   53430: result <= 12'b111101010110;
   53431: result <= 12'b111101010110;
   53432: result <= 12'b111101010101;
   53433: result <= 12'b111101010101;
   53434: result <= 12'b111101010101;
   53435: result <= 12'b111101010101;
   53436: result <= 12'b111101010101;
   53437: result <= 12'b111101010101;
   53438: result <= 12'b111101010101;
   53439: result <= 12'b111101010101;
   53440: result <= 12'b111101010101;
   53441: result <= 12'b111101010101;
   53442: result <= 12'b111101010101;
   53443: result <= 12'b111101010101;
   53444: result <= 12'b111101010101;
   53445: result <= 12'b111101010100;
   53446: result <= 12'b111101010100;
   53447: result <= 12'b111101010100;
   53448: result <= 12'b111101010100;
   53449: result <= 12'b111101010100;
   53450: result <= 12'b111101010100;
   53451: result <= 12'b111101010100;
   53452: result <= 12'b111101010100;
   53453: result <= 12'b111101010100;
   53454: result <= 12'b111101010100;
   53455: result <= 12'b111101010100;
   53456: result <= 12'b111101010100;
   53457: result <= 12'b111101010100;
   53458: result <= 12'b111101010011;
   53459: result <= 12'b111101010011;
   53460: result <= 12'b111101010011;
   53461: result <= 12'b111101010011;
   53462: result <= 12'b111101010011;
   53463: result <= 12'b111101010011;
   53464: result <= 12'b111101010011;
   53465: result <= 12'b111101010011;
   53466: result <= 12'b111101010011;
   53467: result <= 12'b111101010011;
   53468: result <= 12'b111101010011;
   53469: result <= 12'b111101010011;
   53470: result <= 12'b111101010010;
   53471: result <= 12'b111101010010;
   53472: result <= 12'b111101010010;
   53473: result <= 12'b111101010010;
   53474: result <= 12'b111101010010;
   53475: result <= 12'b111101010010;
   53476: result <= 12'b111101010010;
   53477: result <= 12'b111101010010;
   53478: result <= 12'b111101010010;
   53479: result <= 12'b111101010010;
   53480: result <= 12'b111101010010;
   53481: result <= 12'b111101010010;
   53482: result <= 12'b111101010010;
   53483: result <= 12'b111101010001;
   53484: result <= 12'b111101010001;
   53485: result <= 12'b111101010001;
   53486: result <= 12'b111101010001;
   53487: result <= 12'b111101010001;
   53488: result <= 12'b111101010001;
   53489: result <= 12'b111101010001;
   53490: result <= 12'b111101010001;
   53491: result <= 12'b111101010001;
   53492: result <= 12'b111101010001;
   53493: result <= 12'b111101010001;
   53494: result <= 12'b111101010001;
   53495: result <= 12'b111101010001;
   53496: result <= 12'b111101010000;
   53497: result <= 12'b111101010000;
   53498: result <= 12'b111101010000;
   53499: result <= 12'b111101010000;
   53500: result <= 12'b111101010000;
   53501: result <= 12'b111101010000;
   53502: result <= 12'b111101010000;
   53503: result <= 12'b111101010000;
   53504: result <= 12'b111101010000;
   53505: result <= 12'b111101010000;
   53506: result <= 12'b111101010000;
   53507: result <= 12'b111101010000;
   53508: result <= 12'b111101001111;
   53509: result <= 12'b111101001111;
   53510: result <= 12'b111101001111;
   53511: result <= 12'b111101001111;
   53512: result <= 12'b111101001111;
   53513: result <= 12'b111101001111;
   53514: result <= 12'b111101001111;
   53515: result <= 12'b111101001111;
   53516: result <= 12'b111101001111;
   53517: result <= 12'b111101001111;
   53518: result <= 12'b111101001111;
   53519: result <= 12'b111101001111;
   53520: result <= 12'b111101001111;
   53521: result <= 12'b111101001110;
   53522: result <= 12'b111101001110;
   53523: result <= 12'b111101001110;
   53524: result <= 12'b111101001110;
   53525: result <= 12'b111101001110;
   53526: result <= 12'b111101001110;
   53527: result <= 12'b111101001110;
   53528: result <= 12'b111101001110;
   53529: result <= 12'b111101001110;
   53530: result <= 12'b111101001110;
   53531: result <= 12'b111101001110;
   53532: result <= 12'b111101001110;
   53533: result <= 12'b111101001101;
   53534: result <= 12'b111101001101;
   53535: result <= 12'b111101001101;
   53536: result <= 12'b111101001101;
   53537: result <= 12'b111101001101;
   53538: result <= 12'b111101001101;
   53539: result <= 12'b111101001101;
   53540: result <= 12'b111101001101;
   53541: result <= 12'b111101001101;
   53542: result <= 12'b111101001101;
   53543: result <= 12'b111101001101;
   53544: result <= 12'b111101001101;
   53545: result <= 12'b111101001101;
   53546: result <= 12'b111101001100;
   53547: result <= 12'b111101001100;
   53548: result <= 12'b111101001100;
   53549: result <= 12'b111101001100;
   53550: result <= 12'b111101001100;
   53551: result <= 12'b111101001100;
   53552: result <= 12'b111101001100;
   53553: result <= 12'b111101001100;
   53554: result <= 12'b111101001100;
   53555: result <= 12'b111101001100;
   53556: result <= 12'b111101001100;
   53557: result <= 12'b111101001100;
   53558: result <= 12'b111101001011;
   53559: result <= 12'b111101001011;
   53560: result <= 12'b111101001011;
   53561: result <= 12'b111101001011;
   53562: result <= 12'b111101001011;
   53563: result <= 12'b111101001011;
   53564: result <= 12'b111101001011;
   53565: result <= 12'b111101001011;
   53566: result <= 12'b111101001011;
   53567: result <= 12'b111101001011;
   53568: result <= 12'b111101001011;
   53569: result <= 12'b111101001011;
   53570: result <= 12'b111101001011;
   53571: result <= 12'b111101001010;
   53572: result <= 12'b111101001010;
   53573: result <= 12'b111101001010;
   53574: result <= 12'b111101001010;
   53575: result <= 12'b111101001010;
   53576: result <= 12'b111101001010;
   53577: result <= 12'b111101001010;
   53578: result <= 12'b111101001010;
   53579: result <= 12'b111101001010;
   53580: result <= 12'b111101001010;
   53581: result <= 12'b111101001010;
   53582: result <= 12'b111101001010;
   53583: result <= 12'b111101001001;
   53584: result <= 12'b111101001001;
   53585: result <= 12'b111101001001;
   53586: result <= 12'b111101001001;
   53587: result <= 12'b111101001001;
   53588: result <= 12'b111101001001;
   53589: result <= 12'b111101001001;
   53590: result <= 12'b111101001001;
   53591: result <= 12'b111101001001;
   53592: result <= 12'b111101001001;
   53593: result <= 12'b111101001001;
   53594: result <= 12'b111101001001;
   53595: result <= 12'b111101001000;
   53596: result <= 12'b111101001000;
   53597: result <= 12'b111101001000;
   53598: result <= 12'b111101001000;
   53599: result <= 12'b111101001000;
   53600: result <= 12'b111101001000;
   53601: result <= 12'b111101001000;
   53602: result <= 12'b111101001000;
   53603: result <= 12'b111101001000;
   53604: result <= 12'b111101001000;
   53605: result <= 12'b111101001000;
   53606: result <= 12'b111101001000;
   53607: result <= 12'b111101001000;
   53608: result <= 12'b111101000111;
   53609: result <= 12'b111101000111;
   53610: result <= 12'b111101000111;
   53611: result <= 12'b111101000111;
   53612: result <= 12'b111101000111;
   53613: result <= 12'b111101000111;
   53614: result <= 12'b111101000111;
   53615: result <= 12'b111101000111;
   53616: result <= 12'b111101000111;
   53617: result <= 12'b111101000111;
   53618: result <= 12'b111101000111;
   53619: result <= 12'b111101000111;
   53620: result <= 12'b111101000110;
   53621: result <= 12'b111101000110;
   53622: result <= 12'b111101000110;
   53623: result <= 12'b111101000110;
   53624: result <= 12'b111101000110;
   53625: result <= 12'b111101000110;
   53626: result <= 12'b111101000110;
   53627: result <= 12'b111101000110;
   53628: result <= 12'b111101000110;
   53629: result <= 12'b111101000110;
   53630: result <= 12'b111101000110;
   53631: result <= 12'b111101000110;
   53632: result <= 12'b111101000101;
   53633: result <= 12'b111101000101;
   53634: result <= 12'b111101000101;
   53635: result <= 12'b111101000101;
   53636: result <= 12'b111101000101;
   53637: result <= 12'b111101000101;
   53638: result <= 12'b111101000101;
   53639: result <= 12'b111101000101;
   53640: result <= 12'b111101000101;
   53641: result <= 12'b111101000101;
   53642: result <= 12'b111101000101;
   53643: result <= 12'b111101000101;
   53644: result <= 12'b111101000100;
   53645: result <= 12'b111101000100;
   53646: result <= 12'b111101000100;
   53647: result <= 12'b111101000100;
   53648: result <= 12'b111101000100;
   53649: result <= 12'b111101000100;
   53650: result <= 12'b111101000100;
   53651: result <= 12'b111101000100;
   53652: result <= 12'b111101000100;
   53653: result <= 12'b111101000100;
   53654: result <= 12'b111101000100;
   53655: result <= 12'b111101000100;
   53656: result <= 12'b111101000100;
   53657: result <= 12'b111101000011;
   53658: result <= 12'b111101000011;
   53659: result <= 12'b111101000011;
   53660: result <= 12'b111101000011;
   53661: result <= 12'b111101000011;
   53662: result <= 12'b111101000011;
   53663: result <= 12'b111101000011;
   53664: result <= 12'b111101000011;
   53665: result <= 12'b111101000011;
   53666: result <= 12'b111101000011;
   53667: result <= 12'b111101000011;
   53668: result <= 12'b111101000011;
   53669: result <= 12'b111101000010;
   53670: result <= 12'b111101000010;
   53671: result <= 12'b111101000010;
   53672: result <= 12'b111101000010;
   53673: result <= 12'b111101000010;
   53674: result <= 12'b111101000010;
   53675: result <= 12'b111101000010;
   53676: result <= 12'b111101000010;
   53677: result <= 12'b111101000010;
   53678: result <= 12'b111101000010;
   53679: result <= 12'b111101000010;
   53680: result <= 12'b111101000010;
   53681: result <= 12'b111101000001;
   53682: result <= 12'b111101000001;
   53683: result <= 12'b111101000001;
   53684: result <= 12'b111101000001;
   53685: result <= 12'b111101000001;
   53686: result <= 12'b111101000001;
   53687: result <= 12'b111101000001;
   53688: result <= 12'b111101000001;
   53689: result <= 12'b111101000001;
   53690: result <= 12'b111101000001;
   53691: result <= 12'b111101000001;
   53692: result <= 12'b111101000001;
   53693: result <= 12'b111101000000;
   53694: result <= 12'b111101000000;
   53695: result <= 12'b111101000000;
   53696: result <= 12'b111101000000;
   53697: result <= 12'b111101000000;
   53698: result <= 12'b111101000000;
   53699: result <= 12'b111101000000;
   53700: result <= 12'b111101000000;
   53701: result <= 12'b111101000000;
   53702: result <= 12'b111101000000;
   53703: result <= 12'b111101000000;
   53704: result <= 12'b111101000000;
   53705: result <= 12'b111100111111;
   53706: result <= 12'b111100111111;
   53707: result <= 12'b111100111111;
   53708: result <= 12'b111100111111;
   53709: result <= 12'b111100111111;
   53710: result <= 12'b111100111111;
   53711: result <= 12'b111100111111;
   53712: result <= 12'b111100111111;
   53713: result <= 12'b111100111111;
   53714: result <= 12'b111100111111;
   53715: result <= 12'b111100111111;
   53716: result <= 12'b111100111111;
   53717: result <= 12'b111100111110;
   53718: result <= 12'b111100111110;
   53719: result <= 12'b111100111110;
   53720: result <= 12'b111100111110;
   53721: result <= 12'b111100111110;
   53722: result <= 12'b111100111110;
   53723: result <= 12'b111100111110;
   53724: result <= 12'b111100111110;
   53725: result <= 12'b111100111110;
   53726: result <= 12'b111100111110;
   53727: result <= 12'b111100111110;
   53728: result <= 12'b111100111110;
   53729: result <= 12'b111100111101;
   53730: result <= 12'b111100111101;
   53731: result <= 12'b111100111101;
   53732: result <= 12'b111100111101;
   53733: result <= 12'b111100111101;
   53734: result <= 12'b111100111101;
   53735: result <= 12'b111100111101;
   53736: result <= 12'b111100111101;
   53737: result <= 12'b111100111101;
   53738: result <= 12'b111100111101;
   53739: result <= 12'b111100111101;
   53740: result <= 12'b111100111101;
   53741: result <= 12'b111100111100;
   53742: result <= 12'b111100111100;
   53743: result <= 12'b111100111100;
   53744: result <= 12'b111100111100;
   53745: result <= 12'b111100111100;
   53746: result <= 12'b111100111100;
   53747: result <= 12'b111100111100;
   53748: result <= 12'b111100111100;
   53749: result <= 12'b111100111100;
   53750: result <= 12'b111100111100;
   53751: result <= 12'b111100111100;
   53752: result <= 12'b111100111100;
   53753: result <= 12'b111100111011;
   53754: result <= 12'b111100111011;
   53755: result <= 12'b111100111011;
   53756: result <= 12'b111100111011;
   53757: result <= 12'b111100111011;
   53758: result <= 12'b111100111011;
   53759: result <= 12'b111100111011;
   53760: result <= 12'b111100111011;
   53761: result <= 12'b111100111011;
   53762: result <= 12'b111100111011;
   53763: result <= 12'b111100111011;
   53764: result <= 12'b111100111011;
   53765: result <= 12'b111100111010;
   53766: result <= 12'b111100111010;
   53767: result <= 12'b111100111010;
   53768: result <= 12'b111100111010;
   53769: result <= 12'b111100111010;
   53770: result <= 12'b111100111010;
   53771: result <= 12'b111100111010;
   53772: result <= 12'b111100111010;
   53773: result <= 12'b111100111010;
   53774: result <= 12'b111100111010;
   53775: result <= 12'b111100111010;
   53776: result <= 12'b111100111010;
   53777: result <= 12'b111100111001;
   53778: result <= 12'b111100111001;
   53779: result <= 12'b111100111001;
   53780: result <= 12'b111100111001;
   53781: result <= 12'b111100111001;
   53782: result <= 12'b111100111001;
   53783: result <= 12'b111100111001;
   53784: result <= 12'b111100111001;
   53785: result <= 12'b111100111001;
   53786: result <= 12'b111100111001;
   53787: result <= 12'b111100111001;
   53788: result <= 12'b111100111001;
   53789: result <= 12'b111100111000;
   53790: result <= 12'b111100111000;
   53791: result <= 12'b111100111000;
   53792: result <= 12'b111100111000;
   53793: result <= 12'b111100111000;
   53794: result <= 12'b111100111000;
   53795: result <= 12'b111100111000;
   53796: result <= 12'b111100111000;
   53797: result <= 12'b111100111000;
   53798: result <= 12'b111100111000;
   53799: result <= 12'b111100111000;
   53800: result <= 12'b111100110111;
   53801: result <= 12'b111100110111;
   53802: result <= 12'b111100110111;
   53803: result <= 12'b111100110111;
   53804: result <= 12'b111100110111;
   53805: result <= 12'b111100110111;
   53806: result <= 12'b111100110111;
   53807: result <= 12'b111100110111;
   53808: result <= 12'b111100110111;
   53809: result <= 12'b111100110111;
   53810: result <= 12'b111100110111;
   53811: result <= 12'b111100110111;
   53812: result <= 12'b111100110110;
   53813: result <= 12'b111100110110;
   53814: result <= 12'b111100110110;
   53815: result <= 12'b111100110110;
   53816: result <= 12'b111100110110;
   53817: result <= 12'b111100110110;
   53818: result <= 12'b111100110110;
   53819: result <= 12'b111100110110;
   53820: result <= 12'b111100110110;
   53821: result <= 12'b111100110110;
   53822: result <= 12'b111100110110;
   53823: result <= 12'b111100110110;
   53824: result <= 12'b111100110101;
   53825: result <= 12'b111100110101;
   53826: result <= 12'b111100110101;
   53827: result <= 12'b111100110101;
   53828: result <= 12'b111100110101;
   53829: result <= 12'b111100110101;
   53830: result <= 12'b111100110101;
   53831: result <= 12'b111100110101;
   53832: result <= 12'b111100110101;
   53833: result <= 12'b111100110101;
   53834: result <= 12'b111100110101;
   53835: result <= 12'b111100110101;
   53836: result <= 12'b111100110100;
   53837: result <= 12'b111100110100;
   53838: result <= 12'b111100110100;
   53839: result <= 12'b111100110100;
   53840: result <= 12'b111100110100;
   53841: result <= 12'b111100110100;
   53842: result <= 12'b111100110100;
   53843: result <= 12'b111100110100;
   53844: result <= 12'b111100110100;
   53845: result <= 12'b111100110100;
   53846: result <= 12'b111100110100;
   53847: result <= 12'b111100110100;
   53848: result <= 12'b111100110011;
   53849: result <= 12'b111100110011;
   53850: result <= 12'b111100110011;
   53851: result <= 12'b111100110011;
   53852: result <= 12'b111100110011;
   53853: result <= 12'b111100110011;
   53854: result <= 12'b111100110011;
   53855: result <= 12'b111100110011;
   53856: result <= 12'b111100110011;
   53857: result <= 12'b111100110011;
   53858: result <= 12'b111100110011;
   53859: result <= 12'b111100110010;
   53860: result <= 12'b111100110010;
   53861: result <= 12'b111100110010;
   53862: result <= 12'b111100110010;
   53863: result <= 12'b111100110010;
   53864: result <= 12'b111100110010;
   53865: result <= 12'b111100110010;
   53866: result <= 12'b111100110010;
   53867: result <= 12'b111100110010;
   53868: result <= 12'b111100110010;
   53869: result <= 12'b111100110010;
   53870: result <= 12'b111100110010;
   53871: result <= 12'b111100110001;
   53872: result <= 12'b111100110001;
   53873: result <= 12'b111100110001;
   53874: result <= 12'b111100110001;
   53875: result <= 12'b111100110001;
   53876: result <= 12'b111100110001;
   53877: result <= 12'b111100110001;
   53878: result <= 12'b111100110001;
   53879: result <= 12'b111100110001;
   53880: result <= 12'b111100110001;
   53881: result <= 12'b111100110001;
   53882: result <= 12'b111100110001;
   53883: result <= 12'b111100110000;
   53884: result <= 12'b111100110000;
   53885: result <= 12'b111100110000;
   53886: result <= 12'b111100110000;
   53887: result <= 12'b111100110000;
   53888: result <= 12'b111100110000;
   53889: result <= 12'b111100110000;
   53890: result <= 12'b111100110000;
   53891: result <= 12'b111100110000;
   53892: result <= 12'b111100110000;
   53893: result <= 12'b111100110000;
   53894: result <= 12'b111100101111;
   53895: result <= 12'b111100101111;
   53896: result <= 12'b111100101111;
   53897: result <= 12'b111100101111;
   53898: result <= 12'b111100101111;
   53899: result <= 12'b111100101111;
   53900: result <= 12'b111100101111;
   53901: result <= 12'b111100101111;
   53902: result <= 12'b111100101111;
   53903: result <= 12'b111100101111;
   53904: result <= 12'b111100101111;
   53905: result <= 12'b111100101111;
   53906: result <= 12'b111100101110;
   53907: result <= 12'b111100101110;
   53908: result <= 12'b111100101110;
   53909: result <= 12'b111100101110;
   53910: result <= 12'b111100101110;
   53911: result <= 12'b111100101110;
   53912: result <= 12'b111100101110;
   53913: result <= 12'b111100101110;
   53914: result <= 12'b111100101110;
   53915: result <= 12'b111100101110;
   53916: result <= 12'b111100101110;
   53917: result <= 12'b111100101101;
   53918: result <= 12'b111100101101;
   53919: result <= 12'b111100101101;
   53920: result <= 12'b111100101101;
   53921: result <= 12'b111100101101;
   53922: result <= 12'b111100101101;
   53923: result <= 12'b111100101101;
   53924: result <= 12'b111100101101;
   53925: result <= 12'b111100101101;
   53926: result <= 12'b111100101101;
   53927: result <= 12'b111100101101;
   53928: result <= 12'b111100101101;
   53929: result <= 12'b111100101100;
   53930: result <= 12'b111100101100;
   53931: result <= 12'b111100101100;
   53932: result <= 12'b111100101100;
   53933: result <= 12'b111100101100;
   53934: result <= 12'b111100101100;
   53935: result <= 12'b111100101100;
   53936: result <= 12'b111100101100;
   53937: result <= 12'b111100101100;
   53938: result <= 12'b111100101100;
   53939: result <= 12'b111100101100;
   53940: result <= 12'b111100101011;
   53941: result <= 12'b111100101011;
   53942: result <= 12'b111100101011;
   53943: result <= 12'b111100101011;
   53944: result <= 12'b111100101011;
   53945: result <= 12'b111100101011;
   53946: result <= 12'b111100101011;
   53947: result <= 12'b111100101011;
   53948: result <= 12'b111100101011;
   53949: result <= 12'b111100101011;
   53950: result <= 12'b111100101011;
   53951: result <= 12'b111100101011;
   53952: result <= 12'b111100101010;
   53953: result <= 12'b111100101010;
   53954: result <= 12'b111100101010;
   53955: result <= 12'b111100101010;
   53956: result <= 12'b111100101010;
   53957: result <= 12'b111100101010;
   53958: result <= 12'b111100101010;
   53959: result <= 12'b111100101010;
   53960: result <= 12'b111100101010;
   53961: result <= 12'b111100101010;
   53962: result <= 12'b111100101010;
   53963: result <= 12'b111100101001;
   53964: result <= 12'b111100101001;
   53965: result <= 12'b111100101001;
   53966: result <= 12'b111100101001;
   53967: result <= 12'b111100101001;
   53968: result <= 12'b111100101001;
   53969: result <= 12'b111100101001;
   53970: result <= 12'b111100101001;
   53971: result <= 12'b111100101001;
   53972: result <= 12'b111100101001;
   53973: result <= 12'b111100101001;
   53974: result <= 12'b111100101001;
   53975: result <= 12'b111100101000;
   53976: result <= 12'b111100101000;
   53977: result <= 12'b111100101000;
   53978: result <= 12'b111100101000;
   53979: result <= 12'b111100101000;
   53980: result <= 12'b111100101000;
   53981: result <= 12'b111100101000;
   53982: result <= 12'b111100101000;
   53983: result <= 12'b111100101000;
   53984: result <= 12'b111100101000;
   53985: result <= 12'b111100101000;
   53986: result <= 12'b111100100111;
   53987: result <= 12'b111100100111;
   53988: result <= 12'b111100100111;
   53989: result <= 12'b111100100111;
   53990: result <= 12'b111100100111;
   53991: result <= 12'b111100100111;
   53992: result <= 12'b111100100111;
   53993: result <= 12'b111100100111;
   53994: result <= 12'b111100100111;
   53995: result <= 12'b111100100111;
   53996: result <= 12'b111100100111;
   53997: result <= 12'b111100100110;
   53998: result <= 12'b111100100110;
   53999: result <= 12'b111100100110;
   54000: result <= 12'b111100100110;
   54001: result <= 12'b111100100110;
   54002: result <= 12'b111100100110;
   54003: result <= 12'b111100100110;
   54004: result <= 12'b111100100110;
   54005: result <= 12'b111100100110;
   54006: result <= 12'b111100100110;
   54007: result <= 12'b111100100110;
   54008: result <= 12'b111100100110;
   54009: result <= 12'b111100100101;
   54010: result <= 12'b111100100101;
   54011: result <= 12'b111100100101;
   54012: result <= 12'b111100100101;
   54013: result <= 12'b111100100101;
   54014: result <= 12'b111100100101;
   54015: result <= 12'b111100100101;
   54016: result <= 12'b111100100101;
   54017: result <= 12'b111100100101;
   54018: result <= 12'b111100100101;
   54019: result <= 12'b111100100101;
   54020: result <= 12'b111100100100;
   54021: result <= 12'b111100100100;
   54022: result <= 12'b111100100100;
   54023: result <= 12'b111100100100;
   54024: result <= 12'b111100100100;
   54025: result <= 12'b111100100100;
   54026: result <= 12'b111100100100;
   54027: result <= 12'b111100100100;
   54028: result <= 12'b111100100100;
   54029: result <= 12'b111100100100;
   54030: result <= 12'b111100100100;
   54031: result <= 12'b111100100011;
   54032: result <= 12'b111100100011;
   54033: result <= 12'b111100100011;
   54034: result <= 12'b111100100011;
   54035: result <= 12'b111100100011;
   54036: result <= 12'b111100100011;
   54037: result <= 12'b111100100011;
   54038: result <= 12'b111100100011;
   54039: result <= 12'b111100100011;
   54040: result <= 12'b111100100011;
   54041: result <= 12'b111100100011;
   54042: result <= 12'b111100100011;
   54043: result <= 12'b111100100010;
   54044: result <= 12'b111100100010;
   54045: result <= 12'b111100100010;
   54046: result <= 12'b111100100010;
   54047: result <= 12'b111100100010;
   54048: result <= 12'b111100100010;
   54049: result <= 12'b111100100010;
   54050: result <= 12'b111100100010;
   54051: result <= 12'b111100100010;
   54052: result <= 12'b111100100010;
   54053: result <= 12'b111100100010;
   54054: result <= 12'b111100100001;
   54055: result <= 12'b111100100001;
   54056: result <= 12'b111100100001;
   54057: result <= 12'b111100100001;
   54058: result <= 12'b111100100001;
   54059: result <= 12'b111100100001;
   54060: result <= 12'b111100100001;
   54061: result <= 12'b111100100001;
   54062: result <= 12'b111100100001;
   54063: result <= 12'b111100100001;
   54064: result <= 12'b111100100001;
   54065: result <= 12'b111100100000;
   54066: result <= 12'b111100100000;
   54067: result <= 12'b111100100000;
   54068: result <= 12'b111100100000;
   54069: result <= 12'b111100100000;
   54070: result <= 12'b111100100000;
   54071: result <= 12'b111100100000;
   54072: result <= 12'b111100100000;
   54073: result <= 12'b111100100000;
   54074: result <= 12'b111100100000;
   54075: result <= 12'b111100100000;
   54076: result <= 12'b111100011111;
   54077: result <= 12'b111100011111;
   54078: result <= 12'b111100011111;
   54079: result <= 12'b111100011111;
   54080: result <= 12'b111100011111;
   54081: result <= 12'b111100011111;
   54082: result <= 12'b111100011111;
   54083: result <= 12'b111100011111;
   54084: result <= 12'b111100011111;
   54085: result <= 12'b111100011111;
   54086: result <= 12'b111100011111;
   54087: result <= 12'b111100011111;
   54088: result <= 12'b111100011110;
   54089: result <= 12'b111100011110;
   54090: result <= 12'b111100011110;
   54091: result <= 12'b111100011110;
   54092: result <= 12'b111100011110;
   54093: result <= 12'b111100011110;
   54094: result <= 12'b111100011110;
   54095: result <= 12'b111100011110;
   54096: result <= 12'b111100011110;
   54097: result <= 12'b111100011110;
   54098: result <= 12'b111100011110;
   54099: result <= 12'b111100011101;
   54100: result <= 12'b111100011101;
   54101: result <= 12'b111100011101;
   54102: result <= 12'b111100011101;
   54103: result <= 12'b111100011101;
   54104: result <= 12'b111100011101;
   54105: result <= 12'b111100011101;
   54106: result <= 12'b111100011101;
   54107: result <= 12'b111100011101;
   54108: result <= 12'b111100011101;
   54109: result <= 12'b111100011101;
   54110: result <= 12'b111100011100;
   54111: result <= 12'b111100011100;
   54112: result <= 12'b111100011100;
   54113: result <= 12'b111100011100;
   54114: result <= 12'b111100011100;
   54115: result <= 12'b111100011100;
   54116: result <= 12'b111100011100;
   54117: result <= 12'b111100011100;
   54118: result <= 12'b111100011100;
   54119: result <= 12'b111100011100;
   54120: result <= 12'b111100011100;
   54121: result <= 12'b111100011011;
   54122: result <= 12'b111100011011;
   54123: result <= 12'b111100011011;
   54124: result <= 12'b111100011011;
   54125: result <= 12'b111100011011;
   54126: result <= 12'b111100011011;
   54127: result <= 12'b111100011011;
   54128: result <= 12'b111100011011;
   54129: result <= 12'b111100011011;
   54130: result <= 12'b111100011011;
   54131: result <= 12'b111100011011;
   54132: result <= 12'b111100011010;
   54133: result <= 12'b111100011010;
   54134: result <= 12'b111100011010;
   54135: result <= 12'b111100011010;
   54136: result <= 12'b111100011010;
   54137: result <= 12'b111100011010;
   54138: result <= 12'b111100011010;
   54139: result <= 12'b111100011010;
   54140: result <= 12'b111100011010;
   54141: result <= 12'b111100011010;
   54142: result <= 12'b111100011010;
   54143: result <= 12'b111100011001;
   54144: result <= 12'b111100011001;
   54145: result <= 12'b111100011001;
   54146: result <= 12'b111100011001;
   54147: result <= 12'b111100011001;
   54148: result <= 12'b111100011001;
   54149: result <= 12'b111100011001;
   54150: result <= 12'b111100011001;
   54151: result <= 12'b111100011001;
   54152: result <= 12'b111100011001;
   54153: result <= 12'b111100011001;
   54154: result <= 12'b111100011000;
   54155: result <= 12'b111100011000;
   54156: result <= 12'b111100011000;
   54157: result <= 12'b111100011000;
   54158: result <= 12'b111100011000;
   54159: result <= 12'b111100011000;
   54160: result <= 12'b111100011000;
   54161: result <= 12'b111100011000;
   54162: result <= 12'b111100011000;
   54163: result <= 12'b111100011000;
   54164: result <= 12'b111100011000;
   54165: result <= 12'b111100010111;
   54166: result <= 12'b111100010111;
   54167: result <= 12'b111100010111;
   54168: result <= 12'b111100010111;
   54169: result <= 12'b111100010111;
   54170: result <= 12'b111100010111;
   54171: result <= 12'b111100010111;
   54172: result <= 12'b111100010111;
   54173: result <= 12'b111100010111;
   54174: result <= 12'b111100010111;
   54175: result <= 12'b111100010111;
   54176: result <= 12'b111100010110;
   54177: result <= 12'b111100010110;
   54178: result <= 12'b111100010110;
   54179: result <= 12'b111100010110;
   54180: result <= 12'b111100010110;
   54181: result <= 12'b111100010110;
   54182: result <= 12'b111100010110;
   54183: result <= 12'b111100010110;
   54184: result <= 12'b111100010110;
   54185: result <= 12'b111100010110;
   54186: result <= 12'b111100010110;
   54187: result <= 12'b111100010101;
   54188: result <= 12'b111100010101;
   54189: result <= 12'b111100010101;
   54190: result <= 12'b111100010101;
   54191: result <= 12'b111100010101;
   54192: result <= 12'b111100010101;
   54193: result <= 12'b111100010101;
   54194: result <= 12'b111100010101;
   54195: result <= 12'b111100010101;
   54196: result <= 12'b111100010101;
   54197: result <= 12'b111100010101;
   54198: result <= 12'b111100010100;
   54199: result <= 12'b111100010100;
   54200: result <= 12'b111100010100;
   54201: result <= 12'b111100010100;
   54202: result <= 12'b111100010100;
   54203: result <= 12'b111100010100;
   54204: result <= 12'b111100010100;
   54205: result <= 12'b111100010100;
   54206: result <= 12'b111100010100;
   54207: result <= 12'b111100010100;
   54208: result <= 12'b111100010100;
   54209: result <= 12'b111100010011;
   54210: result <= 12'b111100010011;
   54211: result <= 12'b111100010011;
   54212: result <= 12'b111100010011;
   54213: result <= 12'b111100010011;
   54214: result <= 12'b111100010011;
   54215: result <= 12'b111100010011;
   54216: result <= 12'b111100010011;
   54217: result <= 12'b111100010011;
   54218: result <= 12'b111100010011;
   54219: result <= 12'b111100010011;
   54220: result <= 12'b111100010010;
   54221: result <= 12'b111100010010;
   54222: result <= 12'b111100010010;
   54223: result <= 12'b111100010010;
   54224: result <= 12'b111100010010;
   54225: result <= 12'b111100010010;
   54226: result <= 12'b111100010010;
   54227: result <= 12'b111100010010;
   54228: result <= 12'b111100010010;
   54229: result <= 12'b111100010010;
   54230: result <= 12'b111100010010;
   54231: result <= 12'b111100010001;
   54232: result <= 12'b111100010001;
   54233: result <= 12'b111100010001;
   54234: result <= 12'b111100010001;
   54235: result <= 12'b111100010001;
   54236: result <= 12'b111100010001;
   54237: result <= 12'b111100010001;
   54238: result <= 12'b111100010001;
   54239: result <= 12'b111100010001;
   54240: result <= 12'b111100010001;
   54241: result <= 12'b111100010001;
   54242: result <= 12'b111100010000;
   54243: result <= 12'b111100010000;
   54244: result <= 12'b111100010000;
   54245: result <= 12'b111100010000;
   54246: result <= 12'b111100010000;
   54247: result <= 12'b111100010000;
   54248: result <= 12'b111100010000;
   54249: result <= 12'b111100010000;
   54250: result <= 12'b111100010000;
   54251: result <= 12'b111100010000;
   54252: result <= 12'b111100010000;
   54253: result <= 12'b111100001111;
   54254: result <= 12'b111100001111;
   54255: result <= 12'b111100001111;
   54256: result <= 12'b111100001111;
   54257: result <= 12'b111100001111;
   54258: result <= 12'b111100001111;
   54259: result <= 12'b111100001111;
   54260: result <= 12'b111100001111;
   54261: result <= 12'b111100001111;
   54262: result <= 12'b111100001111;
   54263: result <= 12'b111100001111;
   54264: result <= 12'b111100001110;
   54265: result <= 12'b111100001110;
   54266: result <= 12'b111100001110;
   54267: result <= 12'b111100001110;
   54268: result <= 12'b111100001110;
   54269: result <= 12'b111100001110;
   54270: result <= 12'b111100001110;
   54271: result <= 12'b111100001110;
   54272: result <= 12'b111100001110;
   54273: result <= 12'b111100001110;
   54274: result <= 12'b111100001101;
   54275: result <= 12'b111100001101;
   54276: result <= 12'b111100001101;
   54277: result <= 12'b111100001101;
   54278: result <= 12'b111100001101;
   54279: result <= 12'b111100001101;
   54280: result <= 12'b111100001101;
   54281: result <= 12'b111100001101;
   54282: result <= 12'b111100001101;
   54283: result <= 12'b111100001101;
   54284: result <= 12'b111100001101;
   54285: result <= 12'b111100001100;
   54286: result <= 12'b111100001100;
   54287: result <= 12'b111100001100;
   54288: result <= 12'b111100001100;
   54289: result <= 12'b111100001100;
   54290: result <= 12'b111100001100;
   54291: result <= 12'b111100001100;
   54292: result <= 12'b111100001100;
   54293: result <= 12'b111100001100;
   54294: result <= 12'b111100001100;
   54295: result <= 12'b111100001100;
   54296: result <= 12'b111100001011;
   54297: result <= 12'b111100001011;
   54298: result <= 12'b111100001011;
   54299: result <= 12'b111100001011;
   54300: result <= 12'b111100001011;
   54301: result <= 12'b111100001011;
   54302: result <= 12'b111100001011;
   54303: result <= 12'b111100001011;
   54304: result <= 12'b111100001011;
   54305: result <= 12'b111100001011;
   54306: result <= 12'b111100001011;
   54307: result <= 12'b111100001010;
   54308: result <= 12'b111100001010;
   54309: result <= 12'b111100001010;
   54310: result <= 12'b111100001010;
   54311: result <= 12'b111100001010;
   54312: result <= 12'b111100001010;
   54313: result <= 12'b111100001010;
   54314: result <= 12'b111100001010;
   54315: result <= 12'b111100001010;
   54316: result <= 12'b111100001010;
   54317: result <= 12'b111100001001;
   54318: result <= 12'b111100001001;
   54319: result <= 12'b111100001001;
   54320: result <= 12'b111100001001;
   54321: result <= 12'b111100001001;
   54322: result <= 12'b111100001001;
   54323: result <= 12'b111100001001;
   54324: result <= 12'b111100001001;
   54325: result <= 12'b111100001001;
   54326: result <= 12'b111100001001;
   54327: result <= 12'b111100001001;
   54328: result <= 12'b111100001000;
   54329: result <= 12'b111100001000;
   54330: result <= 12'b111100001000;
   54331: result <= 12'b111100001000;
   54332: result <= 12'b111100001000;
   54333: result <= 12'b111100001000;
   54334: result <= 12'b111100001000;
   54335: result <= 12'b111100001000;
   54336: result <= 12'b111100001000;
   54337: result <= 12'b111100001000;
   54338: result <= 12'b111100001000;
   54339: result <= 12'b111100000111;
   54340: result <= 12'b111100000111;
   54341: result <= 12'b111100000111;
   54342: result <= 12'b111100000111;
   54343: result <= 12'b111100000111;
   54344: result <= 12'b111100000111;
   54345: result <= 12'b111100000111;
   54346: result <= 12'b111100000111;
   54347: result <= 12'b111100000111;
   54348: result <= 12'b111100000111;
   54349: result <= 12'b111100000110;
   54350: result <= 12'b111100000110;
   54351: result <= 12'b111100000110;
   54352: result <= 12'b111100000110;
   54353: result <= 12'b111100000110;
   54354: result <= 12'b111100000110;
   54355: result <= 12'b111100000110;
   54356: result <= 12'b111100000110;
   54357: result <= 12'b111100000110;
   54358: result <= 12'b111100000110;
   54359: result <= 12'b111100000110;
   54360: result <= 12'b111100000101;
   54361: result <= 12'b111100000101;
   54362: result <= 12'b111100000101;
   54363: result <= 12'b111100000101;
   54364: result <= 12'b111100000101;
   54365: result <= 12'b111100000101;
   54366: result <= 12'b111100000101;
   54367: result <= 12'b111100000101;
   54368: result <= 12'b111100000101;
   54369: result <= 12'b111100000101;
   54370: result <= 12'b111100000101;
   54371: result <= 12'b111100000100;
   54372: result <= 12'b111100000100;
   54373: result <= 12'b111100000100;
   54374: result <= 12'b111100000100;
   54375: result <= 12'b111100000100;
   54376: result <= 12'b111100000100;
   54377: result <= 12'b111100000100;
   54378: result <= 12'b111100000100;
   54379: result <= 12'b111100000100;
   54380: result <= 12'b111100000100;
   54381: result <= 12'b111100000011;
   54382: result <= 12'b111100000011;
   54383: result <= 12'b111100000011;
   54384: result <= 12'b111100000011;
   54385: result <= 12'b111100000011;
   54386: result <= 12'b111100000011;
   54387: result <= 12'b111100000011;
   54388: result <= 12'b111100000011;
   54389: result <= 12'b111100000011;
   54390: result <= 12'b111100000011;
   54391: result <= 12'b111100000011;
   54392: result <= 12'b111100000010;
   54393: result <= 12'b111100000010;
   54394: result <= 12'b111100000010;
   54395: result <= 12'b111100000010;
   54396: result <= 12'b111100000010;
   54397: result <= 12'b111100000010;
   54398: result <= 12'b111100000010;
   54399: result <= 12'b111100000010;
   54400: result <= 12'b111100000010;
   54401: result <= 12'b111100000010;
   54402: result <= 12'b111100000010;
   54403: result <= 12'b111100000001;
   54404: result <= 12'b111100000001;
   54405: result <= 12'b111100000001;
   54406: result <= 12'b111100000001;
   54407: result <= 12'b111100000001;
   54408: result <= 12'b111100000001;
   54409: result <= 12'b111100000001;
   54410: result <= 12'b111100000001;
   54411: result <= 12'b111100000001;
   54412: result <= 12'b111100000001;
   54413: result <= 12'b111100000000;
   54414: result <= 12'b111100000000;
   54415: result <= 12'b111100000000;
   54416: result <= 12'b111100000000;
   54417: result <= 12'b111100000000;
   54418: result <= 12'b111100000000;
   54419: result <= 12'b111100000000;
   54420: result <= 12'b111100000000;
   54421: result <= 12'b111100000000;
   54422: result <= 12'b111100000000;
   54423: result <= 12'b111100000000;
   54424: result <= 12'b111011111111;
   54425: result <= 12'b111011111111;
   54426: result <= 12'b111011111111;
   54427: result <= 12'b111011111111;
   54428: result <= 12'b111011111111;
   54429: result <= 12'b111011111111;
   54430: result <= 12'b111011111111;
   54431: result <= 12'b111011111111;
   54432: result <= 12'b111011111111;
   54433: result <= 12'b111011111111;
   54434: result <= 12'b111011111110;
   54435: result <= 12'b111011111110;
   54436: result <= 12'b111011111110;
   54437: result <= 12'b111011111110;
   54438: result <= 12'b111011111110;
   54439: result <= 12'b111011111110;
   54440: result <= 12'b111011111110;
   54441: result <= 12'b111011111110;
   54442: result <= 12'b111011111110;
   54443: result <= 12'b111011111110;
   54444: result <= 12'b111011111110;
   54445: result <= 12'b111011111101;
   54446: result <= 12'b111011111101;
   54447: result <= 12'b111011111101;
   54448: result <= 12'b111011111101;
   54449: result <= 12'b111011111101;
   54450: result <= 12'b111011111101;
   54451: result <= 12'b111011111101;
   54452: result <= 12'b111011111101;
   54453: result <= 12'b111011111101;
   54454: result <= 12'b111011111101;
   54455: result <= 12'b111011111100;
   54456: result <= 12'b111011111100;
   54457: result <= 12'b111011111100;
   54458: result <= 12'b111011111100;
   54459: result <= 12'b111011111100;
   54460: result <= 12'b111011111100;
   54461: result <= 12'b111011111100;
   54462: result <= 12'b111011111100;
   54463: result <= 12'b111011111100;
   54464: result <= 12'b111011111100;
   54465: result <= 12'b111011111100;
   54466: result <= 12'b111011111011;
   54467: result <= 12'b111011111011;
   54468: result <= 12'b111011111011;
   54469: result <= 12'b111011111011;
   54470: result <= 12'b111011111011;
   54471: result <= 12'b111011111011;
   54472: result <= 12'b111011111011;
   54473: result <= 12'b111011111011;
   54474: result <= 12'b111011111011;
   54475: result <= 12'b111011111011;
   54476: result <= 12'b111011111010;
   54477: result <= 12'b111011111010;
   54478: result <= 12'b111011111010;
   54479: result <= 12'b111011111010;
   54480: result <= 12'b111011111010;
   54481: result <= 12'b111011111010;
   54482: result <= 12'b111011111010;
   54483: result <= 12'b111011111010;
   54484: result <= 12'b111011111010;
   54485: result <= 12'b111011111010;
   54486: result <= 12'b111011111001;
   54487: result <= 12'b111011111001;
   54488: result <= 12'b111011111001;
   54489: result <= 12'b111011111001;
   54490: result <= 12'b111011111001;
   54491: result <= 12'b111011111001;
   54492: result <= 12'b111011111001;
   54493: result <= 12'b111011111001;
   54494: result <= 12'b111011111001;
   54495: result <= 12'b111011111001;
   54496: result <= 12'b111011111001;
   54497: result <= 12'b111011111000;
   54498: result <= 12'b111011111000;
   54499: result <= 12'b111011111000;
   54500: result <= 12'b111011111000;
   54501: result <= 12'b111011111000;
   54502: result <= 12'b111011111000;
   54503: result <= 12'b111011111000;
   54504: result <= 12'b111011111000;
   54505: result <= 12'b111011111000;
   54506: result <= 12'b111011111000;
   54507: result <= 12'b111011110111;
   54508: result <= 12'b111011110111;
   54509: result <= 12'b111011110111;
   54510: result <= 12'b111011110111;
   54511: result <= 12'b111011110111;
   54512: result <= 12'b111011110111;
   54513: result <= 12'b111011110111;
   54514: result <= 12'b111011110111;
   54515: result <= 12'b111011110111;
   54516: result <= 12'b111011110111;
   54517: result <= 12'b111011110111;
   54518: result <= 12'b111011110110;
   54519: result <= 12'b111011110110;
   54520: result <= 12'b111011110110;
   54521: result <= 12'b111011110110;
   54522: result <= 12'b111011110110;
   54523: result <= 12'b111011110110;
   54524: result <= 12'b111011110110;
   54525: result <= 12'b111011110110;
   54526: result <= 12'b111011110110;
   54527: result <= 12'b111011110110;
   54528: result <= 12'b111011110101;
   54529: result <= 12'b111011110101;
   54530: result <= 12'b111011110101;
   54531: result <= 12'b111011110101;
   54532: result <= 12'b111011110101;
   54533: result <= 12'b111011110101;
   54534: result <= 12'b111011110101;
   54535: result <= 12'b111011110101;
   54536: result <= 12'b111011110101;
   54537: result <= 12'b111011110101;
   54538: result <= 12'b111011110100;
   54539: result <= 12'b111011110100;
   54540: result <= 12'b111011110100;
   54541: result <= 12'b111011110100;
   54542: result <= 12'b111011110100;
   54543: result <= 12'b111011110100;
   54544: result <= 12'b111011110100;
   54545: result <= 12'b111011110100;
   54546: result <= 12'b111011110100;
   54547: result <= 12'b111011110100;
   54548: result <= 12'b111011110011;
   54549: result <= 12'b111011110011;
   54550: result <= 12'b111011110011;
   54551: result <= 12'b111011110011;
   54552: result <= 12'b111011110011;
   54553: result <= 12'b111011110011;
   54554: result <= 12'b111011110011;
   54555: result <= 12'b111011110011;
   54556: result <= 12'b111011110011;
   54557: result <= 12'b111011110011;
   54558: result <= 12'b111011110011;
   54559: result <= 12'b111011110010;
   54560: result <= 12'b111011110010;
   54561: result <= 12'b111011110010;
   54562: result <= 12'b111011110010;
   54563: result <= 12'b111011110010;
   54564: result <= 12'b111011110010;
   54565: result <= 12'b111011110010;
   54566: result <= 12'b111011110010;
   54567: result <= 12'b111011110010;
   54568: result <= 12'b111011110010;
   54569: result <= 12'b111011110001;
   54570: result <= 12'b111011110001;
   54571: result <= 12'b111011110001;
   54572: result <= 12'b111011110001;
   54573: result <= 12'b111011110001;
   54574: result <= 12'b111011110001;
   54575: result <= 12'b111011110001;
   54576: result <= 12'b111011110001;
   54577: result <= 12'b111011110001;
   54578: result <= 12'b111011110001;
   54579: result <= 12'b111011110000;
   54580: result <= 12'b111011110000;
   54581: result <= 12'b111011110000;
   54582: result <= 12'b111011110000;
   54583: result <= 12'b111011110000;
   54584: result <= 12'b111011110000;
   54585: result <= 12'b111011110000;
   54586: result <= 12'b111011110000;
   54587: result <= 12'b111011110000;
   54588: result <= 12'b111011110000;
   54589: result <= 12'b111011110000;
   54590: result <= 12'b111011101111;
   54591: result <= 12'b111011101111;
   54592: result <= 12'b111011101111;
   54593: result <= 12'b111011101111;
   54594: result <= 12'b111011101111;
   54595: result <= 12'b111011101111;
   54596: result <= 12'b111011101111;
   54597: result <= 12'b111011101111;
   54598: result <= 12'b111011101111;
   54599: result <= 12'b111011101111;
   54600: result <= 12'b111011101110;
   54601: result <= 12'b111011101110;
   54602: result <= 12'b111011101110;
   54603: result <= 12'b111011101110;
   54604: result <= 12'b111011101110;
   54605: result <= 12'b111011101110;
   54606: result <= 12'b111011101110;
   54607: result <= 12'b111011101110;
   54608: result <= 12'b111011101110;
   54609: result <= 12'b111011101110;
   54610: result <= 12'b111011101101;
   54611: result <= 12'b111011101101;
   54612: result <= 12'b111011101101;
   54613: result <= 12'b111011101101;
   54614: result <= 12'b111011101101;
   54615: result <= 12'b111011101101;
   54616: result <= 12'b111011101101;
   54617: result <= 12'b111011101101;
   54618: result <= 12'b111011101101;
   54619: result <= 12'b111011101101;
   54620: result <= 12'b111011101100;
   54621: result <= 12'b111011101100;
   54622: result <= 12'b111011101100;
   54623: result <= 12'b111011101100;
   54624: result <= 12'b111011101100;
   54625: result <= 12'b111011101100;
   54626: result <= 12'b111011101100;
   54627: result <= 12'b111011101100;
   54628: result <= 12'b111011101100;
   54629: result <= 12'b111011101100;
   54630: result <= 12'b111011101011;
   54631: result <= 12'b111011101011;
   54632: result <= 12'b111011101011;
   54633: result <= 12'b111011101011;
   54634: result <= 12'b111011101011;
   54635: result <= 12'b111011101011;
   54636: result <= 12'b111011101011;
   54637: result <= 12'b111011101011;
   54638: result <= 12'b111011101011;
   54639: result <= 12'b111011101011;
   54640: result <= 12'b111011101010;
   54641: result <= 12'b111011101010;
   54642: result <= 12'b111011101010;
   54643: result <= 12'b111011101010;
   54644: result <= 12'b111011101010;
   54645: result <= 12'b111011101010;
   54646: result <= 12'b111011101010;
   54647: result <= 12'b111011101010;
   54648: result <= 12'b111011101010;
   54649: result <= 12'b111011101010;
   54650: result <= 12'b111011101010;
   54651: result <= 12'b111011101001;
   54652: result <= 12'b111011101001;
   54653: result <= 12'b111011101001;
   54654: result <= 12'b111011101001;
   54655: result <= 12'b111011101001;
   54656: result <= 12'b111011101001;
   54657: result <= 12'b111011101001;
   54658: result <= 12'b111011101001;
   54659: result <= 12'b111011101001;
   54660: result <= 12'b111011101001;
   54661: result <= 12'b111011101000;
   54662: result <= 12'b111011101000;
   54663: result <= 12'b111011101000;
   54664: result <= 12'b111011101000;
   54665: result <= 12'b111011101000;
   54666: result <= 12'b111011101000;
   54667: result <= 12'b111011101000;
   54668: result <= 12'b111011101000;
   54669: result <= 12'b111011101000;
   54670: result <= 12'b111011101000;
   54671: result <= 12'b111011100111;
   54672: result <= 12'b111011100111;
   54673: result <= 12'b111011100111;
   54674: result <= 12'b111011100111;
   54675: result <= 12'b111011100111;
   54676: result <= 12'b111011100111;
   54677: result <= 12'b111011100111;
   54678: result <= 12'b111011100111;
   54679: result <= 12'b111011100111;
   54680: result <= 12'b111011100111;
   54681: result <= 12'b111011100110;
   54682: result <= 12'b111011100110;
   54683: result <= 12'b111011100110;
   54684: result <= 12'b111011100110;
   54685: result <= 12'b111011100110;
   54686: result <= 12'b111011100110;
   54687: result <= 12'b111011100110;
   54688: result <= 12'b111011100110;
   54689: result <= 12'b111011100110;
   54690: result <= 12'b111011100110;
   54691: result <= 12'b111011100101;
   54692: result <= 12'b111011100101;
   54693: result <= 12'b111011100101;
   54694: result <= 12'b111011100101;
   54695: result <= 12'b111011100101;
   54696: result <= 12'b111011100101;
   54697: result <= 12'b111011100101;
   54698: result <= 12'b111011100101;
   54699: result <= 12'b111011100101;
   54700: result <= 12'b111011100101;
   54701: result <= 12'b111011100100;
   54702: result <= 12'b111011100100;
   54703: result <= 12'b111011100100;
   54704: result <= 12'b111011100100;
   54705: result <= 12'b111011100100;
   54706: result <= 12'b111011100100;
   54707: result <= 12'b111011100100;
   54708: result <= 12'b111011100100;
   54709: result <= 12'b111011100100;
   54710: result <= 12'b111011100100;
   54711: result <= 12'b111011100011;
   54712: result <= 12'b111011100011;
   54713: result <= 12'b111011100011;
   54714: result <= 12'b111011100011;
   54715: result <= 12'b111011100011;
   54716: result <= 12'b111011100011;
   54717: result <= 12'b111011100011;
   54718: result <= 12'b111011100011;
   54719: result <= 12'b111011100011;
   54720: result <= 12'b111011100011;
   54721: result <= 12'b111011100010;
   54722: result <= 12'b111011100010;
   54723: result <= 12'b111011100010;
   54724: result <= 12'b111011100010;
   54725: result <= 12'b111011100010;
   54726: result <= 12'b111011100010;
   54727: result <= 12'b111011100010;
   54728: result <= 12'b111011100010;
   54729: result <= 12'b111011100010;
   54730: result <= 12'b111011100010;
   54731: result <= 12'b111011100001;
   54732: result <= 12'b111011100001;
   54733: result <= 12'b111011100001;
   54734: result <= 12'b111011100001;
   54735: result <= 12'b111011100001;
   54736: result <= 12'b111011100001;
   54737: result <= 12'b111011100001;
   54738: result <= 12'b111011100001;
   54739: result <= 12'b111011100001;
   54740: result <= 12'b111011100001;
   54741: result <= 12'b111011100000;
   54742: result <= 12'b111011100000;
   54743: result <= 12'b111011100000;
   54744: result <= 12'b111011100000;
   54745: result <= 12'b111011100000;
   54746: result <= 12'b111011100000;
   54747: result <= 12'b111011100000;
   54748: result <= 12'b111011100000;
   54749: result <= 12'b111011100000;
   54750: result <= 12'b111011100000;
   54751: result <= 12'b111011011111;
   54752: result <= 12'b111011011111;
   54753: result <= 12'b111011011111;
   54754: result <= 12'b111011011111;
   54755: result <= 12'b111011011111;
   54756: result <= 12'b111011011111;
   54757: result <= 12'b111011011111;
   54758: result <= 12'b111011011111;
   54759: result <= 12'b111011011111;
   54760: result <= 12'b111011011111;
   54761: result <= 12'b111011011110;
   54762: result <= 12'b111011011110;
   54763: result <= 12'b111011011110;
   54764: result <= 12'b111011011110;
   54765: result <= 12'b111011011110;
   54766: result <= 12'b111011011110;
   54767: result <= 12'b111011011110;
   54768: result <= 12'b111011011110;
   54769: result <= 12'b111011011110;
   54770: result <= 12'b111011011110;
   54771: result <= 12'b111011011101;
   54772: result <= 12'b111011011101;
   54773: result <= 12'b111011011101;
   54774: result <= 12'b111011011101;
   54775: result <= 12'b111011011101;
   54776: result <= 12'b111011011101;
   54777: result <= 12'b111011011101;
   54778: result <= 12'b111011011101;
   54779: result <= 12'b111011011101;
   54780: result <= 12'b111011011101;
   54781: result <= 12'b111011011100;
   54782: result <= 12'b111011011100;
   54783: result <= 12'b111011011100;
   54784: result <= 12'b111011011100;
   54785: result <= 12'b111011011100;
   54786: result <= 12'b111011011100;
   54787: result <= 12'b111011011100;
   54788: result <= 12'b111011011100;
   54789: result <= 12'b111011011100;
   54790: result <= 12'b111011011100;
   54791: result <= 12'b111011011011;
   54792: result <= 12'b111011011011;
   54793: result <= 12'b111011011011;
   54794: result <= 12'b111011011011;
   54795: result <= 12'b111011011011;
   54796: result <= 12'b111011011011;
   54797: result <= 12'b111011011011;
   54798: result <= 12'b111011011011;
   54799: result <= 12'b111011011011;
   54800: result <= 12'b111011011011;
   54801: result <= 12'b111011011010;
   54802: result <= 12'b111011011010;
   54803: result <= 12'b111011011010;
   54804: result <= 12'b111011011010;
   54805: result <= 12'b111011011010;
   54806: result <= 12'b111011011010;
   54807: result <= 12'b111011011010;
   54808: result <= 12'b111011011010;
   54809: result <= 12'b111011011010;
   54810: result <= 12'b111011011001;
   54811: result <= 12'b111011011001;
   54812: result <= 12'b111011011001;
   54813: result <= 12'b111011011001;
   54814: result <= 12'b111011011001;
   54815: result <= 12'b111011011001;
   54816: result <= 12'b111011011001;
   54817: result <= 12'b111011011001;
   54818: result <= 12'b111011011001;
   54819: result <= 12'b111011011001;
   54820: result <= 12'b111011011000;
   54821: result <= 12'b111011011000;
   54822: result <= 12'b111011011000;
   54823: result <= 12'b111011011000;
   54824: result <= 12'b111011011000;
   54825: result <= 12'b111011011000;
   54826: result <= 12'b111011011000;
   54827: result <= 12'b111011011000;
   54828: result <= 12'b111011011000;
   54829: result <= 12'b111011011000;
   54830: result <= 12'b111011010111;
   54831: result <= 12'b111011010111;
   54832: result <= 12'b111011010111;
   54833: result <= 12'b111011010111;
   54834: result <= 12'b111011010111;
   54835: result <= 12'b111011010111;
   54836: result <= 12'b111011010111;
   54837: result <= 12'b111011010111;
   54838: result <= 12'b111011010111;
   54839: result <= 12'b111011010111;
   54840: result <= 12'b111011010110;
   54841: result <= 12'b111011010110;
   54842: result <= 12'b111011010110;
   54843: result <= 12'b111011010110;
   54844: result <= 12'b111011010110;
   54845: result <= 12'b111011010110;
   54846: result <= 12'b111011010110;
   54847: result <= 12'b111011010110;
   54848: result <= 12'b111011010110;
   54849: result <= 12'b111011010110;
   54850: result <= 12'b111011010101;
   54851: result <= 12'b111011010101;
   54852: result <= 12'b111011010101;
   54853: result <= 12'b111011010101;
   54854: result <= 12'b111011010101;
   54855: result <= 12'b111011010101;
   54856: result <= 12'b111011010101;
   54857: result <= 12'b111011010101;
   54858: result <= 12'b111011010101;
   54859: result <= 12'b111011010101;
   54860: result <= 12'b111011010100;
   54861: result <= 12'b111011010100;
   54862: result <= 12'b111011010100;
   54863: result <= 12'b111011010100;
   54864: result <= 12'b111011010100;
   54865: result <= 12'b111011010100;
   54866: result <= 12'b111011010100;
   54867: result <= 12'b111011010100;
   54868: result <= 12'b111011010100;
   54869: result <= 12'b111011010011;
   54870: result <= 12'b111011010011;
   54871: result <= 12'b111011010011;
   54872: result <= 12'b111011010011;
   54873: result <= 12'b111011010011;
   54874: result <= 12'b111011010011;
   54875: result <= 12'b111011010011;
   54876: result <= 12'b111011010011;
   54877: result <= 12'b111011010011;
   54878: result <= 12'b111011010011;
   54879: result <= 12'b111011010010;
   54880: result <= 12'b111011010010;
   54881: result <= 12'b111011010010;
   54882: result <= 12'b111011010010;
   54883: result <= 12'b111011010010;
   54884: result <= 12'b111011010010;
   54885: result <= 12'b111011010010;
   54886: result <= 12'b111011010010;
   54887: result <= 12'b111011010010;
   54888: result <= 12'b111011010010;
   54889: result <= 12'b111011010001;
   54890: result <= 12'b111011010001;
   54891: result <= 12'b111011010001;
   54892: result <= 12'b111011010001;
   54893: result <= 12'b111011010001;
   54894: result <= 12'b111011010001;
   54895: result <= 12'b111011010001;
   54896: result <= 12'b111011010001;
   54897: result <= 12'b111011010001;
   54898: result <= 12'b111011010001;
   54899: result <= 12'b111011010000;
   54900: result <= 12'b111011010000;
   54901: result <= 12'b111011010000;
   54902: result <= 12'b111011010000;
   54903: result <= 12'b111011010000;
   54904: result <= 12'b111011010000;
   54905: result <= 12'b111011010000;
   54906: result <= 12'b111011010000;
   54907: result <= 12'b111011010000;
   54908: result <= 12'b111011001111;
   54909: result <= 12'b111011001111;
   54910: result <= 12'b111011001111;
   54911: result <= 12'b111011001111;
   54912: result <= 12'b111011001111;
   54913: result <= 12'b111011001111;
   54914: result <= 12'b111011001111;
   54915: result <= 12'b111011001111;
   54916: result <= 12'b111011001111;
   54917: result <= 12'b111011001111;
   54918: result <= 12'b111011001110;
   54919: result <= 12'b111011001110;
   54920: result <= 12'b111011001110;
   54921: result <= 12'b111011001110;
   54922: result <= 12'b111011001110;
   54923: result <= 12'b111011001110;
   54924: result <= 12'b111011001110;
   54925: result <= 12'b111011001110;
   54926: result <= 12'b111011001110;
   54927: result <= 12'b111011001110;
   54928: result <= 12'b111011001101;
   54929: result <= 12'b111011001101;
   54930: result <= 12'b111011001101;
   54931: result <= 12'b111011001101;
   54932: result <= 12'b111011001101;
   54933: result <= 12'b111011001101;
   54934: result <= 12'b111011001101;
   54935: result <= 12'b111011001101;
   54936: result <= 12'b111011001101;
   54937: result <= 12'b111011001100;
   54938: result <= 12'b111011001100;
   54939: result <= 12'b111011001100;
   54940: result <= 12'b111011001100;
   54941: result <= 12'b111011001100;
   54942: result <= 12'b111011001100;
   54943: result <= 12'b111011001100;
   54944: result <= 12'b111011001100;
   54945: result <= 12'b111011001100;
   54946: result <= 12'b111011001100;
   54947: result <= 12'b111011001011;
   54948: result <= 12'b111011001011;
   54949: result <= 12'b111011001011;
   54950: result <= 12'b111011001011;
   54951: result <= 12'b111011001011;
   54952: result <= 12'b111011001011;
   54953: result <= 12'b111011001011;
   54954: result <= 12'b111011001011;
   54955: result <= 12'b111011001011;
   54956: result <= 12'b111011001011;
   54957: result <= 12'b111011001010;
   54958: result <= 12'b111011001010;
   54959: result <= 12'b111011001010;
   54960: result <= 12'b111011001010;
   54961: result <= 12'b111011001010;
   54962: result <= 12'b111011001010;
   54963: result <= 12'b111011001010;
   54964: result <= 12'b111011001010;
   54965: result <= 12'b111011001010;
   54966: result <= 12'b111011001001;
   54967: result <= 12'b111011001001;
   54968: result <= 12'b111011001001;
   54969: result <= 12'b111011001001;
   54970: result <= 12'b111011001001;
   54971: result <= 12'b111011001001;
   54972: result <= 12'b111011001001;
   54973: result <= 12'b111011001001;
   54974: result <= 12'b111011001001;
   54975: result <= 12'b111011001001;
   54976: result <= 12'b111011001000;
   54977: result <= 12'b111011001000;
   54978: result <= 12'b111011001000;
   54979: result <= 12'b111011001000;
   54980: result <= 12'b111011001000;
   54981: result <= 12'b111011001000;
   54982: result <= 12'b111011001000;
   54983: result <= 12'b111011001000;
   54984: result <= 12'b111011001000;
   54985: result <= 12'b111011001000;
   54986: result <= 12'b111011000111;
   54987: result <= 12'b111011000111;
   54988: result <= 12'b111011000111;
   54989: result <= 12'b111011000111;
   54990: result <= 12'b111011000111;
   54991: result <= 12'b111011000111;
   54992: result <= 12'b111011000111;
   54993: result <= 12'b111011000111;
   54994: result <= 12'b111011000111;
   54995: result <= 12'b111011000110;
   54996: result <= 12'b111011000110;
   54997: result <= 12'b111011000110;
   54998: result <= 12'b111011000110;
   54999: result <= 12'b111011000110;
   55000: result <= 12'b111011000110;
   55001: result <= 12'b111011000110;
   55002: result <= 12'b111011000110;
   55003: result <= 12'b111011000110;
   55004: result <= 12'b111011000110;
   55005: result <= 12'b111011000101;
   55006: result <= 12'b111011000101;
   55007: result <= 12'b111011000101;
   55008: result <= 12'b111011000101;
   55009: result <= 12'b111011000101;
   55010: result <= 12'b111011000101;
   55011: result <= 12'b111011000101;
   55012: result <= 12'b111011000101;
   55013: result <= 12'b111011000101;
   55014: result <= 12'b111011000100;
   55015: result <= 12'b111011000100;
   55016: result <= 12'b111011000100;
   55017: result <= 12'b111011000100;
   55018: result <= 12'b111011000100;
   55019: result <= 12'b111011000100;
   55020: result <= 12'b111011000100;
   55021: result <= 12'b111011000100;
   55022: result <= 12'b111011000100;
   55023: result <= 12'b111011000100;
   55024: result <= 12'b111011000011;
   55025: result <= 12'b111011000011;
   55026: result <= 12'b111011000011;
   55027: result <= 12'b111011000011;
   55028: result <= 12'b111011000011;
   55029: result <= 12'b111011000011;
   55030: result <= 12'b111011000011;
   55031: result <= 12'b111011000011;
   55032: result <= 12'b111011000011;
   55033: result <= 12'b111011000010;
   55034: result <= 12'b111011000010;
   55035: result <= 12'b111011000010;
   55036: result <= 12'b111011000010;
   55037: result <= 12'b111011000010;
   55038: result <= 12'b111011000010;
   55039: result <= 12'b111011000010;
   55040: result <= 12'b111011000010;
   55041: result <= 12'b111011000010;
   55042: result <= 12'b111011000010;
   55043: result <= 12'b111011000001;
   55044: result <= 12'b111011000001;
   55045: result <= 12'b111011000001;
   55046: result <= 12'b111011000001;
   55047: result <= 12'b111011000001;
   55048: result <= 12'b111011000001;
   55049: result <= 12'b111011000001;
   55050: result <= 12'b111011000001;
   55051: result <= 12'b111011000001;
   55052: result <= 12'b111011000000;
   55053: result <= 12'b111011000000;
   55054: result <= 12'b111011000000;
   55055: result <= 12'b111011000000;
   55056: result <= 12'b111011000000;
   55057: result <= 12'b111011000000;
   55058: result <= 12'b111011000000;
   55059: result <= 12'b111011000000;
   55060: result <= 12'b111011000000;
   55061: result <= 12'b111011000000;
   55062: result <= 12'b111010111111;
   55063: result <= 12'b111010111111;
   55064: result <= 12'b111010111111;
   55065: result <= 12'b111010111111;
   55066: result <= 12'b111010111111;
   55067: result <= 12'b111010111111;
   55068: result <= 12'b111010111111;
   55069: result <= 12'b111010111111;
   55070: result <= 12'b111010111111;
   55071: result <= 12'b111010111110;
   55072: result <= 12'b111010111110;
   55073: result <= 12'b111010111110;
   55074: result <= 12'b111010111110;
   55075: result <= 12'b111010111110;
   55076: result <= 12'b111010111110;
   55077: result <= 12'b111010111110;
   55078: result <= 12'b111010111110;
   55079: result <= 12'b111010111110;
   55080: result <= 12'b111010111110;
   55081: result <= 12'b111010111101;
   55082: result <= 12'b111010111101;
   55083: result <= 12'b111010111101;
   55084: result <= 12'b111010111101;
   55085: result <= 12'b111010111101;
   55086: result <= 12'b111010111101;
   55087: result <= 12'b111010111101;
   55088: result <= 12'b111010111101;
   55089: result <= 12'b111010111101;
   55090: result <= 12'b111010111100;
   55091: result <= 12'b111010111100;
   55092: result <= 12'b111010111100;
   55093: result <= 12'b111010111100;
   55094: result <= 12'b111010111100;
   55095: result <= 12'b111010111100;
   55096: result <= 12'b111010111100;
   55097: result <= 12'b111010111100;
   55098: result <= 12'b111010111100;
   55099: result <= 12'b111010111100;
   55100: result <= 12'b111010111011;
   55101: result <= 12'b111010111011;
   55102: result <= 12'b111010111011;
   55103: result <= 12'b111010111011;
   55104: result <= 12'b111010111011;
   55105: result <= 12'b111010111011;
   55106: result <= 12'b111010111011;
   55107: result <= 12'b111010111011;
   55108: result <= 12'b111010111011;
   55109: result <= 12'b111010111010;
   55110: result <= 12'b111010111010;
   55111: result <= 12'b111010111010;
   55112: result <= 12'b111010111010;
   55113: result <= 12'b111010111010;
   55114: result <= 12'b111010111010;
   55115: result <= 12'b111010111010;
   55116: result <= 12'b111010111010;
   55117: result <= 12'b111010111010;
   55118: result <= 12'b111010111010;
   55119: result <= 12'b111010111001;
   55120: result <= 12'b111010111001;
   55121: result <= 12'b111010111001;
   55122: result <= 12'b111010111001;
   55123: result <= 12'b111010111001;
   55124: result <= 12'b111010111001;
   55125: result <= 12'b111010111001;
   55126: result <= 12'b111010111001;
   55127: result <= 12'b111010111001;
   55128: result <= 12'b111010111000;
   55129: result <= 12'b111010111000;
   55130: result <= 12'b111010111000;
   55131: result <= 12'b111010111000;
   55132: result <= 12'b111010111000;
   55133: result <= 12'b111010111000;
   55134: result <= 12'b111010111000;
   55135: result <= 12'b111010111000;
   55136: result <= 12'b111010111000;
   55137: result <= 12'b111010110111;
   55138: result <= 12'b111010110111;
   55139: result <= 12'b111010110111;
   55140: result <= 12'b111010110111;
   55141: result <= 12'b111010110111;
   55142: result <= 12'b111010110111;
   55143: result <= 12'b111010110111;
   55144: result <= 12'b111010110111;
   55145: result <= 12'b111010110111;
   55146: result <= 12'b111010110111;
   55147: result <= 12'b111010110110;
   55148: result <= 12'b111010110110;
   55149: result <= 12'b111010110110;
   55150: result <= 12'b111010110110;
   55151: result <= 12'b111010110110;
   55152: result <= 12'b111010110110;
   55153: result <= 12'b111010110110;
   55154: result <= 12'b111010110110;
   55155: result <= 12'b111010110110;
   55156: result <= 12'b111010110101;
   55157: result <= 12'b111010110101;
   55158: result <= 12'b111010110101;
   55159: result <= 12'b111010110101;
   55160: result <= 12'b111010110101;
   55161: result <= 12'b111010110101;
   55162: result <= 12'b111010110101;
   55163: result <= 12'b111010110101;
   55164: result <= 12'b111010110101;
   55165: result <= 12'b111010110101;
   55166: result <= 12'b111010110100;
   55167: result <= 12'b111010110100;
   55168: result <= 12'b111010110100;
   55169: result <= 12'b111010110100;
   55170: result <= 12'b111010110100;
   55171: result <= 12'b111010110100;
   55172: result <= 12'b111010110100;
   55173: result <= 12'b111010110100;
   55174: result <= 12'b111010110100;
   55175: result <= 12'b111010110011;
   55176: result <= 12'b111010110011;
   55177: result <= 12'b111010110011;
   55178: result <= 12'b111010110011;
   55179: result <= 12'b111010110011;
   55180: result <= 12'b111010110011;
   55181: result <= 12'b111010110011;
   55182: result <= 12'b111010110011;
   55183: result <= 12'b111010110011;
   55184: result <= 12'b111010110010;
   55185: result <= 12'b111010110010;
   55186: result <= 12'b111010110010;
   55187: result <= 12'b111010110010;
   55188: result <= 12'b111010110010;
   55189: result <= 12'b111010110010;
   55190: result <= 12'b111010110010;
   55191: result <= 12'b111010110010;
   55192: result <= 12'b111010110010;
   55193: result <= 12'b111010110010;
   55194: result <= 12'b111010110001;
   55195: result <= 12'b111010110001;
   55196: result <= 12'b111010110001;
   55197: result <= 12'b111010110001;
   55198: result <= 12'b111010110001;
   55199: result <= 12'b111010110001;
   55200: result <= 12'b111010110001;
   55201: result <= 12'b111010110001;
   55202: result <= 12'b111010110001;
   55203: result <= 12'b111010110000;
   55204: result <= 12'b111010110000;
   55205: result <= 12'b111010110000;
   55206: result <= 12'b111010110000;
   55207: result <= 12'b111010110000;
   55208: result <= 12'b111010110000;
   55209: result <= 12'b111010110000;
   55210: result <= 12'b111010110000;
   55211: result <= 12'b111010110000;
   55212: result <= 12'b111010101111;
   55213: result <= 12'b111010101111;
   55214: result <= 12'b111010101111;
   55215: result <= 12'b111010101111;
   55216: result <= 12'b111010101111;
   55217: result <= 12'b111010101111;
   55218: result <= 12'b111010101111;
   55219: result <= 12'b111010101111;
   55220: result <= 12'b111010101111;
   55221: result <= 12'b111010101110;
   55222: result <= 12'b111010101110;
   55223: result <= 12'b111010101110;
   55224: result <= 12'b111010101110;
   55225: result <= 12'b111010101110;
   55226: result <= 12'b111010101110;
   55227: result <= 12'b111010101110;
   55228: result <= 12'b111010101110;
   55229: result <= 12'b111010101110;
   55230: result <= 12'b111010101110;
   55231: result <= 12'b111010101101;
   55232: result <= 12'b111010101101;
   55233: result <= 12'b111010101101;
   55234: result <= 12'b111010101101;
   55235: result <= 12'b111010101101;
   55236: result <= 12'b111010101101;
   55237: result <= 12'b111010101101;
   55238: result <= 12'b111010101101;
   55239: result <= 12'b111010101101;
   55240: result <= 12'b111010101100;
   55241: result <= 12'b111010101100;
   55242: result <= 12'b111010101100;
   55243: result <= 12'b111010101100;
   55244: result <= 12'b111010101100;
   55245: result <= 12'b111010101100;
   55246: result <= 12'b111010101100;
   55247: result <= 12'b111010101100;
   55248: result <= 12'b111010101100;
   55249: result <= 12'b111010101011;
   55250: result <= 12'b111010101011;
   55251: result <= 12'b111010101011;
   55252: result <= 12'b111010101011;
   55253: result <= 12'b111010101011;
   55254: result <= 12'b111010101011;
   55255: result <= 12'b111010101011;
   55256: result <= 12'b111010101011;
   55257: result <= 12'b111010101011;
   55258: result <= 12'b111010101010;
   55259: result <= 12'b111010101010;
   55260: result <= 12'b111010101010;
   55261: result <= 12'b111010101010;
   55262: result <= 12'b111010101010;
   55263: result <= 12'b111010101010;
   55264: result <= 12'b111010101010;
   55265: result <= 12'b111010101010;
   55266: result <= 12'b111010101010;
   55267: result <= 12'b111010101010;
   55268: result <= 12'b111010101001;
   55269: result <= 12'b111010101001;
   55270: result <= 12'b111010101001;
   55271: result <= 12'b111010101001;
   55272: result <= 12'b111010101001;
   55273: result <= 12'b111010101001;
   55274: result <= 12'b111010101001;
   55275: result <= 12'b111010101001;
   55276: result <= 12'b111010101001;
   55277: result <= 12'b111010101000;
   55278: result <= 12'b111010101000;
   55279: result <= 12'b111010101000;
   55280: result <= 12'b111010101000;
   55281: result <= 12'b111010101000;
   55282: result <= 12'b111010101000;
   55283: result <= 12'b111010101000;
   55284: result <= 12'b111010101000;
   55285: result <= 12'b111010101000;
   55286: result <= 12'b111010100111;
   55287: result <= 12'b111010100111;
   55288: result <= 12'b111010100111;
   55289: result <= 12'b111010100111;
   55290: result <= 12'b111010100111;
   55291: result <= 12'b111010100111;
   55292: result <= 12'b111010100111;
   55293: result <= 12'b111010100111;
   55294: result <= 12'b111010100111;
   55295: result <= 12'b111010100110;
   55296: result <= 12'b111010100110;
   55297: result <= 12'b111010100110;
   55298: result <= 12'b111010100110;
   55299: result <= 12'b111010100110;
   55300: result <= 12'b111010100110;
   55301: result <= 12'b111010100110;
   55302: result <= 12'b111010100110;
   55303: result <= 12'b111010100110;
   55304: result <= 12'b111010100101;
   55305: result <= 12'b111010100101;
   55306: result <= 12'b111010100101;
   55307: result <= 12'b111010100101;
   55308: result <= 12'b111010100101;
   55309: result <= 12'b111010100101;
   55310: result <= 12'b111010100101;
   55311: result <= 12'b111010100101;
   55312: result <= 12'b111010100101;
   55313: result <= 12'b111010100100;
   55314: result <= 12'b111010100100;
   55315: result <= 12'b111010100100;
   55316: result <= 12'b111010100100;
   55317: result <= 12'b111010100100;
   55318: result <= 12'b111010100100;
   55319: result <= 12'b111010100100;
   55320: result <= 12'b111010100100;
   55321: result <= 12'b111010100100;
   55322: result <= 12'b111010100100;
   55323: result <= 12'b111010100011;
   55324: result <= 12'b111010100011;
   55325: result <= 12'b111010100011;
   55326: result <= 12'b111010100011;
   55327: result <= 12'b111010100011;
   55328: result <= 12'b111010100011;
   55329: result <= 12'b111010100011;
   55330: result <= 12'b111010100011;
   55331: result <= 12'b111010100011;
   55332: result <= 12'b111010100010;
   55333: result <= 12'b111010100010;
   55334: result <= 12'b111010100010;
   55335: result <= 12'b111010100010;
   55336: result <= 12'b111010100010;
   55337: result <= 12'b111010100010;
   55338: result <= 12'b111010100010;
   55339: result <= 12'b111010100010;
   55340: result <= 12'b111010100010;
   55341: result <= 12'b111010100001;
   55342: result <= 12'b111010100001;
   55343: result <= 12'b111010100001;
   55344: result <= 12'b111010100001;
   55345: result <= 12'b111010100001;
   55346: result <= 12'b111010100001;
   55347: result <= 12'b111010100001;
   55348: result <= 12'b111010100001;
   55349: result <= 12'b111010100001;
   55350: result <= 12'b111010100000;
   55351: result <= 12'b111010100000;
   55352: result <= 12'b111010100000;
   55353: result <= 12'b111010100000;
   55354: result <= 12'b111010100000;
   55355: result <= 12'b111010100000;
   55356: result <= 12'b111010100000;
   55357: result <= 12'b111010100000;
   55358: result <= 12'b111010100000;
   55359: result <= 12'b111010011111;
   55360: result <= 12'b111010011111;
   55361: result <= 12'b111010011111;
   55362: result <= 12'b111010011111;
   55363: result <= 12'b111010011111;
   55364: result <= 12'b111010011111;
   55365: result <= 12'b111010011111;
   55366: result <= 12'b111010011111;
   55367: result <= 12'b111010011111;
   55368: result <= 12'b111010011110;
   55369: result <= 12'b111010011110;
   55370: result <= 12'b111010011110;
   55371: result <= 12'b111010011110;
   55372: result <= 12'b111010011110;
   55373: result <= 12'b111010011110;
   55374: result <= 12'b111010011110;
   55375: result <= 12'b111010011110;
   55376: result <= 12'b111010011110;
   55377: result <= 12'b111010011101;
   55378: result <= 12'b111010011101;
   55379: result <= 12'b111010011101;
   55380: result <= 12'b111010011101;
   55381: result <= 12'b111010011101;
   55382: result <= 12'b111010011101;
   55383: result <= 12'b111010011101;
   55384: result <= 12'b111010011101;
   55385: result <= 12'b111010011101;
   55386: result <= 12'b111010011100;
   55387: result <= 12'b111010011100;
   55388: result <= 12'b111010011100;
   55389: result <= 12'b111010011100;
   55390: result <= 12'b111010011100;
   55391: result <= 12'b111010011100;
   55392: result <= 12'b111010011100;
   55393: result <= 12'b111010011100;
   55394: result <= 12'b111010011100;
   55395: result <= 12'b111010011011;
   55396: result <= 12'b111010011011;
   55397: result <= 12'b111010011011;
   55398: result <= 12'b111010011011;
   55399: result <= 12'b111010011011;
   55400: result <= 12'b111010011011;
   55401: result <= 12'b111010011011;
   55402: result <= 12'b111010011011;
   55403: result <= 12'b111010011011;
   55404: result <= 12'b111010011010;
   55405: result <= 12'b111010011010;
   55406: result <= 12'b111010011010;
   55407: result <= 12'b111010011010;
   55408: result <= 12'b111010011010;
   55409: result <= 12'b111010011010;
   55410: result <= 12'b111010011010;
   55411: result <= 12'b111010011010;
   55412: result <= 12'b111010011010;
   55413: result <= 12'b111010011001;
   55414: result <= 12'b111010011001;
   55415: result <= 12'b111010011001;
   55416: result <= 12'b111010011001;
   55417: result <= 12'b111010011001;
   55418: result <= 12'b111010011001;
   55419: result <= 12'b111010011001;
   55420: result <= 12'b111010011001;
   55421: result <= 12'b111010011001;
   55422: result <= 12'b111010011000;
   55423: result <= 12'b111010011000;
   55424: result <= 12'b111010011000;
   55425: result <= 12'b111010011000;
   55426: result <= 12'b111010011000;
   55427: result <= 12'b111010011000;
   55428: result <= 12'b111010011000;
   55429: result <= 12'b111010011000;
   55430: result <= 12'b111010011000;
   55431: result <= 12'b111010010111;
   55432: result <= 12'b111010010111;
   55433: result <= 12'b111010010111;
   55434: result <= 12'b111010010111;
   55435: result <= 12'b111010010111;
   55436: result <= 12'b111010010111;
   55437: result <= 12'b111010010111;
   55438: result <= 12'b111010010111;
   55439: result <= 12'b111010010111;
   55440: result <= 12'b111010010110;
   55441: result <= 12'b111010010110;
   55442: result <= 12'b111010010110;
   55443: result <= 12'b111010010110;
   55444: result <= 12'b111010010110;
   55445: result <= 12'b111010010110;
   55446: result <= 12'b111010010110;
   55447: result <= 12'b111010010110;
   55448: result <= 12'b111010010110;
   55449: result <= 12'b111010010101;
   55450: result <= 12'b111010010101;
   55451: result <= 12'b111010010101;
   55452: result <= 12'b111010010101;
   55453: result <= 12'b111010010101;
   55454: result <= 12'b111010010101;
   55455: result <= 12'b111010010101;
   55456: result <= 12'b111010010101;
   55457: result <= 12'b111010010101;
   55458: result <= 12'b111010010100;
   55459: result <= 12'b111010010100;
   55460: result <= 12'b111010010100;
   55461: result <= 12'b111010010100;
   55462: result <= 12'b111010010100;
   55463: result <= 12'b111010010100;
   55464: result <= 12'b111010010100;
   55465: result <= 12'b111010010100;
   55466: result <= 12'b111010010100;
   55467: result <= 12'b111010010011;
   55468: result <= 12'b111010010011;
   55469: result <= 12'b111010010011;
   55470: result <= 12'b111010010011;
   55471: result <= 12'b111010010011;
   55472: result <= 12'b111010010011;
   55473: result <= 12'b111010010011;
   55474: result <= 12'b111010010011;
   55475: result <= 12'b111010010011;
   55476: result <= 12'b111010010010;
   55477: result <= 12'b111010010010;
   55478: result <= 12'b111010010010;
   55479: result <= 12'b111010010010;
   55480: result <= 12'b111010010010;
   55481: result <= 12'b111010010010;
   55482: result <= 12'b111010010010;
   55483: result <= 12'b111010010010;
   55484: result <= 12'b111010010010;
   55485: result <= 12'b111010010001;
   55486: result <= 12'b111010010001;
   55487: result <= 12'b111010010001;
   55488: result <= 12'b111010010001;
   55489: result <= 12'b111010010001;
   55490: result <= 12'b111010010001;
   55491: result <= 12'b111010010001;
   55492: result <= 12'b111010010001;
   55493: result <= 12'b111010010001;
   55494: result <= 12'b111010010000;
   55495: result <= 12'b111010010000;
   55496: result <= 12'b111010010000;
   55497: result <= 12'b111010010000;
   55498: result <= 12'b111010010000;
   55499: result <= 12'b111010010000;
   55500: result <= 12'b111010010000;
   55501: result <= 12'b111010010000;
   55502: result <= 12'b111010010000;
   55503: result <= 12'b111010001111;
   55504: result <= 12'b111010001111;
   55505: result <= 12'b111010001111;
   55506: result <= 12'b111010001111;
   55507: result <= 12'b111010001111;
   55508: result <= 12'b111010001111;
   55509: result <= 12'b111010001111;
   55510: result <= 12'b111010001111;
   55511: result <= 12'b111010001111;
   55512: result <= 12'b111010001110;
   55513: result <= 12'b111010001110;
   55514: result <= 12'b111010001110;
   55515: result <= 12'b111010001110;
   55516: result <= 12'b111010001110;
   55517: result <= 12'b111010001110;
   55518: result <= 12'b111010001110;
   55519: result <= 12'b111010001110;
   55520: result <= 12'b111010001110;
   55521: result <= 12'b111010001101;
   55522: result <= 12'b111010001101;
   55523: result <= 12'b111010001101;
   55524: result <= 12'b111010001101;
   55525: result <= 12'b111010001101;
   55526: result <= 12'b111010001101;
   55527: result <= 12'b111010001101;
   55528: result <= 12'b111010001101;
   55529: result <= 12'b111010001101;
   55530: result <= 12'b111010001100;
   55531: result <= 12'b111010001100;
   55532: result <= 12'b111010001100;
   55533: result <= 12'b111010001100;
   55534: result <= 12'b111010001100;
   55535: result <= 12'b111010001100;
   55536: result <= 12'b111010001100;
   55537: result <= 12'b111010001100;
   55538: result <= 12'b111010001011;
   55539: result <= 12'b111010001011;
   55540: result <= 12'b111010001011;
   55541: result <= 12'b111010001011;
   55542: result <= 12'b111010001011;
   55543: result <= 12'b111010001011;
   55544: result <= 12'b111010001011;
   55545: result <= 12'b111010001011;
   55546: result <= 12'b111010001011;
   55547: result <= 12'b111010001010;
   55548: result <= 12'b111010001010;
   55549: result <= 12'b111010001010;
   55550: result <= 12'b111010001010;
   55551: result <= 12'b111010001010;
   55552: result <= 12'b111010001010;
   55553: result <= 12'b111010001010;
   55554: result <= 12'b111010001010;
   55555: result <= 12'b111010001010;
   55556: result <= 12'b111010001001;
   55557: result <= 12'b111010001001;
   55558: result <= 12'b111010001001;
   55559: result <= 12'b111010001001;
   55560: result <= 12'b111010001001;
   55561: result <= 12'b111010001001;
   55562: result <= 12'b111010001001;
   55563: result <= 12'b111010001001;
   55564: result <= 12'b111010001001;
   55565: result <= 12'b111010001000;
   55566: result <= 12'b111010001000;
   55567: result <= 12'b111010001000;
   55568: result <= 12'b111010001000;
   55569: result <= 12'b111010001000;
   55570: result <= 12'b111010001000;
   55571: result <= 12'b111010001000;
   55572: result <= 12'b111010001000;
   55573: result <= 12'b111010001000;
   55574: result <= 12'b111010000111;
   55575: result <= 12'b111010000111;
   55576: result <= 12'b111010000111;
   55577: result <= 12'b111010000111;
   55578: result <= 12'b111010000111;
   55579: result <= 12'b111010000111;
   55580: result <= 12'b111010000111;
   55581: result <= 12'b111010000111;
   55582: result <= 12'b111010000111;
   55583: result <= 12'b111010000110;
   55584: result <= 12'b111010000110;
   55585: result <= 12'b111010000110;
   55586: result <= 12'b111010000110;
   55587: result <= 12'b111010000110;
   55588: result <= 12'b111010000110;
   55589: result <= 12'b111010000110;
   55590: result <= 12'b111010000110;
   55591: result <= 12'b111010000101;
   55592: result <= 12'b111010000101;
   55593: result <= 12'b111010000101;
   55594: result <= 12'b111010000101;
   55595: result <= 12'b111010000101;
   55596: result <= 12'b111010000101;
   55597: result <= 12'b111010000101;
   55598: result <= 12'b111010000101;
   55599: result <= 12'b111010000101;
   55600: result <= 12'b111010000100;
   55601: result <= 12'b111010000100;
   55602: result <= 12'b111010000100;
   55603: result <= 12'b111010000100;
   55604: result <= 12'b111010000100;
   55605: result <= 12'b111010000100;
   55606: result <= 12'b111010000100;
   55607: result <= 12'b111010000100;
   55608: result <= 12'b111010000100;
   55609: result <= 12'b111010000011;
   55610: result <= 12'b111010000011;
   55611: result <= 12'b111010000011;
   55612: result <= 12'b111010000011;
   55613: result <= 12'b111010000011;
   55614: result <= 12'b111010000011;
   55615: result <= 12'b111010000011;
   55616: result <= 12'b111010000011;
   55617: result <= 12'b111010000011;
   55618: result <= 12'b111010000010;
   55619: result <= 12'b111010000010;
   55620: result <= 12'b111010000010;
   55621: result <= 12'b111010000010;
   55622: result <= 12'b111010000010;
   55623: result <= 12'b111010000010;
   55624: result <= 12'b111010000010;
   55625: result <= 12'b111010000010;
   55626: result <= 12'b111010000010;
   55627: result <= 12'b111010000001;
   55628: result <= 12'b111010000001;
   55629: result <= 12'b111010000001;
   55630: result <= 12'b111010000001;
   55631: result <= 12'b111010000001;
   55632: result <= 12'b111010000001;
   55633: result <= 12'b111010000001;
   55634: result <= 12'b111010000001;
   55635: result <= 12'b111010000000;
   55636: result <= 12'b111010000000;
   55637: result <= 12'b111010000000;
   55638: result <= 12'b111010000000;
   55639: result <= 12'b111010000000;
   55640: result <= 12'b111010000000;
   55641: result <= 12'b111010000000;
   55642: result <= 12'b111010000000;
   55643: result <= 12'b111010000000;
   55644: result <= 12'b111001111111;
   55645: result <= 12'b111001111111;
   55646: result <= 12'b111001111111;
   55647: result <= 12'b111001111111;
   55648: result <= 12'b111001111111;
   55649: result <= 12'b111001111111;
   55650: result <= 12'b111001111111;
   55651: result <= 12'b111001111111;
   55652: result <= 12'b111001111111;
   55653: result <= 12'b111001111110;
   55654: result <= 12'b111001111110;
   55655: result <= 12'b111001111110;
   55656: result <= 12'b111001111110;
   55657: result <= 12'b111001111110;
   55658: result <= 12'b111001111110;
   55659: result <= 12'b111001111110;
   55660: result <= 12'b111001111110;
   55661: result <= 12'b111001111101;
   55662: result <= 12'b111001111101;
   55663: result <= 12'b111001111101;
   55664: result <= 12'b111001111101;
   55665: result <= 12'b111001111101;
   55666: result <= 12'b111001111101;
   55667: result <= 12'b111001111101;
   55668: result <= 12'b111001111101;
   55669: result <= 12'b111001111101;
   55670: result <= 12'b111001111100;
   55671: result <= 12'b111001111100;
   55672: result <= 12'b111001111100;
   55673: result <= 12'b111001111100;
   55674: result <= 12'b111001111100;
   55675: result <= 12'b111001111100;
   55676: result <= 12'b111001111100;
   55677: result <= 12'b111001111100;
   55678: result <= 12'b111001111100;
   55679: result <= 12'b111001111011;
   55680: result <= 12'b111001111011;
   55681: result <= 12'b111001111011;
   55682: result <= 12'b111001111011;
   55683: result <= 12'b111001111011;
   55684: result <= 12'b111001111011;
   55685: result <= 12'b111001111011;
   55686: result <= 12'b111001111011;
   55687: result <= 12'b111001111011;
   55688: result <= 12'b111001111010;
   55689: result <= 12'b111001111010;
   55690: result <= 12'b111001111010;
   55691: result <= 12'b111001111010;
   55692: result <= 12'b111001111010;
   55693: result <= 12'b111001111010;
   55694: result <= 12'b111001111010;
   55695: result <= 12'b111001111010;
   55696: result <= 12'b111001111001;
   55697: result <= 12'b111001111001;
   55698: result <= 12'b111001111001;
   55699: result <= 12'b111001111001;
   55700: result <= 12'b111001111001;
   55701: result <= 12'b111001111001;
   55702: result <= 12'b111001111001;
   55703: result <= 12'b111001111001;
   55704: result <= 12'b111001111001;
   55705: result <= 12'b111001111000;
   55706: result <= 12'b111001111000;
   55707: result <= 12'b111001111000;
   55708: result <= 12'b111001111000;
   55709: result <= 12'b111001111000;
   55710: result <= 12'b111001111000;
   55711: result <= 12'b111001111000;
   55712: result <= 12'b111001111000;
   55713: result <= 12'b111001111000;
   55714: result <= 12'b111001110111;
   55715: result <= 12'b111001110111;
   55716: result <= 12'b111001110111;
   55717: result <= 12'b111001110111;
   55718: result <= 12'b111001110111;
   55719: result <= 12'b111001110111;
   55720: result <= 12'b111001110111;
   55721: result <= 12'b111001110111;
   55722: result <= 12'b111001110110;
   55723: result <= 12'b111001110110;
   55724: result <= 12'b111001110110;
   55725: result <= 12'b111001110110;
   55726: result <= 12'b111001110110;
   55727: result <= 12'b111001110110;
   55728: result <= 12'b111001110110;
   55729: result <= 12'b111001110110;
   55730: result <= 12'b111001110110;
   55731: result <= 12'b111001110101;
   55732: result <= 12'b111001110101;
   55733: result <= 12'b111001110101;
   55734: result <= 12'b111001110101;
   55735: result <= 12'b111001110101;
   55736: result <= 12'b111001110101;
   55737: result <= 12'b111001110101;
   55738: result <= 12'b111001110101;
   55739: result <= 12'b111001110101;
   55740: result <= 12'b111001110100;
   55741: result <= 12'b111001110100;
   55742: result <= 12'b111001110100;
   55743: result <= 12'b111001110100;
   55744: result <= 12'b111001110100;
   55745: result <= 12'b111001110100;
   55746: result <= 12'b111001110100;
   55747: result <= 12'b111001110100;
   55748: result <= 12'b111001110011;
   55749: result <= 12'b111001110011;
   55750: result <= 12'b111001110011;
   55751: result <= 12'b111001110011;
   55752: result <= 12'b111001110011;
   55753: result <= 12'b111001110011;
   55754: result <= 12'b111001110011;
   55755: result <= 12'b111001110011;
   55756: result <= 12'b111001110011;
   55757: result <= 12'b111001110010;
   55758: result <= 12'b111001110010;
   55759: result <= 12'b111001110010;
   55760: result <= 12'b111001110010;
   55761: result <= 12'b111001110010;
   55762: result <= 12'b111001110010;
   55763: result <= 12'b111001110010;
   55764: result <= 12'b111001110010;
   55765: result <= 12'b111001110001;
   55766: result <= 12'b111001110001;
   55767: result <= 12'b111001110001;
   55768: result <= 12'b111001110001;
   55769: result <= 12'b111001110001;
   55770: result <= 12'b111001110001;
   55771: result <= 12'b111001110001;
   55772: result <= 12'b111001110001;
   55773: result <= 12'b111001110001;
   55774: result <= 12'b111001110000;
   55775: result <= 12'b111001110000;
   55776: result <= 12'b111001110000;
   55777: result <= 12'b111001110000;
   55778: result <= 12'b111001110000;
   55779: result <= 12'b111001110000;
   55780: result <= 12'b111001110000;
   55781: result <= 12'b111001110000;
   55782: result <= 12'b111001110000;
   55783: result <= 12'b111001101111;
   55784: result <= 12'b111001101111;
   55785: result <= 12'b111001101111;
   55786: result <= 12'b111001101111;
   55787: result <= 12'b111001101111;
   55788: result <= 12'b111001101111;
   55789: result <= 12'b111001101111;
   55790: result <= 12'b111001101111;
   55791: result <= 12'b111001101110;
   55792: result <= 12'b111001101110;
   55793: result <= 12'b111001101110;
   55794: result <= 12'b111001101110;
   55795: result <= 12'b111001101110;
   55796: result <= 12'b111001101110;
   55797: result <= 12'b111001101110;
   55798: result <= 12'b111001101110;
   55799: result <= 12'b111001101110;
   55800: result <= 12'b111001101101;
   55801: result <= 12'b111001101101;
   55802: result <= 12'b111001101101;
   55803: result <= 12'b111001101101;
   55804: result <= 12'b111001101101;
   55805: result <= 12'b111001101101;
   55806: result <= 12'b111001101101;
   55807: result <= 12'b111001101101;
   55808: result <= 12'b111001101100;
   55809: result <= 12'b111001101100;
   55810: result <= 12'b111001101100;
   55811: result <= 12'b111001101100;
   55812: result <= 12'b111001101100;
   55813: result <= 12'b111001101100;
   55814: result <= 12'b111001101100;
   55815: result <= 12'b111001101100;
   55816: result <= 12'b111001101100;
   55817: result <= 12'b111001101011;
   55818: result <= 12'b111001101011;
   55819: result <= 12'b111001101011;
   55820: result <= 12'b111001101011;
   55821: result <= 12'b111001101011;
   55822: result <= 12'b111001101011;
   55823: result <= 12'b111001101011;
   55824: result <= 12'b111001101011;
   55825: result <= 12'b111001101010;
   55826: result <= 12'b111001101010;
   55827: result <= 12'b111001101010;
   55828: result <= 12'b111001101010;
   55829: result <= 12'b111001101010;
   55830: result <= 12'b111001101010;
   55831: result <= 12'b111001101010;
   55832: result <= 12'b111001101010;
   55833: result <= 12'b111001101010;
   55834: result <= 12'b111001101001;
   55835: result <= 12'b111001101001;
   55836: result <= 12'b111001101001;
   55837: result <= 12'b111001101001;
   55838: result <= 12'b111001101001;
   55839: result <= 12'b111001101001;
   55840: result <= 12'b111001101001;
   55841: result <= 12'b111001101001;
   55842: result <= 12'b111001101000;
   55843: result <= 12'b111001101000;
   55844: result <= 12'b111001101000;
   55845: result <= 12'b111001101000;
   55846: result <= 12'b111001101000;
   55847: result <= 12'b111001101000;
   55848: result <= 12'b111001101000;
   55849: result <= 12'b111001101000;
   55850: result <= 12'b111001101000;
   55851: result <= 12'b111001100111;
   55852: result <= 12'b111001100111;
   55853: result <= 12'b111001100111;
   55854: result <= 12'b111001100111;
   55855: result <= 12'b111001100111;
   55856: result <= 12'b111001100111;
   55857: result <= 12'b111001100111;
   55858: result <= 12'b111001100111;
   55859: result <= 12'b111001100110;
   55860: result <= 12'b111001100110;
   55861: result <= 12'b111001100110;
   55862: result <= 12'b111001100110;
   55863: result <= 12'b111001100110;
   55864: result <= 12'b111001100110;
   55865: result <= 12'b111001100110;
   55866: result <= 12'b111001100110;
   55867: result <= 12'b111001100110;
   55868: result <= 12'b111001100101;
   55869: result <= 12'b111001100101;
   55870: result <= 12'b111001100101;
   55871: result <= 12'b111001100101;
   55872: result <= 12'b111001100101;
   55873: result <= 12'b111001100101;
   55874: result <= 12'b111001100101;
   55875: result <= 12'b111001100101;
   55876: result <= 12'b111001100100;
   55877: result <= 12'b111001100100;
   55878: result <= 12'b111001100100;
   55879: result <= 12'b111001100100;
   55880: result <= 12'b111001100100;
   55881: result <= 12'b111001100100;
   55882: result <= 12'b111001100100;
   55883: result <= 12'b111001100100;
   55884: result <= 12'b111001100100;
   55885: result <= 12'b111001100011;
   55886: result <= 12'b111001100011;
   55887: result <= 12'b111001100011;
   55888: result <= 12'b111001100011;
   55889: result <= 12'b111001100011;
   55890: result <= 12'b111001100011;
   55891: result <= 12'b111001100011;
   55892: result <= 12'b111001100011;
   55893: result <= 12'b111001100010;
   55894: result <= 12'b111001100010;
   55895: result <= 12'b111001100010;
   55896: result <= 12'b111001100010;
   55897: result <= 12'b111001100010;
   55898: result <= 12'b111001100010;
   55899: result <= 12'b111001100010;
   55900: result <= 12'b111001100010;
   55901: result <= 12'b111001100010;
   55902: result <= 12'b111001100001;
   55903: result <= 12'b111001100001;
   55904: result <= 12'b111001100001;
   55905: result <= 12'b111001100001;
   55906: result <= 12'b111001100001;
   55907: result <= 12'b111001100001;
   55908: result <= 12'b111001100001;
   55909: result <= 12'b111001100001;
   55910: result <= 12'b111001100000;
   55911: result <= 12'b111001100000;
   55912: result <= 12'b111001100000;
   55913: result <= 12'b111001100000;
   55914: result <= 12'b111001100000;
   55915: result <= 12'b111001100000;
   55916: result <= 12'b111001100000;
   55917: result <= 12'b111001100000;
   55918: result <= 12'b111001100000;
   55919: result <= 12'b111001011111;
   55920: result <= 12'b111001011111;
   55921: result <= 12'b111001011111;
   55922: result <= 12'b111001011111;
   55923: result <= 12'b111001011111;
   55924: result <= 12'b111001011111;
   55925: result <= 12'b111001011111;
   55926: result <= 12'b111001011111;
   55927: result <= 12'b111001011110;
   55928: result <= 12'b111001011110;
   55929: result <= 12'b111001011110;
   55930: result <= 12'b111001011110;
   55931: result <= 12'b111001011110;
   55932: result <= 12'b111001011110;
   55933: result <= 12'b111001011110;
   55934: result <= 12'b111001011110;
   55935: result <= 12'b111001011101;
   55936: result <= 12'b111001011101;
   55937: result <= 12'b111001011101;
   55938: result <= 12'b111001011101;
   55939: result <= 12'b111001011101;
   55940: result <= 12'b111001011101;
   55941: result <= 12'b111001011101;
   55942: result <= 12'b111001011101;
   55943: result <= 12'b111001011101;
   55944: result <= 12'b111001011100;
   55945: result <= 12'b111001011100;
   55946: result <= 12'b111001011100;
   55947: result <= 12'b111001011100;
   55948: result <= 12'b111001011100;
   55949: result <= 12'b111001011100;
   55950: result <= 12'b111001011100;
   55951: result <= 12'b111001011100;
   55952: result <= 12'b111001011011;
   55953: result <= 12'b111001011011;
   55954: result <= 12'b111001011011;
   55955: result <= 12'b111001011011;
   55956: result <= 12'b111001011011;
   55957: result <= 12'b111001011011;
   55958: result <= 12'b111001011011;
   55959: result <= 12'b111001011011;
   55960: result <= 12'b111001011011;
   55961: result <= 12'b111001011010;
   55962: result <= 12'b111001011010;
   55963: result <= 12'b111001011010;
   55964: result <= 12'b111001011010;
   55965: result <= 12'b111001011010;
   55966: result <= 12'b111001011010;
   55967: result <= 12'b111001011010;
   55968: result <= 12'b111001011010;
   55969: result <= 12'b111001011001;
   55970: result <= 12'b111001011001;
   55971: result <= 12'b111001011001;
   55972: result <= 12'b111001011001;
   55973: result <= 12'b111001011001;
   55974: result <= 12'b111001011001;
   55975: result <= 12'b111001011001;
   55976: result <= 12'b111001011001;
   55977: result <= 12'b111001011000;
   55978: result <= 12'b111001011000;
   55979: result <= 12'b111001011000;
   55980: result <= 12'b111001011000;
   55981: result <= 12'b111001011000;
   55982: result <= 12'b111001011000;
   55983: result <= 12'b111001011000;
   55984: result <= 12'b111001011000;
   55985: result <= 12'b111001011000;
   55986: result <= 12'b111001010111;
   55987: result <= 12'b111001010111;
   55988: result <= 12'b111001010111;
   55989: result <= 12'b111001010111;
   55990: result <= 12'b111001010111;
   55991: result <= 12'b111001010111;
   55992: result <= 12'b111001010111;
   55993: result <= 12'b111001010111;
   55994: result <= 12'b111001010110;
   55995: result <= 12'b111001010110;
   55996: result <= 12'b111001010110;
   55997: result <= 12'b111001010110;
   55998: result <= 12'b111001010110;
   55999: result <= 12'b111001010110;
   56000: result <= 12'b111001010110;
   56001: result <= 12'b111001010110;
   56002: result <= 12'b111001010101;
   56003: result <= 12'b111001010101;
   56004: result <= 12'b111001010101;
   56005: result <= 12'b111001010101;
   56006: result <= 12'b111001010101;
   56007: result <= 12'b111001010101;
   56008: result <= 12'b111001010101;
   56009: result <= 12'b111001010101;
   56010: result <= 12'b111001010101;
   56011: result <= 12'b111001010100;
   56012: result <= 12'b111001010100;
   56013: result <= 12'b111001010100;
   56014: result <= 12'b111001010100;
   56015: result <= 12'b111001010100;
   56016: result <= 12'b111001010100;
   56017: result <= 12'b111001010100;
   56018: result <= 12'b111001010100;
   56019: result <= 12'b111001010011;
   56020: result <= 12'b111001010011;
   56021: result <= 12'b111001010011;
   56022: result <= 12'b111001010011;
   56023: result <= 12'b111001010011;
   56024: result <= 12'b111001010011;
   56025: result <= 12'b111001010011;
   56026: result <= 12'b111001010011;
   56027: result <= 12'b111001010010;
   56028: result <= 12'b111001010010;
   56029: result <= 12'b111001010010;
   56030: result <= 12'b111001010010;
   56031: result <= 12'b111001010010;
   56032: result <= 12'b111001010010;
   56033: result <= 12'b111001010010;
   56034: result <= 12'b111001010010;
   56035: result <= 12'b111001010010;
   56036: result <= 12'b111001010001;
   56037: result <= 12'b111001010001;
   56038: result <= 12'b111001010001;
   56039: result <= 12'b111001010001;
   56040: result <= 12'b111001010001;
   56041: result <= 12'b111001010001;
   56042: result <= 12'b111001010001;
   56043: result <= 12'b111001010001;
   56044: result <= 12'b111001010000;
   56045: result <= 12'b111001010000;
   56046: result <= 12'b111001010000;
   56047: result <= 12'b111001010000;
   56048: result <= 12'b111001010000;
   56049: result <= 12'b111001010000;
   56050: result <= 12'b111001010000;
   56051: result <= 12'b111001010000;
   56052: result <= 12'b111001001111;
   56053: result <= 12'b111001001111;
   56054: result <= 12'b111001001111;
   56055: result <= 12'b111001001111;
   56056: result <= 12'b111001001111;
   56057: result <= 12'b111001001111;
   56058: result <= 12'b111001001111;
   56059: result <= 12'b111001001111;
   56060: result <= 12'b111001001111;
   56061: result <= 12'b111001001110;
   56062: result <= 12'b111001001110;
   56063: result <= 12'b111001001110;
   56064: result <= 12'b111001001110;
   56065: result <= 12'b111001001110;
   56066: result <= 12'b111001001110;
   56067: result <= 12'b111001001110;
   56068: result <= 12'b111001001110;
   56069: result <= 12'b111001001101;
   56070: result <= 12'b111001001101;
   56071: result <= 12'b111001001101;
   56072: result <= 12'b111001001101;
   56073: result <= 12'b111001001101;
   56074: result <= 12'b111001001101;
   56075: result <= 12'b111001001101;
   56076: result <= 12'b111001001101;
   56077: result <= 12'b111001001100;
   56078: result <= 12'b111001001100;
   56079: result <= 12'b111001001100;
   56080: result <= 12'b111001001100;
   56081: result <= 12'b111001001100;
   56082: result <= 12'b111001001100;
   56083: result <= 12'b111001001100;
   56084: result <= 12'b111001001100;
   56085: result <= 12'b111001001011;
   56086: result <= 12'b111001001011;
   56087: result <= 12'b111001001011;
   56088: result <= 12'b111001001011;
   56089: result <= 12'b111001001011;
   56090: result <= 12'b111001001011;
   56091: result <= 12'b111001001011;
   56092: result <= 12'b111001001011;
   56093: result <= 12'b111001001011;
   56094: result <= 12'b111001001010;
   56095: result <= 12'b111001001010;
   56096: result <= 12'b111001001010;
   56097: result <= 12'b111001001010;
   56098: result <= 12'b111001001010;
   56099: result <= 12'b111001001010;
   56100: result <= 12'b111001001010;
   56101: result <= 12'b111001001010;
   56102: result <= 12'b111001001001;
   56103: result <= 12'b111001001001;
   56104: result <= 12'b111001001001;
   56105: result <= 12'b111001001001;
   56106: result <= 12'b111001001001;
   56107: result <= 12'b111001001001;
   56108: result <= 12'b111001001001;
   56109: result <= 12'b111001001001;
   56110: result <= 12'b111001001000;
   56111: result <= 12'b111001001000;
   56112: result <= 12'b111001001000;
   56113: result <= 12'b111001001000;
   56114: result <= 12'b111001001000;
   56115: result <= 12'b111001001000;
   56116: result <= 12'b111001001000;
   56117: result <= 12'b111001001000;
   56118: result <= 12'b111001000111;
   56119: result <= 12'b111001000111;
   56120: result <= 12'b111001000111;
   56121: result <= 12'b111001000111;
   56122: result <= 12'b111001000111;
   56123: result <= 12'b111001000111;
   56124: result <= 12'b111001000111;
   56125: result <= 12'b111001000111;
   56126: result <= 12'b111001000111;
   56127: result <= 12'b111001000110;
   56128: result <= 12'b111001000110;
   56129: result <= 12'b111001000110;
   56130: result <= 12'b111001000110;
   56131: result <= 12'b111001000110;
   56132: result <= 12'b111001000110;
   56133: result <= 12'b111001000110;
   56134: result <= 12'b111001000110;
   56135: result <= 12'b111001000101;
   56136: result <= 12'b111001000101;
   56137: result <= 12'b111001000101;
   56138: result <= 12'b111001000101;
   56139: result <= 12'b111001000101;
   56140: result <= 12'b111001000101;
   56141: result <= 12'b111001000101;
   56142: result <= 12'b111001000101;
   56143: result <= 12'b111001000100;
   56144: result <= 12'b111001000100;
   56145: result <= 12'b111001000100;
   56146: result <= 12'b111001000100;
   56147: result <= 12'b111001000100;
   56148: result <= 12'b111001000100;
   56149: result <= 12'b111001000100;
   56150: result <= 12'b111001000100;
   56151: result <= 12'b111001000011;
   56152: result <= 12'b111001000011;
   56153: result <= 12'b111001000011;
   56154: result <= 12'b111001000011;
   56155: result <= 12'b111001000011;
   56156: result <= 12'b111001000011;
   56157: result <= 12'b111001000011;
   56158: result <= 12'b111001000011;
   56159: result <= 12'b111001000010;
   56160: result <= 12'b111001000010;
   56161: result <= 12'b111001000010;
   56162: result <= 12'b111001000010;
   56163: result <= 12'b111001000010;
   56164: result <= 12'b111001000010;
   56165: result <= 12'b111001000010;
   56166: result <= 12'b111001000010;
   56167: result <= 12'b111001000010;
   56168: result <= 12'b111001000001;
   56169: result <= 12'b111001000001;
   56170: result <= 12'b111001000001;
   56171: result <= 12'b111001000001;
   56172: result <= 12'b111001000001;
   56173: result <= 12'b111001000001;
   56174: result <= 12'b111001000001;
   56175: result <= 12'b111001000001;
   56176: result <= 12'b111001000000;
   56177: result <= 12'b111001000000;
   56178: result <= 12'b111001000000;
   56179: result <= 12'b111001000000;
   56180: result <= 12'b111001000000;
   56181: result <= 12'b111001000000;
   56182: result <= 12'b111001000000;
   56183: result <= 12'b111001000000;
   56184: result <= 12'b111000111111;
   56185: result <= 12'b111000111111;
   56186: result <= 12'b111000111111;
   56187: result <= 12'b111000111111;
   56188: result <= 12'b111000111111;
   56189: result <= 12'b111000111111;
   56190: result <= 12'b111000111111;
   56191: result <= 12'b111000111111;
   56192: result <= 12'b111000111110;
   56193: result <= 12'b111000111110;
   56194: result <= 12'b111000111110;
   56195: result <= 12'b111000111110;
   56196: result <= 12'b111000111110;
   56197: result <= 12'b111000111110;
   56198: result <= 12'b111000111110;
   56199: result <= 12'b111000111110;
   56200: result <= 12'b111000111101;
   56201: result <= 12'b111000111101;
   56202: result <= 12'b111000111101;
   56203: result <= 12'b111000111101;
   56204: result <= 12'b111000111101;
   56205: result <= 12'b111000111101;
   56206: result <= 12'b111000111101;
   56207: result <= 12'b111000111101;
   56208: result <= 12'b111000111100;
   56209: result <= 12'b111000111100;
   56210: result <= 12'b111000111100;
   56211: result <= 12'b111000111100;
   56212: result <= 12'b111000111100;
   56213: result <= 12'b111000111100;
   56214: result <= 12'b111000111100;
   56215: result <= 12'b111000111100;
   56216: result <= 12'b111000111100;
   56217: result <= 12'b111000111011;
   56218: result <= 12'b111000111011;
   56219: result <= 12'b111000111011;
   56220: result <= 12'b111000111011;
   56221: result <= 12'b111000111011;
   56222: result <= 12'b111000111011;
   56223: result <= 12'b111000111011;
   56224: result <= 12'b111000111011;
   56225: result <= 12'b111000111010;
   56226: result <= 12'b111000111010;
   56227: result <= 12'b111000111010;
   56228: result <= 12'b111000111010;
   56229: result <= 12'b111000111010;
   56230: result <= 12'b111000111010;
   56231: result <= 12'b111000111010;
   56232: result <= 12'b111000111010;
   56233: result <= 12'b111000111001;
   56234: result <= 12'b111000111001;
   56235: result <= 12'b111000111001;
   56236: result <= 12'b111000111001;
   56237: result <= 12'b111000111001;
   56238: result <= 12'b111000111001;
   56239: result <= 12'b111000111001;
   56240: result <= 12'b111000111001;
   56241: result <= 12'b111000111000;
   56242: result <= 12'b111000111000;
   56243: result <= 12'b111000111000;
   56244: result <= 12'b111000111000;
   56245: result <= 12'b111000111000;
   56246: result <= 12'b111000111000;
   56247: result <= 12'b111000111000;
   56248: result <= 12'b111000111000;
   56249: result <= 12'b111000110111;
   56250: result <= 12'b111000110111;
   56251: result <= 12'b111000110111;
   56252: result <= 12'b111000110111;
   56253: result <= 12'b111000110111;
   56254: result <= 12'b111000110111;
   56255: result <= 12'b111000110111;
   56256: result <= 12'b111000110111;
   56257: result <= 12'b111000110110;
   56258: result <= 12'b111000110110;
   56259: result <= 12'b111000110110;
   56260: result <= 12'b111000110110;
   56261: result <= 12'b111000110110;
   56262: result <= 12'b111000110110;
   56263: result <= 12'b111000110110;
   56264: result <= 12'b111000110110;
   56265: result <= 12'b111000110101;
   56266: result <= 12'b111000110101;
   56267: result <= 12'b111000110101;
   56268: result <= 12'b111000110101;
   56269: result <= 12'b111000110101;
   56270: result <= 12'b111000110101;
   56271: result <= 12'b111000110101;
   56272: result <= 12'b111000110101;
   56273: result <= 12'b111000110100;
   56274: result <= 12'b111000110100;
   56275: result <= 12'b111000110100;
   56276: result <= 12'b111000110100;
   56277: result <= 12'b111000110100;
   56278: result <= 12'b111000110100;
   56279: result <= 12'b111000110100;
   56280: result <= 12'b111000110100;
   56281: result <= 12'b111000110011;
   56282: result <= 12'b111000110011;
   56283: result <= 12'b111000110011;
   56284: result <= 12'b111000110011;
   56285: result <= 12'b111000110011;
   56286: result <= 12'b111000110011;
   56287: result <= 12'b111000110011;
   56288: result <= 12'b111000110011;
   56289: result <= 12'b111000110010;
   56290: result <= 12'b111000110010;
   56291: result <= 12'b111000110010;
   56292: result <= 12'b111000110010;
   56293: result <= 12'b111000110010;
   56294: result <= 12'b111000110010;
   56295: result <= 12'b111000110010;
   56296: result <= 12'b111000110010;
   56297: result <= 12'b111000110001;
   56298: result <= 12'b111000110001;
   56299: result <= 12'b111000110001;
   56300: result <= 12'b111000110001;
   56301: result <= 12'b111000110001;
   56302: result <= 12'b111000110001;
   56303: result <= 12'b111000110001;
   56304: result <= 12'b111000110001;
   56305: result <= 12'b111000110000;
   56306: result <= 12'b111000110000;
   56307: result <= 12'b111000110000;
   56308: result <= 12'b111000110000;
   56309: result <= 12'b111000110000;
   56310: result <= 12'b111000110000;
   56311: result <= 12'b111000110000;
   56312: result <= 12'b111000110000;
   56313: result <= 12'b111000101111;
   56314: result <= 12'b111000101111;
   56315: result <= 12'b111000101111;
   56316: result <= 12'b111000101111;
   56317: result <= 12'b111000101111;
   56318: result <= 12'b111000101111;
   56319: result <= 12'b111000101111;
   56320: result <= 12'b111000101111;
   56321: result <= 12'b111000101111;
   56322: result <= 12'b111000101110;
   56323: result <= 12'b111000101110;
   56324: result <= 12'b111000101110;
   56325: result <= 12'b111000101110;
   56326: result <= 12'b111000101110;
   56327: result <= 12'b111000101110;
   56328: result <= 12'b111000101110;
   56329: result <= 12'b111000101110;
   56330: result <= 12'b111000101101;
   56331: result <= 12'b111000101101;
   56332: result <= 12'b111000101101;
   56333: result <= 12'b111000101101;
   56334: result <= 12'b111000101101;
   56335: result <= 12'b111000101101;
   56336: result <= 12'b111000101101;
   56337: result <= 12'b111000101101;
   56338: result <= 12'b111000101100;
   56339: result <= 12'b111000101100;
   56340: result <= 12'b111000101100;
   56341: result <= 12'b111000101100;
   56342: result <= 12'b111000101100;
   56343: result <= 12'b111000101100;
   56344: result <= 12'b111000101100;
   56345: result <= 12'b111000101100;
   56346: result <= 12'b111000101011;
   56347: result <= 12'b111000101011;
   56348: result <= 12'b111000101011;
   56349: result <= 12'b111000101011;
   56350: result <= 12'b111000101011;
   56351: result <= 12'b111000101011;
   56352: result <= 12'b111000101011;
   56353: result <= 12'b111000101011;
   56354: result <= 12'b111000101010;
   56355: result <= 12'b111000101010;
   56356: result <= 12'b111000101010;
   56357: result <= 12'b111000101010;
   56358: result <= 12'b111000101010;
   56359: result <= 12'b111000101010;
   56360: result <= 12'b111000101010;
   56361: result <= 12'b111000101010;
   56362: result <= 12'b111000101001;
   56363: result <= 12'b111000101001;
   56364: result <= 12'b111000101001;
   56365: result <= 12'b111000101001;
   56366: result <= 12'b111000101001;
   56367: result <= 12'b111000101001;
   56368: result <= 12'b111000101001;
   56369: result <= 12'b111000101001;
   56370: result <= 12'b111000101000;
   56371: result <= 12'b111000101000;
   56372: result <= 12'b111000101000;
   56373: result <= 12'b111000101000;
   56374: result <= 12'b111000101000;
   56375: result <= 12'b111000101000;
   56376: result <= 12'b111000101000;
   56377: result <= 12'b111000101000;
   56378: result <= 12'b111000100111;
   56379: result <= 12'b111000100111;
   56380: result <= 12'b111000100111;
   56381: result <= 12'b111000100111;
   56382: result <= 12'b111000100111;
   56383: result <= 12'b111000100111;
   56384: result <= 12'b111000100111;
   56385: result <= 12'b111000100110;
   56386: result <= 12'b111000100110;
   56387: result <= 12'b111000100110;
   56388: result <= 12'b111000100110;
   56389: result <= 12'b111000100110;
   56390: result <= 12'b111000100110;
   56391: result <= 12'b111000100110;
   56392: result <= 12'b111000100110;
   56393: result <= 12'b111000100101;
   56394: result <= 12'b111000100101;
   56395: result <= 12'b111000100101;
   56396: result <= 12'b111000100101;
   56397: result <= 12'b111000100101;
   56398: result <= 12'b111000100101;
   56399: result <= 12'b111000100101;
   56400: result <= 12'b111000100101;
   56401: result <= 12'b111000100100;
   56402: result <= 12'b111000100100;
   56403: result <= 12'b111000100100;
   56404: result <= 12'b111000100100;
   56405: result <= 12'b111000100100;
   56406: result <= 12'b111000100100;
   56407: result <= 12'b111000100100;
   56408: result <= 12'b111000100100;
   56409: result <= 12'b111000100011;
   56410: result <= 12'b111000100011;
   56411: result <= 12'b111000100011;
   56412: result <= 12'b111000100011;
   56413: result <= 12'b111000100011;
   56414: result <= 12'b111000100011;
   56415: result <= 12'b111000100011;
   56416: result <= 12'b111000100011;
   56417: result <= 12'b111000100010;
   56418: result <= 12'b111000100010;
   56419: result <= 12'b111000100010;
   56420: result <= 12'b111000100010;
   56421: result <= 12'b111000100010;
   56422: result <= 12'b111000100010;
   56423: result <= 12'b111000100010;
   56424: result <= 12'b111000100010;
   56425: result <= 12'b111000100001;
   56426: result <= 12'b111000100001;
   56427: result <= 12'b111000100001;
   56428: result <= 12'b111000100001;
   56429: result <= 12'b111000100001;
   56430: result <= 12'b111000100001;
   56431: result <= 12'b111000100001;
   56432: result <= 12'b111000100001;
   56433: result <= 12'b111000100000;
   56434: result <= 12'b111000100000;
   56435: result <= 12'b111000100000;
   56436: result <= 12'b111000100000;
   56437: result <= 12'b111000100000;
   56438: result <= 12'b111000100000;
   56439: result <= 12'b111000100000;
   56440: result <= 12'b111000100000;
   56441: result <= 12'b111000011111;
   56442: result <= 12'b111000011111;
   56443: result <= 12'b111000011111;
   56444: result <= 12'b111000011111;
   56445: result <= 12'b111000011111;
   56446: result <= 12'b111000011111;
   56447: result <= 12'b111000011111;
   56448: result <= 12'b111000011111;
   56449: result <= 12'b111000011110;
   56450: result <= 12'b111000011110;
   56451: result <= 12'b111000011110;
   56452: result <= 12'b111000011110;
   56453: result <= 12'b111000011110;
   56454: result <= 12'b111000011110;
   56455: result <= 12'b111000011110;
   56456: result <= 12'b111000011110;
   56457: result <= 12'b111000011101;
   56458: result <= 12'b111000011101;
   56459: result <= 12'b111000011101;
   56460: result <= 12'b111000011101;
   56461: result <= 12'b111000011101;
   56462: result <= 12'b111000011101;
   56463: result <= 12'b111000011101;
   56464: result <= 12'b111000011101;
   56465: result <= 12'b111000011100;
   56466: result <= 12'b111000011100;
   56467: result <= 12'b111000011100;
   56468: result <= 12'b111000011100;
   56469: result <= 12'b111000011100;
   56470: result <= 12'b111000011100;
   56471: result <= 12'b111000011100;
   56472: result <= 12'b111000011100;
   56473: result <= 12'b111000011011;
   56474: result <= 12'b111000011011;
   56475: result <= 12'b111000011011;
   56476: result <= 12'b111000011011;
   56477: result <= 12'b111000011011;
   56478: result <= 12'b111000011011;
   56479: result <= 12'b111000011011;
   56480: result <= 12'b111000011011;
   56481: result <= 12'b111000011010;
   56482: result <= 12'b111000011010;
   56483: result <= 12'b111000011010;
   56484: result <= 12'b111000011010;
   56485: result <= 12'b111000011010;
   56486: result <= 12'b111000011010;
   56487: result <= 12'b111000011010;
   56488: result <= 12'b111000011001;
   56489: result <= 12'b111000011001;
   56490: result <= 12'b111000011001;
   56491: result <= 12'b111000011001;
   56492: result <= 12'b111000011001;
   56493: result <= 12'b111000011001;
   56494: result <= 12'b111000011001;
   56495: result <= 12'b111000011001;
   56496: result <= 12'b111000011000;
   56497: result <= 12'b111000011000;
   56498: result <= 12'b111000011000;
   56499: result <= 12'b111000011000;
   56500: result <= 12'b111000011000;
   56501: result <= 12'b111000011000;
   56502: result <= 12'b111000011000;
   56503: result <= 12'b111000011000;
   56504: result <= 12'b111000010111;
   56505: result <= 12'b111000010111;
   56506: result <= 12'b111000010111;
   56507: result <= 12'b111000010111;
   56508: result <= 12'b111000010111;
   56509: result <= 12'b111000010111;
   56510: result <= 12'b111000010111;
   56511: result <= 12'b111000010111;
   56512: result <= 12'b111000010110;
   56513: result <= 12'b111000010110;
   56514: result <= 12'b111000010110;
   56515: result <= 12'b111000010110;
   56516: result <= 12'b111000010110;
   56517: result <= 12'b111000010110;
   56518: result <= 12'b111000010110;
   56519: result <= 12'b111000010110;
   56520: result <= 12'b111000010101;
   56521: result <= 12'b111000010101;
   56522: result <= 12'b111000010101;
   56523: result <= 12'b111000010101;
   56524: result <= 12'b111000010101;
   56525: result <= 12'b111000010101;
   56526: result <= 12'b111000010101;
   56527: result <= 12'b111000010101;
   56528: result <= 12'b111000010100;
   56529: result <= 12'b111000010100;
   56530: result <= 12'b111000010100;
   56531: result <= 12'b111000010100;
   56532: result <= 12'b111000010100;
   56533: result <= 12'b111000010100;
   56534: result <= 12'b111000010100;
   56535: result <= 12'b111000010100;
   56536: result <= 12'b111000010011;
   56537: result <= 12'b111000010011;
   56538: result <= 12'b111000010011;
   56539: result <= 12'b111000010011;
   56540: result <= 12'b111000010011;
   56541: result <= 12'b111000010011;
   56542: result <= 12'b111000010011;
   56543: result <= 12'b111000010010;
   56544: result <= 12'b111000010010;
   56545: result <= 12'b111000010010;
   56546: result <= 12'b111000010010;
   56547: result <= 12'b111000010010;
   56548: result <= 12'b111000010010;
   56549: result <= 12'b111000010010;
   56550: result <= 12'b111000010010;
   56551: result <= 12'b111000010001;
   56552: result <= 12'b111000010001;
   56553: result <= 12'b111000010001;
   56554: result <= 12'b111000010001;
   56555: result <= 12'b111000010001;
   56556: result <= 12'b111000010001;
   56557: result <= 12'b111000010001;
   56558: result <= 12'b111000010001;
   56559: result <= 12'b111000010000;
   56560: result <= 12'b111000010000;
   56561: result <= 12'b111000010000;
   56562: result <= 12'b111000010000;
   56563: result <= 12'b111000010000;
   56564: result <= 12'b111000010000;
   56565: result <= 12'b111000010000;
   56566: result <= 12'b111000010000;
   56567: result <= 12'b111000001111;
   56568: result <= 12'b111000001111;
   56569: result <= 12'b111000001111;
   56570: result <= 12'b111000001111;
   56571: result <= 12'b111000001111;
   56572: result <= 12'b111000001111;
   56573: result <= 12'b111000001111;
   56574: result <= 12'b111000001111;
   56575: result <= 12'b111000001110;
   56576: result <= 12'b111000001110;
   56577: result <= 12'b111000001110;
   56578: result <= 12'b111000001110;
   56579: result <= 12'b111000001110;
   56580: result <= 12'b111000001110;
   56581: result <= 12'b111000001110;
   56582: result <= 12'b111000001101;
   56583: result <= 12'b111000001101;
   56584: result <= 12'b111000001101;
   56585: result <= 12'b111000001101;
   56586: result <= 12'b111000001101;
   56587: result <= 12'b111000001101;
   56588: result <= 12'b111000001101;
   56589: result <= 12'b111000001101;
   56590: result <= 12'b111000001100;
   56591: result <= 12'b111000001100;
   56592: result <= 12'b111000001100;
   56593: result <= 12'b111000001100;
   56594: result <= 12'b111000001100;
   56595: result <= 12'b111000001100;
   56596: result <= 12'b111000001100;
   56597: result <= 12'b111000001100;
   56598: result <= 12'b111000001011;
   56599: result <= 12'b111000001011;
   56600: result <= 12'b111000001011;
   56601: result <= 12'b111000001011;
   56602: result <= 12'b111000001011;
   56603: result <= 12'b111000001011;
   56604: result <= 12'b111000001011;
   56605: result <= 12'b111000001011;
   56606: result <= 12'b111000001010;
   56607: result <= 12'b111000001010;
   56608: result <= 12'b111000001010;
   56609: result <= 12'b111000001010;
   56610: result <= 12'b111000001010;
   56611: result <= 12'b111000001010;
   56612: result <= 12'b111000001010;
   56613: result <= 12'b111000001010;
   56614: result <= 12'b111000001001;
   56615: result <= 12'b111000001001;
   56616: result <= 12'b111000001001;
   56617: result <= 12'b111000001001;
   56618: result <= 12'b111000001001;
   56619: result <= 12'b111000001001;
   56620: result <= 12'b111000001001;
   56621: result <= 12'b111000001000;
   56622: result <= 12'b111000001000;
   56623: result <= 12'b111000001000;
   56624: result <= 12'b111000001000;
   56625: result <= 12'b111000001000;
   56626: result <= 12'b111000001000;
   56627: result <= 12'b111000001000;
   56628: result <= 12'b111000001000;
   56629: result <= 12'b111000000111;
   56630: result <= 12'b111000000111;
   56631: result <= 12'b111000000111;
   56632: result <= 12'b111000000111;
   56633: result <= 12'b111000000111;
   56634: result <= 12'b111000000111;
   56635: result <= 12'b111000000111;
   56636: result <= 12'b111000000111;
   56637: result <= 12'b111000000110;
   56638: result <= 12'b111000000110;
   56639: result <= 12'b111000000110;
   56640: result <= 12'b111000000110;
   56641: result <= 12'b111000000110;
   56642: result <= 12'b111000000110;
   56643: result <= 12'b111000000110;
   56644: result <= 12'b111000000110;
   56645: result <= 12'b111000000101;
   56646: result <= 12'b111000000101;
   56647: result <= 12'b111000000101;
   56648: result <= 12'b111000000101;
   56649: result <= 12'b111000000101;
   56650: result <= 12'b111000000101;
   56651: result <= 12'b111000000101;
   56652: result <= 12'b111000000100;
   56653: result <= 12'b111000000100;
   56654: result <= 12'b111000000100;
   56655: result <= 12'b111000000100;
   56656: result <= 12'b111000000100;
   56657: result <= 12'b111000000100;
   56658: result <= 12'b111000000100;
   56659: result <= 12'b111000000100;
   56660: result <= 12'b111000000011;
   56661: result <= 12'b111000000011;
   56662: result <= 12'b111000000011;
   56663: result <= 12'b111000000011;
   56664: result <= 12'b111000000011;
   56665: result <= 12'b111000000011;
   56666: result <= 12'b111000000011;
   56667: result <= 12'b111000000011;
   56668: result <= 12'b111000000010;
   56669: result <= 12'b111000000010;
   56670: result <= 12'b111000000010;
   56671: result <= 12'b111000000010;
   56672: result <= 12'b111000000010;
   56673: result <= 12'b111000000010;
   56674: result <= 12'b111000000010;
   56675: result <= 12'b111000000001;
   56676: result <= 12'b111000000001;
   56677: result <= 12'b111000000001;
   56678: result <= 12'b111000000001;
   56679: result <= 12'b111000000001;
   56680: result <= 12'b111000000001;
   56681: result <= 12'b111000000001;
   56682: result <= 12'b111000000001;
   56683: result <= 12'b111000000000;
   56684: result <= 12'b111000000000;
   56685: result <= 12'b111000000000;
   56686: result <= 12'b111000000000;
   56687: result <= 12'b111000000000;
   56688: result <= 12'b111000000000;
   56689: result <= 12'b111000000000;
   56690: result <= 12'b111000000000;
   56691: result <= 12'b110111111111;
   56692: result <= 12'b110111111111;
   56693: result <= 12'b110111111111;
   56694: result <= 12'b110111111111;
   56695: result <= 12'b110111111111;
   56696: result <= 12'b110111111111;
   56697: result <= 12'b110111111111;
   56698: result <= 12'b110111111111;
   56699: result <= 12'b110111111110;
   56700: result <= 12'b110111111110;
   56701: result <= 12'b110111111110;
   56702: result <= 12'b110111111110;
   56703: result <= 12'b110111111110;
   56704: result <= 12'b110111111110;
   56705: result <= 12'b110111111110;
   56706: result <= 12'b110111111101;
   56707: result <= 12'b110111111101;
   56708: result <= 12'b110111111101;
   56709: result <= 12'b110111111101;
   56710: result <= 12'b110111111101;
   56711: result <= 12'b110111111101;
   56712: result <= 12'b110111111101;
   56713: result <= 12'b110111111101;
   56714: result <= 12'b110111111100;
   56715: result <= 12'b110111111100;
   56716: result <= 12'b110111111100;
   56717: result <= 12'b110111111100;
   56718: result <= 12'b110111111100;
   56719: result <= 12'b110111111100;
   56720: result <= 12'b110111111100;
   56721: result <= 12'b110111111100;
   56722: result <= 12'b110111111011;
   56723: result <= 12'b110111111011;
   56724: result <= 12'b110111111011;
   56725: result <= 12'b110111111011;
   56726: result <= 12'b110111111011;
   56727: result <= 12'b110111111011;
   56728: result <= 12'b110111111011;
   56729: result <= 12'b110111111010;
   56730: result <= 12'b110111111010;
   56731: result <= 12'b110111111010;
   56732: result <= 12'b110111111010;
   56733: result <= 12'b110111111010;
   56734: result <= 12'b110111111010;
   56735: result <= 12'b110111111010;
   56736: result <= 12'b110111111010;
   56737: result <= 12'b110111111001;
   56738: result <= 12'b110111111001;
   56739: result <= 12'b110111111001;
   56740: result <= 12'b110111111001;
   56741: result <= 12'b110111111001;
   56742: result <= 12'b110111111001;
   56743: result <= 12'b110111111001;
   56744: result <= 12'b110111111001;
   56745: result <= 12'b110111111000;
   56746: result <= 12'b110111111000;
   56747: result <= 12'b110111111000;
   56748: result <= 12'b110111111000;
   56749: result <= 12'b110111111000;
   56750: result <= 12'b110111111000;
   56751: result <= 12'b110111111000;
   56752: result <= 12'b110111110111;
   56753: result <= 12'b110111110111;
   56754: result <= 12'b110111110111;
   56755: result <= 12'b110111110111;
   56756: result <= 12'b110111110111;
   56757: result <= 12'b110111110111;
   56758: result <= 12'b110111110111;
   56759: result <= 12'b110111110111;
   56760: result <= 12'b110111110110;
   56761: result <= 12'b110111110110;
   56762: result <= 12'b110111110110;
   56763: result <= 12'b110111110110;
   56764: result <= 12'b110111110110;
   56765: result <= 12'b110111110110;
   56766: result <= 12'b110111110110;
   56767: result <= 12'b110111110110;
   56768: result <= 12'b110111110101;
   56769: result <= 12'b110111110101;
   56770: result <= 12'b110111110101;
   56771: result <= 12'b110111110101;
   56772: result <= 12'b110111110101;
   56773: result <= 12'b110111110101;
   56774: result <= 12'b110111110101;
   56775: result <= 12'b110111110100;
   56776: result <= 12'b110111110100;
   56777: result <= 12'b110111110100;
   56778: result <= 12'b110111110100;
   56779: result <= 12'b110111110100;
   56780: result <= 12'b110111110100;
   56781: result <= 12'b110111110100;
   56782: result <= 12'b110111110100;
   56783: result <= 12'b110111110011;
   56784: result <= 12'b110111110011;
   56785: result <= 12'b110111110011;
   56786: result <= 12'b110111110011;
   56787: result <= 12'b110111110011;
   56788: result <= 12'b110111110011;
   56789: result <= 12'b110111110011;
   56790: result <= 12'b110111110010;
   56791: result <= 12'b110111110010;
   56792: result <= 12'b110111110010;
   56793: result <= 12'b110111110010;
   56794: result <= 12'b110111110010;
   56795: result <= 12'b110111110010;
   56796: result <= 12'b110111110010;
   56797: result <= 12'b110111110010;
   56798: result <= 12'b110111110001;
   56799: result <= 12'b110111110001;
   56800: result <= 12'b110111110001;
   56801: result <= 12'b110111110001;
   56802: result <= 12'b110111110001;
   56803: result <= 12'b110111110001;
   56804: result <= 12'b110111110001;
   56805: result <= 12'b110111110001;
   56806: result <= 12'b110111110000;
   56807: result <= 12'b110111110000;
   56808: result <= 12'b110111110000;
   56809: result <= 12'b110111110000;
   56810: result <= 12'b110111110000;
   56811: result <= 12'b110111110000;
   56812: result <= 12'b110111110000;
   56813: result <= 12'b110111101111;
   56814: result <= 12'b110111101111;
   56815: result <= 12'b110111101111;
   56816: result <= 12'b110111101111;
   56817: result <= 12'b110111101111;
   56818: result <= 12'b110111101111;
   56819: result <= 12'b110111101111;
   56820: result <= 12'b110111101111;
   56821: result <= 12'b110111101110;
   56822: result <= 12'b110111101110;
   56823: result <= 12'b110111101110;
   56824: result <= 12'b110111101110;
   56825: result <= 12'b110111101110;
   56826: result <= 12'b110111101110;
   56827: result <= 12'b110111101110;
   56828: result <= 12'b110111101101;
   56829: result <= 12'b110111101101;
   56830: result <= 12'b110111101101;
   56831: result <= 12'b110111101101;
   56832: result <= 12'b110111101101;
   56833: result <= 12'b110111101101;
   56834: result <= 12'b110111101101;
   56835: result <= 12'b110111101101;
   56836: result <= 12'b110111101100;
   56837: result <= 12'b110111101100;
   56838: result <= 12'b110111101100;
   56839: result <= 12'b110111101100;
   56840: result <= 12'b110111101100;
   56841: result <= 12'b110111101100;
   56842: result <= 12'b110111101100;
   56843: result <= 12'b110111101100;
   56844: result <= 12'b110111101011;
   56845: result <= 12'b110111101011;
   56846: result <= 12'b110111101011;
   56847: result <= 12'b110111101011;
   56848: result <= 12'b110111101011;
   56849: result <= 12'b110111101011;
   56850: result <= 12'b110111101011;
   56851: result <= 12'b110111101010;
   56852: result <= 12'b110111101010;
   56853: result <= 12'b110111101010;
   56854: result <= 12'b110111101010;
   56855: result <= 12'b110111101010;
   56856: result <= 12'b110111101010;
   56857: result <= 12'b110111101010;
   56858: result <= 12'b110111101010;
   56859: result <= 12'b110111101001;
   56860: result <= 12'b110111101001;
   56861: result <= 12'b110111101001;
   56862: result <= 12'b110111101001;
   56863: result <= 12'b110111101001;
   56864: result <= 12'b110111101001;
   56865: result <= 12'b110111101001;
   56866: result <= 12'b110111101000;
   56867: result <= 12'b110111101000;
   56868: result <= 12'b110111101000;
   56869: result <= 12'b110111101000;
   56870: result <= 12'b110111101000;
   56871: result <= 12'b110111101000;
   56872: result <= 12'b110111101000;
   56873: result <= 12'b110111101000;
   56874: result <= 12'b110111100111;
   56875: result <= 12'b110111100111;
   56876: result <= 12'b110111100111;
   56877: result <= 12'b110111100111;
   56878: result <= 12'b110111100111;
   56879: result <= 12'b110111100111;
   56880: result <= 12'b110111100111;
   56881: result <= 12'b110111100110;
   56882: result <= 12'b110111100110;
   56883: result <= 12'b110111100110;
   56884: result <= 12'b110111100110;
   56885: result <= 12'b110111100110;
   56886: result <= 12'b110111100110;
   56887: result <= 12'b110111100110;
   56888: result <= 12'b110111100110;
   56889: result <= 12'b110111100101;
   56890: result <= 12'b110111100101;
   56891: result <= 12'b110111100101;
   56892: result <= 12'b110111100101;
   56893: result <= 12'b110111100101;
   56894: result <= 12'b110111100101;
   56895: result <= 12'b110111100101;
   56896: result <= 12'b110111100101;
   56897: result <= 12'b110111100100;
   56898: result <= 12'b110111100100;
   56899: result <= 12'b110111100100;
   56900: result <= 12'b110111100100;
   56901: result <= 12'b110111100100;
   56902: result <= 12'b110111100100;
   56903: result <= 12'b110111100100;
   56904: result <= 12'b110111100011;
   56905: result <= 12'b110111100011;
   56906: result <= 12'b110111100011;
   56907: result <= 12'b110111100011;
   56908: result <= 12'b110111100011;
   56909: result <= 12'b110111100011;
   56910: result <= 12'b110111100011;
   56911: result <= 12'b110111100011;
   56912: result <= 12'b110111100010;
   56913: result <= 12'b110111100010;
   56914: result <= 12'b110111100010;
   56915: result <= 12'b110111100010;
   56916: result <= 12'b110111100010;
   56917: result <= 12'b110111100010;
   56918: result <= 12'b110111100010;
   56919: result <= 12'b110111100001;
   56920: result <= 12'b110111100001;
   56921: result <= 12'b110111100001;
   56922: result <= 12'b110111100001;
   56923: result <= 12'b110111100001;
   56924: result <= 12'b110111100001;
   56925: result <= 12'b110111100001;
   56926: result <= 12'b110111100001;
   56927: result <= 12'b110111100000;
   56928: result <= 12'b110111100000;
   56929: result <= 12'b110111100000;
   56930: result <= 12'b110111100000;
   56931: result <= 12'b110111100000;
   56932: result <= 12'b110111100000;
   56933: result <= 12'b110111100000;
   56934: result <= 12'b110111011111;
   56935: result <= 12'b110111011111;
   56936: result <= 12'b110111011111;
   56937: result <= 12'b110111011111;
   56938: result <= 12'b110111011111;
   56939: result <= 12'b110111011111;
   56940: result <= 12'b110111011111;
   56941: result <= 12'b110111011111;
   56942: result <= 12'b110111011110;
   56943: result <= 12'b110111011110;
   56944: result <= 12'b110111011110;
   56945: result <= 12'b110111011110;
   56946: result <= 12'b110111011110;
   56947: result <= 12'b110111011110;
   56948: result <= 12'b110111011110;
   56949: result <= 12'b110111011101;
   56950: result <= 12'b110111011101;
   56951: result <= 12'b110111011101;
   56952: result <= 12'b110111011101;
   56953: result <= 12'b110111011101;
   56954: result <= 12'b110111011101;
   56955: result <= 12'b110111011101;
   56956: result <= 12'b110111011101;
   56957: result <= 12'b110111011100;
   56958: result <= 12'b110111011100;
   56959: result <= 12'b110111011100;
   56960: result <= 12'b110111011100;
   56961: result <= 12'b110111011100;
   56962: result <= 12'b110111011100;
   56963: result <= 12'b110111011100;
   56964: result <= 12'b110111011011;
   56965: result <= 12'b110111011011;
   56966: result <= 12'b110111011011;
   56967: result <= 12'b110111011011;
   56968: result <= 12'b110111011011;
   56969: result <= 12'b110111011011;
   56970: result <= 12'b110111011011;
   56971: result <= 12'b110111011011;
   56972: result <= 12'b110111011010;
   56973: result <= 12'b110111011010;
   56974: result <= 12'b110111011010;
   56975: result <= 12'b110111011010;
   56976: result <= 12'b110111011010;
   56977: result <= 12'b110111011010;
   56978: result <= 12'b110111011010;
   56979: result <= 12'b110111011001;
   56980: result <= 12'b110111011001;
   56981: result <= 12'b110111011001;
   56982: result <= 12'b110111011001;
   56983: result <= 12'b110111011001;
   56984: result <= 12'b110111011001;
   56985: result <= 12'b110111011001;
   56986: result <= 12'b110111011000;
   56987: result <= 12'b110111011000;
   56988: result <= 12'b110111011000;
   56989: result <= 12'b110111011000;
   56990: result <= 12'b110111011000;
   56991: result <= 12'b110111011000;
   56992: result <= 12'b110111011000;
   56993: result <= 12'b110111011000;
   56994: result <= 12'b110111010111;
   56995: result <= 12'b110111010111;
   56996: result <= 12'b110111010111;
   56997: result <= 12'b110111010111;
   56998: result <= 12'b110111010111;
   56999: result <= 12'b110111010111;
   57000: result <= 12'b110111010111;
   57001: result <= 12'b110111010110;
   57002: result <= 12'b110111010110;
   57003: result <= 12'b110111010110;
   57004: result <= 12'b110111010110;
   57005: result <= 12'b110111010110;
   57006: result <= 12'b110111010110;
   57007: result <= 12'b110111010110;
   57008: result <= 12'b110111010110;
   57009: result <= 12'b110111010101;
   57010: result <= 12'b110111010101;
   57011: result <= 12'b110111010101;
   57012: result <= 12'b110111010101;
   57013: result <= 12'b110111010101;
   57014: result <= 12'b110111010101;
   57015: result <= 12'b110111010101;
   57016: result <= 12'b110111010100;
   57017: result <= 12'b110111010100;
   57018: result <= 12'b110111010100;
   57019: result <= 12'b110111010100;
   57020: result <= 12'b110111010100;
   57021: result <= 12'b110111010100;
   57022: result <= 12'b110111010100;
   57023: result <= 12'b110111010100;
   57024: result <= 12'b110111010011;
   57025: result <= 12'b110111010011;
   57026: result <= 12'b110111010011;
   57027: result <= 12'b110111010011;
   57028: result <= 12'b110111010011;
   57029: result <= 12'b110111010011;
   57030: result <= 12'b110111010011;
   57031: result <= 12'b110111010010;
   57032: result <= 12'b110111010010;
   57033: result <= 12'b110111010010;
   57034: result <= 12'b110111010010;
   57035: result <= 12'b110111010010;
   57036: result <= 12'b110111010010;
   57037: result <= 12'b110111010010;
   57038: result <= 12'b110111010010;
   57039: result <= 12'b110111010001;
   57040: result <= 12'b110111010001;
   57041: result <= 12'b110111010001;
   57042: result <= 12'b110111010001;
   57043: result <= 12'b110111010001;
   57044: result <= 12'b110111010001;
   57045: result <= 12'b110111010001;
   57046: result <= 12'b110111010000;
   57047: result <= 12'b110111010000;
   57048: result <= 12'b110111010000;
   57049: result <= 12'b110111010000;
   57050: result <= 12'b110111010000;
   57051: result <= 12'b110111010000;
   57052: result <= 12'b110111010000;
   57053: result <= 12'b110111001111;
   57054: result <= 12'b110111001111;
   57055: result <= 12'b110111001111;
   57056: result <= 12'b110111001111;
   57057: result <= 12'b110111001111;
   57058: result <= 12'b110111001111;
   57059: result <= 12'b110111001111;
   57060: result <= 12'b110111001111;
   57061: result <= 12'b110111001110;
   57062: result <= 12'b110111001110;
   57063: result <= 12'b110111001110;
   57064: result <= 12'b110111001110;
   57065: result <= 12'b110111001110;
   57066: result <= 12'b110111001110;
   57067: result <= 12'b110111001110;
   57068: result <= 12'b110111001101;
   57069: result <= 12'b110111001101;
   57070: result <= 12'b110111001101;
   57071: result <= 12'b110111001101;
   57072: result <= 12'b110111001101;
   57073: result <= 12'b110111001101;
   57074: result <= 12'b110111001101;
   57075: result <= 12'b110111001101;
   57076: result <= 12'b110111001100;
   57077: result <= 12'b110111001100;
   57078: result <= 12'b110111001100;
   57079: result <= 12'b110111001100;
   57080: result <= 12'b110111001100;
   57081: result <= 12'b110111001100;
   57082: result <= 12'b110111001100;
   57083: result <= 12'b110111001011;
   57084: result <= 12'b110111001011;
   57085: result <= 12'b110111001011;
   57086: result <= 12'b110111001011;
   57087: result <= 12'b110111001011;
   57088: result <= 12'b110111001011;
   57089: result <= 12'b110111001011;
   57090: result <= 12'b110111001010;
   57091: result <= 12'b110111001010;
   57092: result <= 12'b110111001010;
   57093: result <= 12'b110111001010;
   57094: result <= 12'b110111001010;
   57095: result <= 12'b110111001010;
   57096: result <= 12'b110111001010;
   57097: result <= 12'b110111001010;
   57098: result <= 12'b110111001001;
   57099: result <= 12'b110111001001;
   57100: result <= 12'b110111001001;
   57101: result <= 12'b110111001001;
   57102: result <= 12'b110111001001;
   57103: result <= 12'b110111001001;
   57104: result <= 12'b110111001001;
   57105: result <= 12'b110111001000;
   57106: result <= 12'b110111001000;
   57107: result <= 12'b110111001000;
   57108: result <= 12'b110111001000;
   57109: result <= 12'b110111001000;
   57110: result <= 12'b110111001000;
   57111: result <= 12'b110111001000;
   57112: result <= 12'b110111001000;
   57113: result <= 12'b110111000111;
   57114: result <= 12'b110111000111;
   57115: result <= 12'b110111000111;
   57116: result <= 12'b110111000111;
   57117: result <= 12'b110111000111;
   57118: result <= 12'b110111000111;
   57119: result <= 12'b110111000111;
   57120: result <= 12'b110111000110;
   57121: result <= 12'b110111000110;
   57122: result <= 12'b110111000110;
   57123: result <= 12'b110111000110;
   57124: result <= 12'b110111000110;
   57125: result <= 12'b110111000110;
   57126: result <= 12'b110111000110;
   57127: result <= 12'b110111000101;
   57128: result <= 12'b110111000101;
   57129: result <= 12'b110111000101;
   57130: result <= 12'b110111000101;
   57131: result <= 12'b110111000101;
   57132: result <= 12'b110111000101;
   57133: result <= 12'b110111000101;
   57134: result <= 12'b110111000101;
   57135: result <= 12'b110111000100;
   57136: result <= 12'b110111000100;
   57137: result <= 12'b110111000100;
   57138: result <= 12'b110111000100;
   57139: result <= 12'b110111000100;
   57140: result <= 12'b110111000100;
   57141: result <= 12'b110111000100;
   57142: result <= 12'b110111000011;
   57143: result <= 12'b110111000011;
   57144: result <= 12'b110111000011;
   57145: result <= 12'b110111000011;
   57146: result <= 12'b110111000011;
   57147: result <= 12'b110111000011;
   57148: result <= 12'b110111000011;
   57149: result <= 12'b110111000010;
   57150: result <= 12'b110111000010;
   57151: result <= 12'b110111000010;
   57152: result <= 12'b110111000010;
   57153: result <= 12'b110111000010;
   57154: result <= 12'b110111000010;
   57155: result <= 12'b110111000010;
   57156: result <= 12'b110111000010;
   57157: result <= 12'b110111000001;
   57158: result <= 12'b110111000001;
   57159: result <= 12'b110111000001;
   57160: result <= 12'b110111000001;
   57161: result <= 12'b110111000001;
   57162: result <= 12'b110111000001;
   57163: result <= 12'b110111000001;
   57164: result <= 12'b110111000000;
   57165: result <= 12'b110111000000;
   57166: result <= 12'b110111000000;
   57167: result <= 12'b110111000000;
   57168: result <= 12'b110111000000;
   57169: result <= 12'b110111000000;
   57170: result <= 12'b110111000000;
   57171: result <= 12'b110110111111;
   57172: result <= 12'b110110111111;
   57173: result <= 12'b110110111111;
   57174: result <= 12'b110110111111;
   57175: result <= 12'b110110111111;
   57176: result <= 12'b110110111111;
   57177: result <= 12'b110110111111;
   57178: result <= 12'b110110111111;
   57179: result <= 12'b110110111110;
   57180: result <= 12'b110110111110;
   57181: result <= 12'b110110111110;
   57182: result <= 12'b110110111110;
   57183: result <= 12'b110110111110;
   57184: result <= 12'b110110111110;
   57185: result <= 12'b110110111110;
   57186: result <= 12'b110110111101;
   57187: result <= 12'b110110111101;
   57188: result <= 12'b110110111101;
   57189: result <= 12'b110110111101;
   57190: result <= 12'b110110111101;
   57191: result <= 12'b110110111101;
   57192: result <= 12'b110110111101;
   57193: result <= 12'b110110111100;
   57194: result <= 12'b110110111100;
   57195: result <= 12'b110110111100;
   57196: result <= 12'b110110111100;
   57197: result <= 12'b110110111100;
   57198: result <= 12'b110110111100;
   57199: result <= 12'b110110111100;
   57200: result <= 12'b110110111100;
   57201: result <= 12'b110110111011;
   57202: result <= 12'b110110111011;
   57203: result <= 12'b110110111011;
   57204: result <= 12'b110110111011;
   57205: result <= 12'b110110111011;
   57206: result <= 12'b110110111011;
   57207: result <= 12'b110110111011;
   57208: result <= 12'b110110111010;
   57209: result <= 12'b110110111010;
   57210: result <= 12'b110110111010;
   57211: result <= 12'b110110111010;
   57212: result <= 12'b110110111010;
   57213: result <= 12'b110110111010;
   57214: result <= 12'b110110111010;
   57215: result <= 12'b110110111001;
   57216: result <= 12'b110110111001;
   57217: result <= 12'b110110111001;
   57218: result <= 12'b110110111001;
   57219: result <= 12'b110110111001;
   57220: result <= 12'b110110111001;
   57221: result <= 12'b110110111001;
   57222: result <= 12'b110110111000;
   57223: result <= 12'b110110111000;
   57224: result <= 12'b110110111000;
   57225: result <= 12'b110110111000;
   57226: result <= 12'b110110111000;
   57227: result <= 12'b110110111000;
   57228: result <= 12'b110110111000;
   57229: result <= 12'b110110111000;
   57230: result <= 12'b110110110111;
   57231: result <= 12'b110110110111;
   57232: result <= 12'b110110110111;
   57233: result <= 12'b110110110111;
   57234: result <= 12'b110110110111;
   57235: result <= 12'b110110110111;
   57236: result <= 12'b110110110111;
   57237: result <= 12'b110110110110;
   57238: result <= 12'b110110110110;
   57239: result <= 12'b110110110110;
   57240: result <= 12'b110110110110;
   57241: result <= 12'b110110110110;
   57242: result <= 12'b110110110110;
   57243: result <= 12'b110110110110;
   57244: result <= 12'b110110110101;
   57245: result <= 12'b110110110101;
   57246: result <= 12'b110110110101;
   57247: result <= 12'b110110110101;
   57248: result <= 12'b110110110101;
   57249: result <= 12'b110110110101;
   57250: result <= 12'b110110110101;
   57251: result <= 12'b110110110101;
   57252: result <= 12'b110110110100;
   57253: result <= 12'b110110110100;
   57254: result <= 12'b110110110100;
   57255: result <= 12'b110110110100;
   57256: result <= 12'b110110110100;
   57257: result <= 12'b110110110100;
   57258: result <= 12'b110110110100;
   57259: result <= 12'b110110110011;
   57260: result <= 12'b110110110011;
   57261: result <= 12'b110110110011;
   57262: result <= 12'b110110110011;
   57263: result <= 12'b110110110011;
   57264: result <= 12'b110110110011;
   57265: result <= 12'b110110110011;
   57266: result <= 12'b110110110010;
   57267: result <= 12'b110110110010;
   57268: result <= 12'b110110110010;
   57269: result <= 12'b110110110010;
   57270: result <= 12'b110110110010;
   57271: result <= 12'b110110110010;
   57272: result <= 12'b110110110010;
   57273: result <= 12'b110110110001;
   57274: result <= 12'b110110110001;
   57275: result <= 12'b110110110001;
   57276: result <= 12'b110110110001;
   57277: result <= 12'b110110110001;
   57278: result <= 12'b110110110001;
   57279: result <= 12'b110110110001;
   57280: result <= 12'b110110110001;
   57281: result <= 12'b110110110000;
   57282: result <= 12'b110110110000;
   57283: result <= 12'b110110110000;
   57284: result <= 12'b110110110000;
   57285: result <= 12'b110110110000;
   57286: result <= 12'b110110110000;
   57287: result <= 12'b110110110000;
   57288: result <= 12'b110110101111;
   57289: result <= 12'b110110101111;
   57290: result <= 12'b110110101111;
   57291: result <= 12'b110110101111;
   57292: result <= 12'b110110101111;
   57293: result <= 12'b110110101111;
   57294: result <= 12'b110110101111;
   57295: result <= 12'b110110101110;
   57296: result <= 12'b110110101110;
   57297: result <= 12'b110110101110;
   57298: result <= 12'b110110101110;
   57299: result <= 12'b110110101110;
   57300: result <= 12'b110110101110;
   57301: result <= 12'b110110101110;
   57302: result <= 12'b110110101101;
   57303: result <= 12'b110110101101;
   57304: result <= 12'b110110101101;
   57305: result <= 12'b110110101101;
   57306: result <= 12'b110110101101;
   57307: result <= 12'b110110101101;
   57308: result <= 12'b110110101101;
   57309: result <= 12'b110110101101;
   57310: result <= 12'b110110101100;
   57311: result <= 12'b110110101100;
   57312: result <= 12'b110110101100;
   57313: result <= 12'b110110101100;
   57314: result <= 12'b110110101100;
   57315: result <= 12'b110110101100;
   57316: result <= 12'b110110101100;
   57317: result <= 12'b110110101011;
   57318: result <= 12'b110110101011;
   57319: result <= 12'b110110101011;
   57320: result <= 12'b110110101011;
   57321: result <= 12'b110110101011;
   57322: result <= 12'b110110101011;
   57323: result <= 12'b110110101011;
   57324: result <= 12'b110110101010;
   57325: result <= 12'b110110101010;
   57326: result <= 12'b110110101010;
   57327: result <= 12'b110110101010;
   57328: result <= 12'b110110101010;
   57329: result <= 12'b110110101010;
   57330: result <= 12'b110110101010;
   57331: result <= 12'b110110101001;
   57332: result <= 12'b110110101001;
   57333: result <= 12'b110110101001;
   57334: result <= 12'b110110101001;
   57335: result <= 12'b110110101001;
   57336: result <= 12'b110110101001;
   57337: result <= 12'b110110101001;
   57338: result <= 12'b110110101000;
   57339: result <= 12'b110110101000;
   57340: result <= 12'b110110101000;
   57341: result <= 12'b110110101000;
   57342: result <= 12'b110110101000;
   57343: result <= 12'b110110101000;
   57344: result <= 12'b110110101000;
   57345: result <= 12'b110110101000;
   57346: result <= 12'b110110100111;
   57347: result <= 12'b110110100111;
   57348: result <= 12'b110110100111;
   57349: result <= 12'b110110100111;
   57350: result <= 12'b110110100111;
   57351: result <= 12'b110110100111;
   57352: result <= 12'b110110100111;
   57353: result <= 12'b110110100110;
   57354: result <= 12'b110110100110;
   57355: result <= 12'b110110100110;
   57356: result <= 12'b110110100110;
   57357: result <= 12'b110110100110;
   57358: result <= 12'b110110100110;
   57359: result <= 12'b110110100110;
   57360: result <= 12'b110110100101;
   57361: result <= 12'b110110100101;
   57362: result <= 12'b110110100101;
   57363: result <= 12'b110110100101;
   57364: result <= 12'b110110100101;
   57365: result <= 12'b110110100101;
   57366: result <= 12'b110110100101;
   57367: result <= 12'b110110100100;
   57368: result <= 12'b110110100100;
   57369: result <= 12'b110110100100;
   57370: result <= 12'b110110100100;
   57371: result <= 12'b110110100100;
   57372: result <= 12'b110110100100;
   57373: result <= 12'b110110100100;
   57374: result <= 12'b110110100011;
   57375: result <= 12'b110110100011;
   57376: result <= 12'b110110100011;
   57377: result <= 12'b110110100011;
   57378: result <= 12'b110110100011;
   57379: result <= 12'b110110100011;
   57380: result <= 12'b110110100011;
   57381: result <= 12'b110110100011;
   57382: result <= 12'b110110100010;
   57383: result <= 12'b110110100010;
   57384: result <= 12'b110110100010;
   57385: result <= 12'b110110100010;
   57386: result <= 12'b110110100010;
   57387: result <= 12'b110110100010;
   57388: result <= 12'b110110100010;
   57389: result <= 12'b110110100001;
   57390: result <= 12'b110110100001;
   57391: result <= 12'b110110100001;
   57392: result <= 12'b110110100001;
   57393: result <= 12'b110110100001;
   57394: result <= 12'b110110100001;
   57395: result <= 12'b110110100001;
   57396: result <= 12'b110110100000;
   57397: result <= 12'b110110100000;
   57398: result <= 12'b110110100000;
   57399: result <= 12'b110110100000;
   57400: result <= 12'b110110100000;
   57401: result <= 12'b110110100000;
   57402: result <= 12'b110110100000;
   57403: result <= 12'b110110011111;
   57404: result <= 12'b110110011111;
   57405: result <= 12'b110110011111;
   57406: result <= 12'b110110011111;
   57407: result <= 12'b110110011111;
   57408: result <= 12'b110110011111;
   57409: result <= 12'b110110011111;
   57410: result <= 12'b110110011110;
   57411: result <= 12'b110110011110;
   57412: result <= 12'b110110011110;
   57413: result <= 12'b110110011110;
   57414: result <= 12'b110110011110;
   57415: result <= 12'b110110011110;
   57416: result <= 12'b110110011110;
   57417: result <= 12'b110110011101;
   57418: result <= 12'b110110011101;
   57419: result <= 12'b110110011101;
   57420: result <= 12'b110110011101;
   57421: result <= 12'b110110011101;
   57422: result <= 12'b110110011101;
   57423: result <= 12'b110110011101;
   57424: result <= 12'b110110011101;
   57425: result <= 12'b110110011100;
   57426: result <= 12'b110110011100;
   57427: result <= 12'b110110011100;
   57428: result <= 12'b110110011100;
   57429: result <= 12'b110110011100;
   57430: result <= 12'b110110011100;
   57431: result <= 12'b110110011100;
   57432: result <= 12'b110110011011;
   57433: result <= 12'b110110011011;
   57434: result <= 12'b110110011011;
   57435: result <= 12'b110110011011;
   57436: result <= 12'b110110011011;
   57437: result <= 12'b110110011011;
   57438: result <= 12'b110110011011;
   57439: result <= 12'b110110011010;
   57440: result <= 12'b110110011010;
   57441: result <= 12'b110110011010;
   57442: result <= 12'b110110011010;
   57443: result <= 12'b110110011010;
   57444: result <= 12'b110110011010;
   57445: result <= 12'b110110011010;
   57446: result <= 12'b110110011001;
   57447: result <= 12'b110110011001;
   57448: result <= 12'b110110011001;
   57449: result <= 12'b110110011001;
   57450: result <= 12'b110110011001;
   57451: result <= 12'b110110011001;
   57452: result <= 12'b110110011001;
   57453: result <= 12'b110110011000;
   57454: result <= 12'b110110011000;
   57455: result <= 12'b110110011000;
   57456: result <= 12'b110110011000;
   57457: result <= 12'b110110011000;
   57458: result <= 12'b110110011000;
   57459: result <= 12'b110110011000;
   57460: result <= 12'b110110010111;
   57461: result <= 12'b110110010111;
   57462: result <= 12'b110110010111;
   57463: result <= 12'b110110010111;
   57464: result <= 12'b110110010111;
   57465: result <= 12'b110110010111;
   57466: result <= 12'b110110010111;
   57467: result <= 12'b110110010110;
   57468: result <= 12'b110110010110;
   57469: result <= 12'b110110010110;
   57470: result <= 12'b110110010110;
   57471: result <= 12'b110110010110;
   57472: result <= 12'b110110010110;
   57473: result <= 12'b110110010110;
   57474: result <= 12'b110110010101;
   57475: result <= 12'b110110010101;
   57476: result <= 12'b110110010101;
   57477: result <= 12'b110110010101;
   57478: result <= 12'b110110010101;
   57479: result <= 12'b110110010101;
   57480: result <= 12'b110110010101;
   57481: result <= 12'b110110010101;
   57482: result <= 12'b110110010100;
   57483: result <= 12'b110110010100;
   57484: result <= 12'b110110010100;
   57485: result <= 12'b110110010100;
   57486: result <= 12'b110110010100;
   57487: result <= 12'b110110010100;
   57488: result <= 12'b110110010100;
   57489: result <= 12'b110110010011;
   57490: result <= 12'b110110010011;
   57491: result <= 12'b110110010011;
   57492: result <= 12'b110110010011;
   57493: result <= 12'b110110010011;
   57494: result <= 12'b110110010011;
   57495: result <= 12'b110110010011;
   57496: result <= 12'b110110010010;
   57497: result <= 12'b110110010010;
   57498: result <= 12'b110110010010;
   57499: result <= 12'b110110010010;
   57500: result <= 12'b110110010010;
   57501: result <= 12'b110110010010;
   57502: result <= 12'b110110010010;
   57503: result <= 12'b110110010001;
   57504: result <= 12'b110110010001;
   57505: result <= 12'b110110010001;
   57506: result <= 12'b110110010001;
   57507: result <= 12'b110110010001;
   57508: result <= 12'b110110010001;
   57509: result <= 12'b110110010001;
   57510: result <= 12'b110110010000;
   57511: result <= 12'b110110010000;
   57512: result <= 12'b110110010000;
   57513: result <= 12'b110110010000;
   57514: result <= 12'b110110010000;
   57515: result <= 12'b110110010000;
   57516: result <= 12'b110110010000;
   57517: result <= 12'b110110001111;
   57518: result <= 12'b110110001111;
   57519: result <= 12'b110110001111;
   57520: result <= 12'b110110001111;
   57521: result <= 12'b110110001111;
   57522: result <= 12'b110110001111;
   57523: result <= 12'b110110001111;
   57524: result <= 12'b110110001110;
   57525: result <= 12'b110110001110;
   57526: result <= 12'b110110001110;
   57527: result <= 12'b110110001110;
   57528: result <= 12'b110110001110;
   57529: result <= 12'b110110001110;
   57530: result <= 12'b110110001110;
   57531: result <= 12'b110110001101;
   57532: result <= 12'b110110001101;
   57533: result <= 12'b110110001101;
   57534: result <= 12'b110110001101;
   57535: result <= 12'b110110001101;
   57536: result <= 12'b110110001101;
   57537: result <= 12'b110110001101;
   57538: result <= 12'b110110001100;
   57539: result <= 12'b110110001100;
   57540: result <= 12'b110110001100;
   57541: result <= 12'b110110001100;
   57542: result <= 12'b110110001100;
   57543: result <= 12'b110110001100;
   57544: result <= 12'b110110001100;
   57545: result <= 12'b110110001011;
   57546: result <= 12'b110110001011;
   57547: result <= 12'b110110001011;
   57548: result <= 12'b110110001011;
   57549: result <= 12'b110110001011;
   57550: result <= 12'b110110001011;
   57551: result <= 12'b110110001011;
   57552: result <= 12'b110110001010;
   57553: result <= 12'b110110001010;
   57554: result <= 12'b110110001010;
   57555: result <= 12'b110110001010;
   57556: result <= 12'b110110001010;
   57557: result <= 12'b110110001010;
   57558: result <= 12'b110110001010;
   57559: result <= 12'b110110001001;
   57560: result <= 12'b110110001001;
   57561: result <= 12'b110110001001;
   57562: result <= 12'b110110001001;
   57563: result <= 12'b110110001001;
   57564: result <= 12'b110110001001;
   57565: result <= 12'b110110001001;
   57566: result <= 12'b110110001001;
   57567: result <= 12'b110110001000;
   57568: result <= 12'b110110001000;
   57569: result <= 12'b110110001000;
   57570: result <= 12'b110110001000;
   57571: result <= 12'b110110001000;
   57572: result <= 12'b110110001000;
   57573: result <= 12'b110110001000;
   57574: result <= 12'b110110000111;
   57575: result <= 12'b110110000111;
   57576: result <= 12'b110110000111;
   57577: result <= 12'b110110000111;
   57578: result <= 12'b110110000111;
   57579: result <= 12'b110110000111;
   57580: result <= 12'b110110000111;
   57581: result <= 12'b110110000110;
   57582: result <= 12'b110110000110;
   57583: result <= 12'b110110000110;
   57584: result <= 12'b110110000110;
   57585: result <= 12'b110110000110;
   57586: result <= 12'b110110000110;
   57587: result <= 12'b110110000110;
   57588: result <= 12'b110110000101;
   57589: result <= 12'b110110000101;
   57590: result <= 12'b110110000101;
   57591: result <= 12'b110110000101;
   57592: result <= 12'b110110000101;
   57593: result <= 12'b110110000101;
   57594: result <= 12'b110110000101;
   57595: result <= 12'b110110000100;
   57596: result <= 12'b110110000100;
   57597: result <= 12'b110110000100;
   57598: result <= 12'b110110000100;
   57599: result <= 12'b110110000100;
   57600: result <= 12'b110110000100;
   57601: result <= 12'b110110000100;
   57602: result <= 12'b110110000011;
   57603: result <= 12'b110110000011;
   57604: result <= 12'b110110000011;
   57605: result <= 12'b110110000011;
   57606: result <= 12'b110110000011;
   57607: result <= 12'b110110000011;
   57608: result <= 12'b110110000011;
   57609: result <= 12'b110110000010;
   57610: result <= 12'b110110000010;
   57611: result <= 12'b110110000010;
   57612: result <= 12'b110110000010;
   57613: result <= 12'b110110000010;
   57614: result <= 12'b110110000010;
   57615: result <= 12'b110110000010;
   57616: result <= 12'b110110000001;
   57617: result <= 12'b110110000001;
   57618: result <= 12'b110110000001;
   57619: result <= 12'b110110000001;
   57620: result <= 12'b110110000001;
   57621: result <= 12'b110110000001;
   57622: result <= 12'b110110000001;
   57623: result <= 12'b110110000000;
   57624: result <= 12'b110110000000;
   57625: result <= 12'b110110000000;
   57626: result <= 12'b110110000000;
   57627: result <= 12'b110110000000;
   57628: result <= 12'b110110000000;
   57629: result <= 12'b110110000000;
   57630: result <= 12'b110101111111;
   57631: result <= 12'b110101111111;
   57632: result <= 12'b110101111111;
   57633: result <= 12'b110101111111;
   57634: result <= 12'b110101111111;
   57635: result <= 12'b110101111111;
   57636: result <= 12'b110101111111;
   57637: result <= 12'b110101111110;
   57638: result <= 12'b110101111110;
   57639: result <= 12'b110101111110;
   57640: result <= 12'b110101111110;
   57641: result <= 12'b110101111110;
   57642: result <= 12'b110101111110;
   57643: result <= 12'b110101111110;
   57644: result <= 12'b110101111101;
   57645: result <= 12'b110101111101;
   57646: result <= 12'b110101111101;
   57647: result <= 12'b110101111101;
   57648: result <= 12'b110101111101;
   57649: result <= 12'b110101111101;
   57650: result <= 12'b110101111101;
   57651: result <= 12'b110101111100;
   57652: result <= 12'b110101111100;
   57653: result <= 12'b110101111100;
   57654: result <= 12'b110101111100;
   57655: result <= 12'b110101111100;
   57656: result <= 12'b110101111100;
   57657: result <= 12'b110101111100;
   57658: result <= 12'b110101111011;
   57659: result <= 12'b110101111011;
   57660: result <= 12'b110101111011;
   57661: result <= 12'b110101111011;
   57662: result <= 12'b110101111011;
   57663: result <= 12'b110101111011;
   57664: result <= 12'b110101111011;
   57665: result <= 12'b110101111010;
   57666: result <= 12'b110101111010;
   57667: result <= 12'b110101111010;
   57668: result <= 12'b110101111010;
   57669: result <= 12'b110101111010;
   57670: result <= 12'b110101111010;
   57671: result <= 12'b110101111010;
   57672: result <= 12'b110101111001;
   57673: result <= 12'b110101111001;
   57674: result <= 12'b110101111001;
   57675: result <= 12'b110101111001;
   57676: result <= 12'b110101111001;
   57677: result <= 12'b110101111001;
   57678: result <= 12'b110101111001;
   57679: result <= 12'b110101111000;
   57680: result <= 12'b110101111000;
   57681: result <= 12'b110101111000;
   57682: result <= 12'b110101111000;
   57683: result <= 12'b110101111000;
   57684: result <= 12'b110101111000;
   57685: result <= 12'b110101111000;
   57686: result <= 12'b110101110111;
   57687: result <= 12'b110101110111;
   57688: result <= 12'b110101110111;
   57689: result <= 12'b110101110111;
   57690: result <= 12'b110101110111;
   57691: result <= 12'b110101110111;
   57692: result <= 12'b110101110111;
   57693: result <= 12'b110101110110;
   57694: result <= 12'b110101110110;
   57695: result <= 12'b110101110110;
   57696: result <= 12'b110101110110;
   57697: result <= 12'b110101110110;
   57698: result <= 12'b110101110110;
   57699: result <= 12'b110101110110;
   57700: result <= 12'b110101110101;
   57701: result <= 12'b110101110101;
   57702: result <= 12'b110101110101;
   57703: result <= 12'b110101110101;
   57704: result <= 12'b110101110101;
   57705: result <= 12'b110101110101;
   57706: result <= 12'b110101110101;
   57707: result <= 12'b110101110100;
   57708: result <= 12'b110101110100;
   57709: result <= 12'b110101110100;
   57710: result <= 12'b110101110100;
   57711: result <= 12'b110101110100;
   57712: result <= 12'b110101110100;
   57713: result <= 12'b110101110100;
   57714: result <= 12'b110101110011;
   57715: result <= 12'b110101110011;
   57716: result <= 12'b110101110011;
   57717: result <= 12'b110101110011;
   57718: result <= 12'b110101110011;
   57719: result <= 12'b110101110011;
   57720: result <= 12'b110101110011;
   57721: result <= 12'b110101110010;
   57722: result <= 12'b110101110010;
   57723: result <= 12'b110101110010;
   57724: result <= 12'b110101110010;
   57725: result <= 12'b110101110010;
   57726: result <= 12'b110101110010;
   57727: result <= 12'b110101110010;
   57728: result <= 12'b110101110001;
   57729: result <= 12'b110101110001;
   57730: result <= 12'b110101110001;
   57731: result <= 12'b110101110001;
   57732: result <= 12'b110101110001;
   57733: result <= 12'b110101110001;
   57734: result <= 12'b110101110001;
   57735: result <= 12'b110101110000;
   57736: result <= 12'b110101110000;
   57737: result <= 12'b110101110000;
   57738: result <= 12'b110101110000;
   57739: result <= 12'b110101110000;
   57740: result <= 12'b110101110000;
   57741: result <= 12'b110101101111;
   57742: result <= 12'b110101101111;
   57743: result <= 12'b110101101111;
   57744: result <= 12'b110101101111;
   57745: result <= 12'b110101101111;
   57746: result <= 12'b110101101111;
   57747: result <= 12'b110101101111;
   57748: result <= 12'b110101101110;
   57749: result <= 12'b110101101110;
   57750: result <= 12'b110101101110;
   57751: result <= 12'b110101101110;
   57752: result <= 12'b110101101110;
   57753: result <= 12'b110101101110;
   57754: result <= 12'b110101101110;
   57755: result <= 12'b110101101101;
   57756: result <= 12'b110101101101;
   57757: result <= 12'b110101101101;
   57758: result <= 12'b110101101101;
   57759: result <= 12'b110101101101;
   57760: result <= 12'b110101101101;
   57761: result <= 12'b110101101101;
   57762: result <= 12'b110101101100;
   57763: result <= 12'b110101101100;
   57764: result <= 12'b110101101100;
   57765: result <= 12'b110101101100;
   57766: result <= 12'b110101101100;
   57767: result <= 12'b110101101100;
   57768: result <= 12'b110101101100;
   57769: result <= 12'b110101101011;
   57770: result <= 12'b110101101011;
   57771: result <= 12'b110101101011;
   57772: result <= 12'b110101101011;
   57773: result <= 12'b110101101011;
   57774: result <= 12'b110101101011;
   57775: result <= 12'b110101101011;
   57776: result <= 12'b110101101010;
   57777: result <= 12'b110101101010;
   57778: result <= 12'b110101101010;
   57779: result <= 12'b110101101010;
   57780: result <= 12'b110101101010;
   57781: result <= 12'b110101101010;
   57782: result <= 12'b110101101010;
   57783: result <= 12'b110101101001;
   57784: result <= 12'b110101101001;
   57785: result <= 12'b110101101001;
   57786: result <= 12'b110101101001;
   57787: result <= 12'b110101101001;
   57788: result <= 12'b110101101001;
   57789: result <= 12'b110101101001;
   57790: result <= 12'b110101101000;
   57791: result <= 12'b110101101000;
   57792: result <= 12'b110101101000;
   57793: result <= 12'b110101101000;
   57794: result <= 12'b110101101000;
   57795: result <= 12'b110101101000;
   57796: result <= 12'b110101101000;
   57797: result <= 12'b110101100111;
   57798: result <= 12'b110101100111;
   57799: result <= 12'b110101100111;
   57800: result <= 12'b110101100111;
   57801: result <= 12'b110101100111;
   57802: result <= 12'b110101100111;
   57803: result <= 12'b110101100111;
   57804: result <= 12'b110101100110;
   57805: result <= 12'b110101100110;
   57806: result <= 12'b110101100110;
   57807: result <= 12'b110101100110;
   57808: result <= 12'b110101100110;
   57809: result <= 12'b110101100110;
   57810: result <= 12'b110101100110;
   57811: result <= 12'b110101100101;
   57812: result <= 12'b110101100101;
   57813: result <= 12'b110101100101;
   57814: result <= 12'b110101100101;
   57815: result <= 12'b110101100101;
   57816: result <= 12'b110101100101;
   57817: result <= 12'b110101100101;
   57818: result <= 12'b110101100100;
   57819: result <= 12'b110101100100;
   57820: result <= 12'b110101100100;
   57821: result <= 12'b110101100100;
   57822: result <= 12'b110101100100;
   57823: result <= 12'b110101100100;
   57824: result <= 12'b110101100100;
   57825: result <= 12'b110101100011;
   57826: result <= 12'b110101100011;
   57827: result <= 12'b110101100011;
   57828: result <= 12'b110101100011;
   57829: result <= 12'b110101100011;
   57830: result <= 12'b110101100011;
   57831: result <= 12'b110101100010;
   57832: result <= 12'b110101100010;
   57833: result <= 12'b110101100010;
   57834: result <= 12'b110101100010;
   57835: result <= 12'b110101100010;
   57836: result <= 12'b110101100010;
   57837: result <= 12'b110101100010;
   57838: result <= 12'b110101100001;
   57839: result <= 12'b110101100001;
   57840: result <= 12'b110101100001;
   57841: result <= 12'b110101100001;
   57842: result <= 12'b110101100001;
   57843: result <= 12'b110101100001;
   57844: result <= 12'b110101100001;
   57845: result <= 12'b110101100000;
   57846: result <= 12'b110101100000;
   57847: result <= 12'b110101100000;
   57848: result <= 12'b110101100000;
   57849: result <= 12'b110101100000;
   57850: result <= 12'b110101100000;
   57851: result <= 12'b110101100000;
   57852: result <= 12'b110101011111;
   57853: result <= 12'b110101011111;
   57854: result <= 12'b110101011111;
   57855: result <= 12'b110101011111;
   57856: result <= 12'b110101011111;
   57857: result <= 12'b110101011111;
   57858: result <= 12'b110101011111;
   57859: result <= 12'b110101011110;
   57860: result <= 12'b110101011110;
   57861: result <= 12'b110101011110;
   57862: result <= 12'b110101011110;
   57863: result <= 12'b110101011110;
   57864: result <= 12'b110101011110;
   57865: result <= 12'b110101011110;
   57866: result <= 12'b110101011101;
   57867: result <= 12'b110101011101;
   57868: result <= 12'b110101011101;
   57869: result <= 12'b110101011101;
   57870: result <= 12'b110101011101;
   57871: result <= 12'b110101011101;
   57872: result <= 12'b110101011101;
   57873: result <= 12'b110101011100;
   57874: result <= 12'b110101011100;
   57875: result <= 12'b110101011100;
   57876: result <= 12'b110101011100;
   57877: result <= 12'b110101011100;
   57878: result <= 12'b110101011100;
   57879: result <= 12'b110101011100;
   57880: result <= 12'b110101011011;
   57881: result <= 12'b110101011011;
   57882: result <= 12'b110101011011;
   57883: result <= 12'b110101011011;
   57884: result <= 12'b110101011011;
   57885: result <= 12'b110101011011;
   57886: result <= 12'b110101011010;
   57887: result <= 12'b110101011010;
   57888: result <= 12'b110101011010;
   57889: result <= 12'b110101011010;
   57890: result <= 12'b110101011010;
   57891: result <= 12'b110101011010;
   57892: result <= 12'b110101011010;
   57893: result <= 12'b110101011001;
   57894: result <= 12'b110101011001;
   57895: result <= 12'b110101011001;
   57896: result <= 12'b110101011001;
   57897: result <= 12'b110101011001;
   57898: result <= 12'b110101011001;
   57899: result <= 12'b110101011001;
   57900: result <= 12'b110101011000;
   57901: result <= 12'b110101011000;
   57902: result <= 12'b110101011000;
   57903: result <= 12'b110101011000;
   57904: result <= 12'b110101011000;
   57905: result <= 12'b110101011000;
   57906: result <= 12'b110101011000;
   57907: result <= 12'b110101010111;
   57908: result <= 12'b110101010111;
   57909: result <= 12'b110101010111;
   57910: result <= 12'b110101010111;
   57911: result <= 12'b110101010111;
   57912: result <= 12'b110101010111;
   57913: result <= 12'b110101010111;
   57914: result <= 12'b110101010110;
   57915: result <= 12'b110101010110;
   57916: result <= 12'b110101010110;
   57917: result <= 12'b110101010110;
   57918: result <= 12'b110101010110;
   57919: result <= 12'b110101010110;
   57920: result <= 12'b110101010110;
   57921: result <= 12'b110101010101;
   57922: result <= 12'b110101010101;
   57923: result <= 12'b110101010101;
   57924: result <= 12'b110101010101;
   57925: result <= 12'b110101010101;
   57926: result <= 12'b110101010101;
   57927: result <= 12'b110101010100;
   57928: result <= 12'b110101010100;
   57929: result <= 12'b110101010100;
   57930: result <= 12'b110101010100;
   57931: result <= 12'b110101010100;
   57932: result <= 12'b110101010100;
   57933: result <= 12'b110101010100;
   57934: result <= 12'b110101010011;
   57935: result <= 12'b110101010011;
   57936: result <= 12'b110101010011;
   57937: result <= 12'b110101010011;
   57938: result <= 12'b110101010011;
   57939: result <= 12'b110101010011;
   57940: result <= 12'b110101010011;
   57941: result <= 12'b110101010010;
   57942: result <= 12'b110101010010;
   57943: result <= 12'b110101010010;
   57944: result <= 12'b110101010010;
   57945: result <= 12'b110101010010;
   57946: result <= 12'b110101010010;
   57947: result <= 12'b110101010010;
   57948: result <= 12'b110101010001;
   57949: result <= 12'b110101010001;
   57950: result <= 12'b110101010001;
   57951: result <= 12'b110101010001;
   57952: result <= 12'b110101010001;
   57953: result <= 12'b110101010001;
   57954: result <= 12'b110101010001;
   57955: result <= 12'b110101010000;
   57956: result <= 12'b110101010000;
   57957: result <= 12'b110101010000;
   57958: result <= 12'b110101010000;
   57959: result <= 12'b110101010000;
   57960: result <= 12'b110101010000;
   57961: result <= 12'b110101010000;
   57962: result <= 12'b110101001111;
   57963: result <= 12'b110101001111;
   57964: result <= 12'b110101001111;
   57965: result <= 12'b110101001111;
   57966: result <= 12'b110101001111;
   57967: result <= 12'b110101001111;
   57968: result <= 12'b110101001110;
   57969: result <= 12'b110101001110;
   57970: result <= 12'b110101001110;
   57971: result <= 12'b110101001110;
   57972: result <= 12'b110101001110;
   57973: result <= 12'b110101001110;
   57974: result <= 12'b110101001110;
   57975: result <= 12'b110101001101;
   57976: result <= 12'b110101001101;
   57977: result <= 12'b110101001101;
   57978: result <= 12'b110101001101;
   57979: result <= 12'b110101001101;
   57980: result <= 12'b110101001101;
   57981: result <= 12'b110101001101;
   57982: result <= 12'b110101001100;
   57983: result <= 12'b110101001100;
   57984: result <= 12'b110101001100;
   57985: result <= 12'b110101001100;
   57986: result <= 12'b110101001100;
   57987: result <= 12'b110101001100;
   57988: result <= 12'b110101001100;
   57989: result <= 12'b110101001011;
   57990: result <= 12'b110101001011;
   57991: result <= 12'b110101001011;
   57992: result <= 12'b110101001011;
   57993: result <= 12'b110101001011;
   57994: result <= 12'b110101001011;
   57995: result <= 12'b110101001011;
   57996: result <= 12'b110101001010;
   57997: result <= 12'b110101001010;
   57998: result <= 12'b110101001010;
   57999: result <= 12'b110101001010;
   58000: result <= 12'b110101001010;
   58001: result <= 12'b110101001010;
   58002: result <= 12'b110101001001;
   58003: result <= 12'b110101001001;
   58004: result <= 12'b110101001001;
   58005: result <= 12'b110101001001;
   58006: result <= 12'b110101001001;
   58007: result <= 12'b110101001001;
   58008: result <= 12'b110101001001;
   58009: result <= 12'b110101001000;
   58010: result <= 12'b110101001000;
   58011: result <= 12'b110101001000;
   58012: result <= 12'b110101001000;
   58013: result <= 12'b110101001000;
   58014: result <= 12'b110101001000;
   58015: result <= 12'b110101001000;
   58016: result <= 12'b110101000111;
   58017: result <= 12'b110101000111;
   58018: result <= 12'b110101000111;
   58019: result <= 12'b110101000111;
   58020: result <= 12'b110101000111;
   58021: result <= 12'b110101000111;
   58022: result <= 12'b110101000111;
   58023: result <= 12'b110101000110;
   58024: result <= 12'b110101000110;
   58025: result <= 12'b110101000110;
   58026: result <= 12'b110101000110;
   58027: result <= 12'b110101000110;
   58028: result <= 12'b110101000110;
   58029: result <= 12'b110101000101;
   58030: result <= 12'b110101000101;
   58031: result <= 12'b110101000101;
   58032: result <= 12'b110101000101;
   58033: result <= 12'b110101000101;
   58034: result <= 12'b110101000101;
   58035: result <= 12'b110101000101;
   58036: result <= 12'b110101000100;
   58037: result <= 12'b110101000100;
   58038: result <= 12'b110101000100;
   58039: result <= 12'b110101000100;
   58040: result <= 12'b110101000100;
   58041: result <= 12'b110101000100;
   58042: result <= 12'b110101000100;
   58043: result <= 12'b110101000011;
   58044: result <= 12'b110101000011;
   58045: result <= 12'b110101000011;
   58046: result <= 12'b110101000011;
   58047: result <= 12'b110101000011;
   58048: result <= 12'b110101000011;
   58049: result <= 12'b110101000011;
   58050: result <= 12'b110101000010;
   58051: result <= 12'b110101000010;
   58052: result <= 12'b110101000010;
   58053: result <= 12'b110101000010;
   58054: result <= 12'b110101000010;
   58055: result <= 12'b110101000010;
   58056: result <= 12'b110101000010;
   58057: result <= 12'b110101000001;
   58058: result <= 12'b110101000001;
   58059: result <= 12'b110101000001;
   58060: result <= 12'b110101000001;
   58061: result <= 12'b110101000001;
   58062: result <= 12'b110101000001;
   58063: result <= 12'b110101000000;
   58064: result <= 12'b110101000000;
   58065: result <= 12'b110101000000;
   58066: result <= 12'b110101000000;
   58067: result <= 12'b110101000000;
   58068: result <= 12'b110101000000;
   58069: result <= 12'b110101000000;
   58070: result <= 12'b110100111111;
   58071: result <= 12'b110100111111;
   58072: result <= 12'b110100111111;
   58073: result <= 12'b110100111111;
   58074: result <= 12'b110100111111;
   58075: result <= 12'b110100111111;
   58076: result <= 12'b110100111111;
   58077: result <= 12'b110100111110;
   58078: result <= 12'b110100111110;
   58079: result <= 12'b110100111110;
   58080: result <= 12'b110100111110;
   58081: result <= 12'b110100111110;
   58082: result <= 12'b110100111110;
   58083: result <= 12'b110100111110;
   58084: result <= 12'b110100111101;
   58085: result <= 12'b110100111101;
   58086: result <= 12'b110100111101;
   58087: result <= 12'b110100111101;
   58088: result <= 12'b110100111101;
   58089: result <= 12'b110100111101;
   58090: result <= 12'b110100111100;
   58091: result <= 12'b110100111100;
   58092: result <= 12'b110100111100;
   58093: result <= 12'b110100111100;
   58094: result <= 12'b110100111100;
   58095: result <= 12'b110100111100;
   58096: result <= 12'b110100111100;
   58097: result <= 12'b110100111011;
   58098: result <= 12'b110100111011;
   58099: result <= 12'b110100111011;
   58100: result <= 12'b110100111011;
   58101: result <= 12'b110100111011;
   58102: result <= 12'b110100111011;
   58103: result <= 12'b110100111011;
   58104: result <= 12'b110100111010;
   58105: result <= 12'b110100111010;
   58106: result <= 12'b110100111010;
   58107: result <= 12'b110100111010;
   58108: result <= 12'b110100111010;
   58109: result <= 12'b110100111010;
   58110: result <= 12'b110100111001;
   58111: result <= 12'b110100111001;
   58112: result <= 12'b110100111001;
   58113: result <= 12'b110100111001;
   58114: result <= 12'b110100111001;
   58115: result <= 12'b110100111001;
   58116: result <= 12'b110100111001;
   58117: result <= 12'b110100111000;
   58118: result <= 12'b110100111000;
   58119: result <= 12'b110100111000;
   58120: result <= 12'b110100111000;
   58121: result <= 12'b110100111000;
   58122: result <= 12'b110100111000;
   58123: result <= 12'b110100111000;
   58124: result <= 12'b110100110111;
   58125: result <= 12'b110100110111;
   58126: result <= 12'b110100110111;
   58127: result <= 12'b110100110111;
   58128: result <= 12'b110100110111;
   58129: result <= 12'b110100110111;
   58130: result <= 12'b110100110111;
   58131: result <= 12'b110100110110;
   58132: result <= 12'b110100110110;
   58133: result <= 12'b110100110110;
   58134: result <= 12'b110100110110;
   58135: result <= 12'b110100110110;
   58136: result <= 12'b110100110110;
   58137: result <= 12'b110100110101;
   58138: result <= 12'b110100110101;
   58139: result <= 12'b110100110101;
   58140: result <= 12'b110100110101;
   58141: result <= 12'b110100110101;
   58142: result <= 12'b110100110101;
   58143: result <= 12'b110100110101;
   58144: result <= 12'b110100110100;
   58145: result <= 12'b110100110100;
   58146: result <= 12'b110100110100;
   58147: result <= 12'b110100110100;
   58148: result <= 12'b110100110100;
   58149: result <= 12'b110100110100;
   58150: result <= 12'b110100110100;
   58151: result <= 12'b110100110011;
   58152: result <= 12'b110100110011;
   58153: result <= 12'b110100110011;
   58154: result <= 12'b110100110011;
   58155: result <= 12'b110100110011;
   58156: result <= 12'b110100110011;
   58157: result <= 12'b110100110010;
   58158: result <= 12'b110100110010;
   58159: result <= 12'b110100110010;
   58160: result <= 12'b110100110010;
   58161: result <= 12'b110100110010;
   58162: result <= 12'b110100110010;
   58163: result <= 12'b110100110010;
   58164: result <= 12'b110100110001;
   58165: result <= 12'b110100110001;
   58166: result <= 12'b110100110001;
   58167: result <= 12'b110100110001;
   58168: result <= 12'b110100110001;
   58169: result <= 12'b110100110001;
   58170: result <= 12'b110100110001;
   58171: result <= 12'b110100110000;
   58172: result <= 12'b110100110000;
   58173: result <= 12'b110100110000;
   58174: result <= 12'b110100110000;
   58175: result <= 12'b110100110000;
   58176: result <= 12'b110100110000;
   58177: result <= 12'b110100110000;
   58178: result <= 12'b110100101111;
   58179: result <= 12'b110100101111;
   58180: result <= 12'b110100101111;
   58181: result <= 12'b110100101111;
   58182: result <= 12'b110100101111;
   58183: result <= 12'b110100101111;
   58184: result <= 12'b110100101110;
   58185: result <= 12'b110100101110;
   58186: result <= 12'b110100101110;
   58187: result <= 12'b110100101110;
   58188: result <= 12'b110100101110;
   58189: result <= 12'b110100101110;
   58190: result <= 12'b110100101110;
   58191: result <= 12'b110100101101;
   58192: result <= 12'b110100101101;
   58193: result <= 12'b110100101101;
   58194: result <= 12'b110100101101;
   58195: result <= 12'b110100101101;
   58196: result <= 12'b110100101101;
   58197: result <= 12'b110100101101;
   58198: result <= 12'b110100101100;
   58199: result <= 12'b110100101100;
   58200: result <= 12'b110100101100;
   58201: result <= 12'b110100101100;
   58202: result <= 12'b110100101100;
   58203: result <= 12'b110100101100;
   58204: result <= 12'b110100101011;
   58205: result <= 12'b110100101011;
   58206: result <= 12'b110100101011;
   58207: result <= 12'b110100101011;
   58208: result <= 12'b110100101011;
   58209: result <= 12'b110100101011;
   58210: result <= 12'b110100101011;
   58211: result <= 12'b110100101010;
   58212: result <= 12'b110100101010;
   58213: result <= 12'b110100101010;
   58214: result <= 12'b110100101010;
   58215: result <= 12'b110100101010;
   58216: result <= 12'b110100101010;
   58217: result <= 12'b110100101010;
   58218: result <= 12'b110100101001;
   58219: result <= 12'b110100101001;
   58220: result <= 12'b110100101001;
   58221: result <= 12'b110100101001;
   58222: result <= 12'b110100101001;
   58223: result <= 12'b110100101001;
   58224: result <= 12'b110100101000;
   58225: result <= 12'b110100101000;
   58226: result <= 12'b110100101000;
   58227: result <= 12'b110100101000;
   58228: result <= 12'b110100101000;
   58229: result <= 12'b110100101000;
   58230: result <= 12'b110100101000;
   58231: result <= 12'b110100100111;
   58232: result <= 12'b110100100111;
   58233: result <= 12'b110100100111;
   58234: result <= 12'b110100100111;
   58235: result <= 12'b110100100111;
   58236: result <= 12'b110100100111;
   58237: result <= 12'b110100100111;
   58238: result <= 12'b110100100110;
   58239: result <= 12'b110100100110;
   58240: result <= 12'b110100100110;
   58241: result <= 12'b110100100110;
   58242: result <= 12'b110100100110;
   58243: result <= 12'b110100100110;
   58244: result <= 12'b110100100101;
   58245: result <= 12'b110100100101;
   58246: result <= 12'b110100100101;
   58247: result <= 12'b110100100101;
   58248: result <= 12'b110100100101;
   58249: result <= 12'b110100100101;
   58250: result <= 12'b110100100101;
   58251: result <= 12'b110100100100;
   58252: result <= 12'b110100100100;
   58253: result <= 12'b110100100100;
   58254: result <= 12'b110100100100;
   58255: result <= 12'b110100100100;
   58256: result <= 12'b110100100100;
   58257: result <= 12'b110100100100;
   58258: result <= 12'b110100100011;
   58259: result <= 12'b110100100011;
   58260: result <= 12'b110100100011;
   58261: result <= 12'b110100100011;
   58262: result <= 12'b110100100011;
   58263: result <= 12'b110100100011;
   58264: result <= 12'b110100100010;
   58265: result <= 12'b110100100010;
   58266: result <= 12'b110100100010;
   58267: result <= 12'b110100100010;
   58268: result <= 12'b110100100010;
   58269: result <= 12'b110100100010;
   58270: result <= 12'b110100100010;
   58271: result <= 12'b110100100001;
   58272: result <= 12'b110100100001;
   58273: result <= 12'b110100100001;
   58274: result <= 12'b110100100001;
   58275: result <= 12'b110100100001;
   58276: result <= 12'b110100100001;
   58277: result <= 12'b110100100000;
   58278: result <= 12'b110100100000;
   58279: result <= 12'b110100100000;
   58280: result <= 12'b110100100000;
   58281: result <= 12'b110100100000;
   58282: result <= 12'b110100100000;
   58283: result <= 12'b110100100000;
   58284: result <= 12'b110100011111;
   58285: result <= 12'b110100011111;
   58286: result <= 12'b110100011111;
   58287: result <= 12'b110100011111;
   58288: result <= 12'b110100011111;
   58289: result <= 12'b110100011111;
   58290: result <= 12'b110100011111;
   58291: result <= 12'b110100011110;
   58292: result <= 12'b110100011110;
   58293: result <= 12'b110100011110;
   58294: result <= 12'b110100011110;
   58295: result <= 12'b110100011110;
   58296: result <= 12'b110100011110;
   58297: result <= 12'b110100011101;
   58298: result <= 12'b110100011101;
   58299: result <= 12'b110100011101;
   58300: result <= 12'b110100011101;
   58301: result <= 12'b110100011101;
   58302: result <= 12'b110100011101;
   58303: result <= 12'b110100011101;
   58304: result <= 12'b110100011100;
   58305: result <= 12'b110100011100;
   58306: result <= 12'b110100011100;
   58307: result <= 12'b110100011100;
   58308: result <= 12'b110100011100;
   58309: result <= 12'b110100011100;
   58310: result <= 12'b110100011100;
   58311: result <= 12'b110100011011;
   58312: result <= 12'b110100011011;
   58313: result <= 12'b110100011011;
   58314: result <= 12'b110100011011;
   58315: result <= 12'b110100011011;
   58316: result <= 12'b110100011011;
   58317: result <= 12'b110100011010;
   58318: result <= 12'b110100011010;
   58319: result <= 12'b110100011010;
   58320: result <= 12'b110100011010;
   58321: result <= 12'b110100011010;
   58322: result <= 12'b110100011010;
   58323: result <= 12'b110100011010;
   58324: result <= 12'b110100011001;
   58325: result <= 12'b110100011001;
   58326: result <= 12'b110100011001;
   58327: result <= 12'b110100011001;
   58328: result <= 12'b110100011001;
   58329: result <= 12'b110100011001;
   58330: result <= 12'b110100011000;
   58331: result <= 12'b110100011000;
   58332: result <= 12'b110100011000;
   58333: result <= 12'b110100011000;
   58334: result <= 12'b110100011000;
   58335: result <= 12'b110100011000;
   58336: result <= 12'b110100011000;
   58337: result <= 12'b110100010111;
   58338: result <= 12'b110100010111;
   58339: result <= 12'b110100010111;
   58340: result <= 12'b110100010111;
   58341: result <= 12'b110100010111;
   58342: result <= 12'b110100010111;
   58343: result <= 12'b110100010111;
   58344: result <= 12'b110100010110;
   58345: result <= 12'b110100010110;
   58346: result <= 12'b110100010110;
   58347: result <= 12'b110100010110;
   58348: result <= 12'b110100010110;
   58349: result <= 12'b110100010110;
   58350: result <= 12'b110100010101;
   58351: result <= 12'b110100010101;
   58352: result <= 12'b110100010101;
   58353: result <= 12'b110100010101;
   58354: result <= 12'b110100010101;
   58355: result <= 12'b110100010101;
   58356: result <= 12'b110100010101;
   58357: result <= 12'b110100010100;
   58358: result <= 12'b110100010100;
   58359: result <= 12'b110100010100;
   58360: result <= 12'b110100010100;
   58361: result <= 12'b110100010100;
   58362: result <= 12'b110100010100;
   58363: result <= 12'b110100010011;
   58364: result <= 12'b110100010011;
   58365: result <= 12'b110100010011;
   58366: result <= 12'b110100010011;
   58367: result <= 12'b110100010011;
   58368: result <= 12'b110100010011;
   58369: result <= 12'b110100010011;
   58370: result <= 12'b110100010010;
   58371: result <= 12'b110100010010;
   58372: result <= 12'b110100010010;
   58373: result <= 12'b110100010010;
   58374: result <= 12'b110100010010;
   58375: result <= 12'b110100010010;
   58376: result <= 12'b110100010010;
   58377: result <= 12'b110100010001;
   58378: result <= 12'b110100010001;
   58379: result <= 12'b110100010001;
   58380: result <= 12'b110100010001;
   58381: result <= 12'b110100010001;
   58382: result <= 12'b110100010001;
   58383: result <= 12'b110100010000;
   58384: result <= 12'b110100010000;
   58385: result <= 12'b110100010000;
   58386: result <= 12'b110100010000;
   58387: result <= 12'b110100010000;
   58388: result <= 12'b110100010000;
   58389: result <= 12'b110100010000;
   58390: result <= 12'b110100001111;
   58391: result <= 12'b110100001111;
   58392: result <= 12'b110100001111;
   58393: result <= 12'b110100001111;
   58394: result <= 12'b110100001111;
   58395: result <= 12'b110100001111;
   58396: result <= 12'b110100001110;
   58397: result <= 12'b110100001110;
   58398: result <= 12'b110100001110;
   58399: result <= 12'b110100001110;
   58400: result <= 12'b110100001110;
   58401: result <= 12'b110100001110;
   58402: result <= 12'b110100001110;
   58403: result <= 12'b110100001101;
   58404: result <= 12'b110100001101;
   58405: result <= 12'b110100001101;
   58406: result <= 12'b110100001101;
   58407: result <= 12'b110100001101;
   58408: result <= 12'b110100001101;
   58409: result <= 12'b110100001101;
   58410: result <= 12'b110100001100;
   58411: result <= 12'b110100001100;
   58412: result <= 12'b110100001100;
   58413: result <= 12'b110100001100;
   58414: result <= 12'b110100001100;
   58415: result <= 12'b110100001100;
   58416: result <= 12'b110100001011;
   58417: result <= 12'b110100001011;
   58418: result <= 12'b110100001011;
   58419: result <= 12'b110100001011;
   58420: result <= 12'b110100001011;
   58421: result <= 12'b110100001011;
   58422: result <= 12'b110100001011;
   58423: result <= 12'b110100001010;
   58424: result <= 12'b110100001010;
   58425: result <= 12'b110100001010;
   58426: result <= 12'b110100001010;
   58427: result <= 12'b110100001010;
   58428: result <= 12'b110100001010;
   58429: result <= 12'b110100001001;
   58430: result <= 12'b110100001001;
   58431: result <= 12'b110100001001;
   58432: result <= 12'b110100001001;
   58433: result <= 12'b110100001001;
   58434: result <= 12'b110100001001;
   58435: result <= 12'b110100001001;
   58436: result <= 12'b110100001000;
   58437: result <= 12'b110100001000;
   58438: result <= 12'b110100001000;
   58439: result <= 12'b110100001000;
   58440: result <= 12'b110100001000;
   58441: result <= 12'b110100001000;
   58442: result <= 12'b110100000111;
   58443: result <= 12'b110100000111;
   58444: result <= 12'b110100000111;
   58445: result <= 12'b110100000111;
   58446: result <= 12'b110100000111;
   58447: result <= 12'b110100000111;
   58448: result <= 12'b110100000111;
   58449: result <= 12'b110100000110;
   58450: result <= 12'b110100000110;
   58451: result <= 12'b110100000110;
   58452: result <= 12'b110100000110;
   58453: result <= 12'b110100000110;
   58454: result <= 12'b110100000110;
   58455: result <= 12'b110100000101;
   58456: result <= 12'b110100000101;
   58457: result <= 12'b110100000101;
   58458: result <= 12'b110100000101;
   58459: result <= 12'b110100000101;
   58460: result <= 12'b110100000101;
   58461: result <= 12'b110100000101;
   58462: result <= 12'b110100000100;
   58463: result <= 12'b110100000100;
   58464: result <= 12'b110100000100;
   58465: result <= 12'b110100000100;
   58466: result <= 12'b110100000100;
   58467: result <= 12'b110100000100;
   58468: result <= 12'b110100000011;
   58469: result <= 12'b110100000011;
   58470: result <= 12'b110100000011;
   58471: result <= 12'b110100000011;
   58472: result <= 12'b110100000011;
   58473: result <= 12'b110100000011;
   58474: result <= 12'b110100000011;
   58475: result <= 12'b110100000010;
   58476: result <= 12'b110100000010;
   58477: result <= 12'b110100000010;
   58478: result <= 12'b110100000010;
   58479: result <= 12'b110100000010;
   58480: result <= 12'b110100000010;
   58481: result <= 12'b110100000010;
   58482: result <= 12'b110100000001;
   58483: result <= 12'b110100000001;
   58484: result <= 12'b110100000001;
   58485: result <= 12'b110100000001;
   58486: result <= 12'b110100000001;
   58487: result <= 12'b110100000001;
   58488: result <= 12'b110100000000;
   58489: result <= 12'b110100000000;
   58490: result <= 12'b110100000000;
   58491: result <= 12'b110100000000;
   58492: result <= 12'b110100000000;
   58493: result <= 12'b110100000000;
   58494: result <= 12'b110100000000;
   58495: result <= 12'b110011111111;
   58496: result <= 12'b110011111111;
   58497: result <= 12'b110011111111;
   58498: result <= 12'b110011111111;
   58499: result <= 12'b110011111111;
   58500: result <= 12'b110011111111;
   58501: result <= 12'b110011111110;
   58502: result <= 12'b110011111110;
   58503: result <= 12'b110011111110;
   58504: result <= 12'b110011111110;
   58505: result <= 12'b110011111110;
   58506: result <= 12'b110011111110;
   58507: result <= 12'b110011111110;
   58508: result <= 12'b110011111101;
   58509: result <= 12'b110011111101;
   58510: result <= 12'b110011111101;
   58511: result <= 12'b110011111101;
   58512: result <= 12'b110011111101;
   58513: result <= 12'b110011111101;
   58514: result <= 12'b110011111100;
   58515: result <= 12'b110011111100;
   58516: result <= 12'b110011111100;
   58517: result <= 12'b110011111100;
   58518: result <= 12'b110011111100;
   58519: result <= 12'b110011111100;
   58520: result <= 12'b110011111100;
   58521: result <= 12'b110011111011;
   58522: result <= 12'b110011111011;
   58523: result <= 12'b110011111011;
   58524: result <= 12'b110011111011;
   58525: result <= 12'b110011111011;
   58526: result <= 12'b110011111011;
   58527: result <= 12'b110011111010;
   58528: result <= 12'b110011111010;
   58529: result <= 12'b110011111010;
   58530: result <= 12'b110011111010;
   58531: result <= 12'b110011111010;
   58532: result <= 12'b110011111010;
   58533: result <= 12'b110011111010;
   58534: result <= 12'b110011111001;
   58535: result <= 12'b110011111001;
   58536: result <= 12'b110011111001;
   58537: result <= 12'b110011111001;
   58538: result <= 12'b110011111001;
   58539: result <= 12'b110011111001;
   58540: result <= 12'b110011111000;
   58541: result <= 12'b110011111000;
   58542: result <= 12'b110011111000;
   58543: result <= 12'b110011111000;
   58544: result <= 12'b110011111000;
   58545: result <= 12'b110011111000;
   58546: result <= 12'b110011111000;
   58547: result <= 12'b110011110111;
   58548: result <= 12'b110011110111;
   58549: result <= 12'b110011110111;
   58550: result <= 12'b110011110111;
   58551: result <= 12'b110011110111;
   58552: result <= 12'b110011110111;
   58553: result <= 12'b110011110110;
   58554: result <= 12'b110011110110;
   58555: result <= 12'b110011110110;
   58556: result <= 12'b110011110110;
   58557: result <= 12'b110011110110;
   58558: result <= 12'b110011110110;
   58559: result <= 12'b110011110110;
   58560: result <= 12'b110011110101;
   58561: result <= 12'b110011110101;
   58562: result <= 12'b110011110101;
   58563: result <= 12'b110011110101;
   58564: result <= 12'b110011110101;
   58565: result <= 12'b110011110101;
   58566: result <= 12'b110011110100;
   58567: result <= 12'b110011110100;
   58568: result <= 12'b110011110100;
   58569: result <= 12'b110011110100;
   58570: result <= 12'b110011110100;
   58571: result <= 12'b110011110100;
   58572: result <= 12'b110011110100;
   58573: result <= 12'b110011110011;
   58574: result <= 12'b110011110011;
   58575: result <= 12'b110011110011;
   58576: result <= 12'b110011110011;
   58577: result <= 12'b110011110011;
   58578: result <= 12'b110011110011;
   58579: result <= 12'b110011110010;
   58580: result <= 12'b110011110010;
   58581: result <= 12'b110011110010;
   58582: result <= 12'b110011110010;
   58583: result <= 12'b110011110010;
   58584: result <= 12'b110011110010;
   58585: result <= 12'b110011110010;
   58586: result <= 12'b110011110001;
   58587: result <= 12'b110011110001;
   58588: result <= 12'b110011110001;
   58589: result <= 12'b110011110001;
   58590: result <= 12'b110011110001;
   58591: result <= 12'b110011110001;
   58592: result <= 12'b110011110000;
   58593: result <= 12'b110011110000;
   58594: result <= 12'b110011110000;
   58595: result <= 12'b110011110000;
   58596: result <= 12'b110011110000;
   58597: result <= 12'b110011110000;
   58598: result <= 12'b110011110000;
   58599: result <= 12'b110011101111;
   58600: result <= 12'b110011101111;
   58601: result <= 12'b110011101111;
   58602: result <= 12'b110011101111;
   58603: result <= 12'b110011101111;
   58604: result <= 12'b110011101111;
   58605: result <= 12'b110011101110;
   58606: result <= 12'b110011101110;
   58607: result <= 12'b110011101110;
   58608: result <= 12'b110011101110;
   58609: result <= 12'b110011101110;
   58610: result <= 12'b110011101110;
   58611: result <= 12'b110011101110;
   58612: result <= 12'b110011101101;
   58613: result <= 12'b110011101101;
   58614: result <= 12'b110011101101;
   58615: result <= 12'b110011101101;
   58616: result <= 12'b110011101101;
   58617: result <= 12'b110011101101;
   58618: result <= 12'b110011101100;
   58619: result <= 12'b110011101100;
   58620: result <= 12'b110011101100;
   58621: result <= 12'b110011101100;
   58622: result <= 12'b110011101100;
   58623: result <= 12'b110011101100;
   58624: result <= 12'b110011101011;
   58625: result <= 12'b110011101011;
   58626: result <= 12'b110011101011;
   58627: result <= 12'b110011101011;
   58628: result <= 12'b110011101011;
   58629: result <= 12'b110011101011;
   58630: result <= 12'b110011101011;
   58631: result <= 12'b110011101010;
   58632: result <= 12'b110011101010;
   58633: result <= 12'b110011101010;
   58634: result <= 12'b110011101010;
   58635: result <= 12'b110011101010;
   58636: result <= 12'b110011101010;
   58637: result <= 12'b110011101001;
   58638: result <= 12'b110011101001;
   58639: result <= 12'b110011101001;
   58640: result <= 12'b110011101001;
   58641: result <= 12'b110011101001;
   58642: result <= 12'b110011101001;
   58643: result <= 12'b110011101001;
   58644: result <= 12'b110011101000;
   58645: result <= 12'b110011101000;
   58646: result <= 12'b110011101000;
   58647: result <= 12'b110011101000;
   58648: result <= 12'b110011101000;
   58649: result <= 12'b110011101000;
   58650: result <= 12'b110011100111;
   58651: result <= 12'b110011100111;
   58652: result <= 12'b110011100111;
   58653: result <= 12'b110011100111;
   58654: result <= 12'b110011100111;
   58655: result <= 12'b110011100111;
   58656: result <= 12'b110011100111;
   58657: result <= 12'b110011100110;
   58658: result <= 12'b110011100110;
   58659: result <= 12'b110011100110;
   58660: result <= 12'b110011100110;
   58661: result <= 12'b110011100110;
   58662: result <= 12'b110011100110;
   58663: result <= 12'b110011100101;
   58664: result <= 12'b110011100101;
   58665: result <= 12'b110011100101;
   58666: result <= 12'b110011100101;
   58667: result <= 12'b110011100101;
   58668: result <= 12'b110011100101;
   58669: result <= 12'b110011100101;
   58670: result <= 12'b110011100100;
   58671: result <= 12'b110011100100;
   58672: result <= 12'b110011100100;
   58673: result <= 12'b110011100100;
   58674: result <= 12'b110011100100;
   58675: result <= 12'b110011100100;
   58676: result <= 12'b110011100011;
   58677: result <= 12'b110011100011;
   58678: result <= 12'b110011100011;
   58679: result <= 12'b110011100011;
   58680: result <= 12'b110011100011;
   58681: result <= 12'b110011100011;
   58682: result <= 12'b110011100010;
   58683: result <= 12'b110011100010;
   58684: result <= 12'b110011100010;
   58685: result <= 12'b110011100010;
   58686: result <= 12'b110011100010;
   58687: result <= 12'b110011100010;
   58688: result <= 12'b110011100010;
   58689: result <= 12'b110011100001;
   58690: result <= 12'b110011100001;
   58691: result <= 12'b110011100001;
   58692: result <= 12'b110011100001;
   58693: result <= 12'b110011100001;
   58694: result <= 12'b110011100001;
   58695: result <= 12'b110011100000;
   58696: result <= 12'b110011100000;
   58697: result <= 12'b110011100000;
   58698: result <= 12'b110011100000;
   58699: result <= 12'b110011100000;
   58700: result <= 12'b110011100000;
   58701: result <= 12'b110011100000;
   58702: result <= 12'b110011011111;
   58703: result <= 12'b110011011111;
   58704: result <= 12'b110011011111;
   58705: result <= 12'b110011011111;
   58706: result <= 12'b110011011111;
   58707: result <= 12'b110011011111;
   58708: result <= 12'b110011011110;
   58709: result <= 12'b110011011110;
   58710: result <= 12'b110011011110;
   58711: result <= 12'b110011011110;
   58712: result <= 12'b110011011110;
   58713: result <= 12'b110011011110;
   58714: result <= 12'b110011011110;
   58715: result <= 12'b110011011101;
   58716: result <= 12'b110011011101;
   58717: result <= 12'b110011011101;
   58718: result <= 12'b110011011101;
   58719: result <= 12'b110011011101;
   58720: result <= 12'b110011011101;
   58721: result <= 12'b110011011100;
   58722: result <= 12'b110011011100;
   58723: result <= 12'b110011011100;
   58724: result <= 12'b110011011100;
   58725: result <= 12'b110011011100;
   58726: result <= 12'b110011011100;
   58727: result <= 12'b110011011011;
   58728: result <= 12'b110011011011;
   58729: result <= 12'b110011011011;
   58730: result <= 12'b110011011011;
   58731: result <= 12'b110011011011;
   58732: result <= 12'b110011011011;
   58733: result <= 12'b110011011011;
   58734: result <= 12'b110011011010;
   58735: result <= 12'b110011011010;
   58736: result <= 12'b110011011010;
   58737: result <= 12'b110011011010;
   58738: result <= 12'b110011011010;
   58739: result <= 12'b110011011010;
   58740: result <= 12'b110011011001;
   58741: result <= 12'b110011011001;
   58742: result <= 12'b110011011001;
   58743: result <= 12'b110011011001;
   58744: result <= 12'b110011011001;
   58745: result <= 12'b110011011001;
   58746: result <= 12'b110011011001;
   58747: result <= 12'b110011011000;
   58748: result <= 12'b110011011000;
   58749: result <= 12'b110011011000;
   58750: result <= 12'b110011011000;
   58751: result <= 12'b110011011000;
   58752: result <= 12'b110011011000;
   58753: result <= 12'b110011010111;
   58754: result <= 12'b110011010111;
   58755: result <= 12'b110011010111;
   58756: result <= 12'b110011010111;
   58757: result <= 12'b110011010111;
   58758: result <= 12'b110011010111;
   58759: result <= 12'b110011010110;
   58760: result <= 12'b110011010110;
   58761: result <= 12'b110011010110;
   58762: result <= 12'b110011010110;
   58763: result <= 12'b110011010110;
   58764: result <= 12'b110011010110;
   58765: result <= 12'b110011010110;
   58766: result <= 12'b110011010101;
   58767: result <= 12'b110011010101;
   58768: result <= 12'b110011010101;
   58769: result <= 12'b110011010101;
   58770: result <= 12'b110011010101;
   58771: result <= 12'b110011010101;
   58772: result <= 12'b110011010100;
   58773: result <= 12'b110011010100;
   58774: result <= 12'b110011010100;
   58775: result <= 12'b110011010100;
   58776: result <= 12'b110011010100;
   58777: result <= 12'b110011010100;
   58778: result <= 12'b110011010100;
   58779: result <= 12'b110011010011;
   58780: result <= 12'b110011010011;
   58781: result <= 12'b110011010011;
   58782: result <= 12'b110011010011;
   58783: result <= 12'b110011010011;
   58784: result <= 12'b110011010011;
   58785: result <= 12'b110011010010;
   58786: result <= 12'b110011010010;
   58787: result <= 12'b110011010010;
   58788: result <= 12'b110011010010;
   58789: result <= 12'b110011010010;
   58790: result <= 12'b110011010010;
   58791: result <= 12'b110011010001;
   58792: result <= 12'b110011010001;
   58793: result <= 12'b110011010001;
   58794: result <= 12'b110011010001;
   58795: result <= 12'b110011010001;
   58796: result <= 12'b110011010001;
   58797: result <= 12'b110011010001;
   58798: result <= 12'b110011010000;
   58799: result <= 12'b110011010000;
   58800: result <= 12'b110011010000;
   58801: result <= 12'b110011010000;
   58802: result <= 12'b110011010000;
   58803: result <= 12'b110011010000;
   58804: result <= 12'b110011001111;
   58805: result <= 12'b110011001111;
   58806: result <= 12'b110011001111;
   58807: result <= 12'b110011001111;
   58808: result <= 12'b110011001111;
   58809: result <= 12'b110011001111;
   58810: result <= 12'b110011001111;
   58811: result <= 12'b110011001110;
   58812: result <= 12'b110011001110;
   58813: result <= 12'b110011001110;
   58814: result <= 12'b110011001110;
   58815: result <= 12'b110011001110;
   58816: result <= 12'b110011001110;
   58817: result <= 12'b110011001101;
   58818: result <= 12'b110011001101;
   58819: result <= 12'b110011001101;
   58820: result <= 12'b110011001101;
   58821: result <= 12'b110011001101;
   58822: result <= 12'b110011001101;
   58823: result <= 12'b110011001100;
   58824: result <= 12'b110011001100;
   58825: result <= 12'b110011001100;
   58826: result <= 12'b110011001100;
   58827: result <= 12'b110011001100;
   58828: result <= 12'b110011001100;
   58829: result <= 12'b110011001100;
   58830: result <= 12'b110011001011;
   58831: result <= 12'b110011001011;
   58832: result <= 12'b110011001011;
   58833: result <= 12'b110011001011;
   58834: result <= 12'b110011001011;
   58835: result <= 12'b110011001011;
   58836: result <= 12'b110011001010;
   58837: result <= 12'b110011001010;
   58838: result <= 12'b110011001010;
   58839: result <= 12'b110011001010;
   58840: result <= 12'b110011001010;
   58841: result <= 12'b110011001010;
   58842: result <= 12'b110011001001;
   58843: result <= 12'b110011001001;
   58844: result <= 12'b110011001001;
   58845: result <= 12'b110011001001;
   58846: result <= 12'b110011001001;
   58847: result <= 12'b110011001001;
   58848: result <= 12'b110011001001;
   58849: result <= 12'b110011001000;
   58850: result <= 12'b110011001000;
   58851: result <= 12'b110011001000;
   58852: result <= 12'b110011001000;
   58853: result <= 12'b110011001000;
   58854: result <= 12'b110011001000;
   58855: result <= 12'b110011000111;
   58856: result <= 12'b110011000111;
   58857: result <= 12'b110011000111;
   58858: result <= 12'b110011000111;
   58859: result <= 12'b110011000111;
   58860: result <= 12'b110011000111;
   58861: result <= 12'b110011000110;
   58862: result <= 12'b110011000110;
   58863: result <= 12'b110011000110;
   58864: result <= 12'b110011000110;
   58865: result <= 12'b110011000110;
   58866: result <= 12'b110011000110;
   58867: result <= 12'b110011000110;
   58868: result <= 12'b110011000101;
   58869: result <= 12'b110011000101;
   58870: result <= 12'b110011000101;
   58871: result <= 12'b110011000101;
   58872: result <= 12'b110011000101;
   58873: result <= 12'b110011000101;
   58874: result <= 12'b110011000100;
   58875: result <= 12'b110011000100;
   58876: result <= 12'b110011000100;
   58877: result <= 12'b110011000100;
   58878: result <= 12'b110011000100;
   58879: result <= 12'b110011000100;
   58880: result <= 12'b110011000011;
   58881: result <= 12'b110011000011;
   58882: result <= 12'b110011000011;
   58883: result <= 12'b110011000011;
   58884: result <= 12'b110011000011;
   58885: result <= 12'b110011000011;
   58886: result <= 12'b110011000011;
   58887: result <= 12'b110011000010;
   58888: result <= 12'b110011000010;
   58889: result <= 12'b110011000010;
   58890: result <= 12'b110011000010;
   58891: result <= 12'b110011000010;
   58892: result <= 12'b110011000010;
   58893: result <= 12'b110011000001;
   58894: result <= 12'b110011000001;
   58895: result <= 12'b110011000001;
   58896: result <= 12'b110011000001;
   58897: result <= 12'b110011000001;
   58898: result <= 12'b110011000001;
   58899: result <= 12'b110011000000;
   58900: result <= 12'b110011000000;
   58901: result <= 12'b110011000000;
   58902: result <= 12'b110011000000;
   58903: result <= 12'b110011000000;
   58904: result <= 12'b110011000000;
   58905: result <= 12'b110011000000;
   58906: result <= 12'b110010111111;
   58907: result <= 12'b110010111111;
   58908: result <= 12'b110010111111;
   58909: result <= 12'b110010111111;
   58910: result <= 12'b110010111111;
   58911: result <= 12'b110010111111;
   58912: result <= 12'b110010111110;
   58913: result <= 12'b110010111110;
   58914: result <= 12'b110010111110;
   58915: result <= 12'b110010111110;
   58916: result <= 12'b110010111110;
   58917: result <= 12'b110010111110;
   58918: result <= 12'b110010111101;
   58919: result <= 12'b110010111101;
   58920: result <= 12'b110010111101;
   58921: result <= 12'b110010111101;
   58922: result <= 12'b110010111101;
   58923: result <= 12'b110010111101;
   58924: result <= 12'b110010111101;
   58925: result <= 12'b110010111100;
   58926: result <= 12'b110010111100;
   58927: result <= 12'b110010111100;
   58928: result <= 12'b110010111100;
   58929: result <= 12'b110010111100;
   58930: result <= 12'b110010111100;
   58931: result <= 12'b110010111011;
   58932: result <= 12'b110010111011;
   58933: result <= 12'b110010111011;
   58934: result <= 12'b110010111011;
   58935: result <= 12'b110010111011;
   58936: result <= 12'b110010111011;
   58937: result <= 12'b110010111010;
   58938: result <= 12'b110010111010;
   58939: result <= 12'b110010111010;
   58940: result <= 12'b110010111010;
   58941: result <= 12'b110010111010;
   58942: result <= 12'b110010111010;
   58943: result <= 12'b110010111010;
   58944: result <= 12'b110010111001;
   58945: result <= 12'b110010111001;
   58946: result <= 12'b110010111001;
   58947: result <= 12'b110010111001;
   58948: result <= 12'b110010111001;
   58949: result <= 12'b110010111001;
   58950: result <= 12'b110010111000;
   58951: result <= 12'b110010111000;
   58952: result <= 12'b110010111000;
   58953: result <= 12'b110010111000;
   58954: result <= 12'b110010111000;
   58955: result <= 12'b110010111000;
   58956: result <= 12'b110010110111;
   58957: result <= 12'b110010110111;
   58958: result <= 12'b110010110111;
   58959: result <= 12'b110010110111;
   58960: result <= 12'b110010110111;
   58961: result <= 12'b110010110111;
   58962: result <= 12'b110010110111;
   58963: result <= 12'b110010110110;
   58964: result <= 12'b110010110110;
   58965: result <= 12'b110010110110;
   58966: result <= 12'b110010110110;
   58967: result <= 12'b110010110110;
   58968: result <= 12'b110010110110;
   58969: result <= 12'b110010110101;
   58970: result <= 12'b110010110101;
   58971: result <= 12'b110010110101;
   58972: result <= 12'b110010110101;
   58973: result <= 12'b110010110101;
   58974: result <= 12'b110010110101;
   58975: result <= 12'b110010110100;
   58976: result <= 12'b110010110100;
   58977: result <= 12'b110010110100;
   58978: result <= 12'b110010110100;
   58979: result <= 12'b110010110100;
   58980: result <= 12'b110010110100;
   58981: result <= 12'b110010110100;
   58982: result <= 12'b110010110011;
   58983: result <= 12'b110010110011;
   58984: result <= 12'b110010110011;
   58985: result <= 12'b110010110011;
   58986: result <= 12'b110010110011;
   58987: result <= 12'b110010110011;
   58988: result <= 12'b110010110010;
   58989: result <= 12'b110010110010;
   58990: result <= 12'b110010110010;
   58991: result <= 12'b110010110010;
   58992: result <= 12'b110010110010;
   58993: result <= 12'b110010110010;
   58994: result <= 12'b110010110001;
   58995: result <= 12'b110010110001;
   58996: result <= 12'b110010110001;
   58997: result <= 12'b110010110001;
   58998: result <= 12'b110010110001;
   58999: result <= 12'b110010110001;
   59000: result <= 12'b110010110000;
   59001: result <= 12'b110010110000;
   59002: result <= 12'b110010110000;
   59003: result <= 12'b110010110000;
   59004: result <= 12'b110010110000;
   59005: result <= 12'b110010110000;
   59006: result <= 12'b110010110000;
   59007: result <= 12'b110010101111;
   59008: result <= 12'b110010101111;
   59009: result <= 12'b110010101111;
   59010: result <= 12'b110010101111;
   59011: result <= 12'b110010101111;
   59012: result <= 12'b110010101111;
   59013: result <= 12'b110010101110;
   59014: result <= 12'b110010101110;
   59015: result <= 12'b110010101110;
   59016: result <= 12'b110010101110;
   59017: result <= 12'b110010101110;
   59018: result <= 12'b110010101110;
   59019: result <= 12'b110010101101;
   59020: result <= 12'b110010101101;
   59021: result <= 12'b110010101101;
   59022: result <= 12'b110010101101;
   59023: result <= 12'b110010101101;
   59024: result <= 12'b110010101101;
   59025: result <= 12'b110010101101;
   59026: result <= 12'b110010101100;
   59027: result <= 12'b110010101100;
   59028: result <= 12'b110010101100;
   59029: result <= 12'b110010101100;
   59030: result <= 12'b110010101100;
   59031: result <= 12'b110010101100;
   59032: result <= 12'b110010101011;
   59033: result <= 12'b110010101011;
   59034: result <= 12'b110010101011;
   59035: result <= 12'b110010101011;
   59036: result <= 12'b110010101011;
   59037: result <= 12'b110010101011;
   59038: result <= 12'b110010101010;
   59039: result <= 12'b110010101010;
   59040: result <= 12'b110010101010;
   59041: result <= 12'b110010101010;
   59042: result <= 12'b110010101010;
   59043: result <= 12'b110010101010;
   59044: result <= 12'b110010101001;
   59045: result <= 12'b110010101001;
   59046: result <= 12'b110010101001;
   59047: result <= 12'b110010101001;
   59048: result <= 12'b110010101001;
   59049: result <= 12'b110010101001;
   59050: result <= 12'b110010101001;
   59051: result <= 12'b110010101000;
   59052: result <= 12'b110010101000;
   59053: result <= 12'b110010101000;
   59054: result <= 12'b110010101000;
   59055: result <= 12'b110010101000;
   59056: result <= 12'b110010101000;
   59057: result <= 12'b110010100111;
   59058: result <= 12'b110010100111;
   59059: result <= 12'b110010100111;
   59060: result <= 12'b110010100111;
   59061: result <= 12'b110010100111;
   59062: result <= 12'b110010100111;
   59063: result <= 12'b110010100110;
   59064: result <= 12'b110010100110;
   59065: result <= 12'b110010100110;
   59066: result <= 12'b110010100110;
   59067: result <= 12'b110010100110;
   59068: result <= 12'b110010100110;
   59069: result <= 12'b110010100101;
   59070: result <= 12'b110010100101;
   59071: result <= 12'b110010100101;
   59072: result <= 12'b110010100101;
   59073: result <= 12'b110010100101;
   59074: result <= 12'b110010100101;
   59075: result <= 12'b110010100101;
   59076: result <= 12'b110010100100;
   59077: result <= 12'b110010100100;
   59078: result <= 12'b110010100100;
   59079: result <= 12'b110010100100;
   59080: result <= 12'b110010100100;
   59081: result <= 12'b110010100100;
   59082: result <= 12'b110010100011;
   59083: result <= 12'b110010100011;
   59084: result <= 12'b110010100011;
   59085: result <= 12'b110010100011;
   59086: result <= 12'b110010100011;
   59087: result <= 12'b110010100011;
   59088: result <= 12'b110010100010;
   59089: result <= 12'b110010100010;
   59090: result <= 12'b110010100010;
   59091: result <= 12'b110010100010;
   59092: result <= 12'b110010100010;
   59093: result <= 12'b110010100010;
   59094: result <= 12'b110010100001;
   59095: result <= 12'b110010100001;
   59096: result <= 12'b110010100001;
   59097: result <= 12'b110010100001;
   59098: result <= 12'b110010100001;
   59099: result <= 12'b110010100001;
   59100: result <= 12'b110010100001;
   59101: result <= 12'b110010100000;
   59102: result <= 12'b110010100000;
   59103: result <= 12'b110010100000;
   59104: result <= 12'b110010100000;
   59105: result <= 12'b110010100000;
   59106: result <= 12'b110010100000;
   59107: result <= 12'b110010011111;
   59108: result <= 12'b110010011111;
   59109: result <= 12'b110010011111;
   59110: result <= 12'b110010011111;
   59111: result <= 12'b110010011111;
   59112: result <= 12'b110010011111;
   59113: result <= 12'b110010011110;
   59114: result <= 12'b110010011110;
   59115: result <= 12'b110010011110;
   59116: result <= 12'b110010011110;
   59117: result <= 12'b110010011110;
   59118: result <= 12'b110010011110;
   59119: result <= 12'b110010011101;
   59120: result <= 12'b110010011101;
   59121: result <= 12'b110010011101;
   59122: result <= 12'b110010011101;
   59123: result <= 12'b110010011101;
   59124: result <= 12'b110010011101;
   59125: result <= 12'b110010011101;
   59126: result <= 12'b110010011100;
   59127: result <= 12'b110010011100;
   59128: result <= 12'b110010011100;
   59129: result <= 12'b110010011100;
   59130: result <= 12'b110010011100;
   59131: result <= 12'b110010011100;
   59132: result <= 12'b110010011011;
   59133: result <= 12'b110010011011;
   59134: result <= 12'b110010011011;
   59135: result <= 12'b110010011011;
   59136: result <= 12'b110010011011;
   59137: result <= 12'b110010011011;
   59138: result <= 12'b110010011010;
   59139: result <= 12'b110010011010;
   59140: result <= 12'b110010011010;
   59141: result <= 12'b110010011010;
   59142: result <= 12'b110010011010;
   59143: result <= 12'b110010011010;
   59144: result <= 12'b110010011001;
   59145: result <= 12'b110010011001;
   59146: result <= 12'b110010011001;
   59147: result <= 12'b110010011001;
   59148: result <= 12'b110010011001;
   59149: result <= 12'b110010011001;
   59150: result <= 12'b110010011001;
   59151: result <= 12'b110010011000;
   59152: result <= 12'b110010011000;
   59153: result <= 12'b110010011000;
   59154: result <= 12'b110010011000;
   59155: result <= 12'b110010011000;
   59156: result <= 12'b110010011000;
   59157: result <= 12'b110010010111;
   59158: result <= 12'b110010010111;
   59159: result <= 12'b110010010111;
   59160: result <= 12'b110010010111;
   59161: result <= 12'b110010010111;
   59162: result <= 12'b110010010111;
   59163: result <= 12'b110010010110;
   59164: result <= 12'b110010010110;
   59165: result <= 12'b110010010110;
   59166: result <= 12'b110010010110;
   59167: result <= 12'b110010010110;
   59168: result <= 12'b110010010110;
   59169: result <= 12'b110010010101;
   59170: result <= 12'b110010010101;
   59171: result <= 12'b110010010101;
   59172: result <= 12'b110010010101;
   59173: result <= 12'b110010010101;
   59174: result <= 12'b110010010101;
   59175: result <= 12'b110010010100;
   59176: result <= 12'b110010010100;
   59177: result <= 12'b110010010100;
   59178: result <= 12'b110010010100;
   59179: result <= 12'b110010010100;
   59180: result <= 12'b110010010100;
   59181: result <= 12'b110010010100;
   59182: result <= 12'b110010010011;
   59183: result <= 12'b110010010011;
   59184: result <= 12'b110010010011;
   59185: result <= 12'b110010010011;
   59186: result <= 12'b110010010011;
   59187: result <= 12'b110010010011;
   59188: result <= 12'b110010010010;
   59189: result <= 12'b110010010010;
   59190: result <= 12'b110010010010;
   59191: result <= 12'b110010010010;
   59192: result <= 12'b110010010010;
   59193: result <= 12'b110010010010;
   59194: result <= 12'b110010010001;
   59195: result <= 12'b110010010001;
   59196: result <= 12'b110010010001;
   59197: result <= 12'b110010010001;
   59198: result <= 12'b110010010001;
   59199: result <= 12'b110010010001;
   59200: result <= 12'b110010010000;
   59201: result <= 12'b110010010000;
   59202: result <= 12'b110010010000;
   59203: result <= 12'b110010010000;
   59204: result <= 12'b110010010000;
   59205: result <= 12'b110010010000;
   59206: result <= 12'b110010001111;
   59207: result <= 12'b110010001111;
   59208: result <= 12'b110010001111;
   59209: result <= 12'b110010001111;
   59210: result <= 12'b110010001111;
   59211: result <= 12'b110010001111;
   59212: result <= 12'b110010001111;
   59213: result <= 12'b110010001110;
   59214: result <= 12'b110010001110;
   59215: result <= 12'b110010001110;
   59216: result <= 12'b110010001110;
   59217: result <= 12'b110010001110;
   59218: result <= 12'b110010001110;
   59219: result <= 12'b110010001101;
   59220: result <= 12'b110010001101;
   59221: result <= 12'b110010001101;
   59222: result <= 12'b110010001101;
   59223: result <= 12'b110010001101;
   59224: result <= 12'b110010001101;
   59225: result <= 12'b110010001100;
   59226: result <= 12'b110010001100;
   59227: result <= 12'b110010001100;
   59228: result <= 12'b110010001100;
   59229: result <= 12'b110010001100;
   59230: result <= 12'b110010001100;
   59231: result <= 12'b110010001011;
   59232: result <= 12'b110010001011;
   59233: result <= 12'b110010001011;
   59234: result <= 12'b110010001011;
   59235: result <= 12'b110010001011;
   59236: result <= 12'b110010001011;
   59237: result <= 12'b110010001010;
   59238: result <= 12'b110010001010;
   59239: result <= 12'b110010001010;
   59240: result <= 12'b110010001010;
   59241: result <= 12'b110010001010;
   59242: result <= 12'b110010001010;
   59243: result <= 12'b110010001010;
   59244: result <= 12'b110010001001;
   59245: result <= 12'b110010001001;
   59246: result <= 12'b110010001001;
   59247: result <= 12'b110010001001;
   59248: result <= 12'b110010001001;
   59249: result <= 12'b110010001001;
   59250: result <= 12'b110010001000;
   59251: result <= 12'b110010001000;
   59252: result <= 12'b110010001000;
   59253: result <= 12'b110010001000;
   59254: result <= 12'b110010001000;
   59255: result <= 12'b110010001000;
   59256: result <= 12'b110010000111;
   59257: result <= 12'b110010000111;
   59258: result <= 12'b110010000111;
   59259: result <= 12'b110010000111;
   59260: result <= 12'b110010000111;
   59261: result <= 12'b110010000111;
   59262: result <= 12'b110010000110;
   59263: result <= 12'b110010000110;
   59264: result <= 12'b110010000110;
   59265: result <= 12'b110010000110;
   59266: result <= 12'b110010000110;
   59267: result <= 12'b110010000110;
   59268: result <= 12'b110010000101;
   59269: result <= 12'b110010000101;
   59270: result <= 12'b110010000101;
   59271: result <= 12'b110010000101;
   59272: result <= 12'b110010000101;
   59273: result <= 12'b110010000101;
   59274: result <= 12'b110010000100;
   59275: result <= 12'b110010000100;
   59276: result <= 12'b110010000100;
   59277: result <= 12'b110010000100;
   59278: result <= 12'b110010000100;
   59279: result <= 12'b110010000100;
   59280: result <= 12'b110010000100;
   59281: result <= 12'b110010000011;
   59282: result <= 12'b110010000011;
   59283: result <= 12'b110010000011;
   59284: result <= 12'b110010000011;
   59285: result <= 12'b110010000011;
   59286: result <= 12'b110010000011;
   59287: result <= 12'b110010000010;
   59288: result <= 12'b110010000010;
   59289: result <= 12'b110010000010;
   59290: result <= 12'b110010000010;
   59291: result <= 12'b110010000010;
   59292: result <= 12'b110010000010;
   59293: result <= 12'b110010000001;
   59294: result <= 12'b110010000001;
   59295: result <= 12'b110010000001;
   59296: result <= 12'b110010000001;
   59297: result <= 12'b110010000001;
   59298: result <= 12'b110010000001;
   59299: result <= 12'b110010000000;
   59300: result <= 12'b110010000000;
   59301: result <= 12'b110010000000;
   59302: result <= 12'b110010000000;
   59303: result <= 12'b110010000000;
   59304: result <= 12'b110010000000;
   59305: result <= 12'b110001111111;
   59306: result <= 12'b110001111111;
   59307: result <= 12'b110001111111;
   59308: result <= 12'b110001111111;
   59309: result <= 12'b110001111111;
   59310: result <= 12'b110001111111;
   59311: result <= 12'b110001111110;
   59312: result <= 12'b110001111110;
   59313: result <= 12'b110001111110;
   59314: result <= 12'b110001111110;
   59315: result <= 12'b110001111110;
   59316: result <= 12'b110001111110;
   59317: result <= 12'b110001111110;
   59318: result <= 12'b110001111101;
   59319: result <= 12'b110001111101;
   59320: result <= 12'b110001111101;
   59321: result <= 12'b110001111101;
   59322: result <= 12'b110001111101;
   59323: result <= 12'b110001111101;
   59324: result <= 12'b110001111100;
   59325: result <= 12'b110001111100;
   59326: result <= 12'b110001111100;
   59327: result <= 12'b110001111100;
   59328: result <= 12'b110001111100;
   59329: result <= 12'b110001111100;
   59330: result <= 12'b110001111011;
   59331: result <= 12'b110001111011;
   59332: result <= 12'b110001111011;
   59333: result <= 12'b110001111011;
   59334: result <= 12'b110001111011;
   59335: result <= 12'b110001111011;
   59336: result <= 12'b110001111010;
   59337: result <= 12'b110001111010;
   59338: result <= 12'b110001111010;
   59339: result <= 12'b110001111010;
   59340: result <= 12'b110001111010;
   59341: result <= 12'b110001111010;
   59342: result <= 12'b110001111001;
   59343: result <= 12'b110001111001;
   59344: result <= 12'b110001111001;
   59345: result <= 12'b110001111001;
   59346: result <= 12'b110001111001;
   59347: result <= 12'b110001111001;
   59348: result <= 12'b110001111000;
   59349: result <= 12'b110001111000;
   59350: result <= 12'b110001111000;
   59351: result <= 12'b110001111000;
   59352: result <= 12'b110001111000;
   59353: result <= 12'b110001111000;
   59354: result <= 12'b110001111000;
   59355: result <= 12'b110001110111;
   59356: result <= 12'b110001110111;
   59357: result <= 12'b110001110111;
   59358: result <= 12'b110001110111;
   59359: result <= 12'b110001110111;
   59360: result <= 12'b110001110111;
   59361: result <= 12'b110001110110;
   59362: result <= 12'b110001110110;
   59363: result <= 12'b110001110110;
   59364: result <= 12'b110001110110;
   59365: result <= 12'b110001110110;
   59366: result <= 12'b110001110110;
   59367: result <= 12'b110001110101;
   59368: result <= 12'b110001110101;
   59369: result <= 12'b110001110101;
   59370: result <= 12'b110001110101;
   59371: result <= 12'b110001110101;
   59372: result <= 12'b110001110101;
   59373: result <= 12'b110001110100;
   59374: result <= 12'b110001110100;
   59375: result <= 12'b110001110100;
   59376: result <= 12'b110001110100;
   59377: result <= 12'b110001110100;
   59378: result <= 12'b110001110100;
   59379: result <= 12'b110001110011;
   59380: result <= 12'b110001110011;
   59381: result <= 12'b110001110011;
   59382: result <= 12'b110001110011;
   59383: result <= 12'b110001110011;
   59384: result <= 12'b110001110011;
   59385: result <= 12'b110001110010;
   59386: result <= 12'b110001110010;
   59387: result <= 12'b110001110010;
   59388: result <= 12'b110001110010;
   59389: result <= 12'b110001110010;
   59390: result <= 12'b110001110010;
   59391: result <= 12'b110001110001;
   59392: result <= 12'b110001110001;
   59393: result <= 12'b110001110001;
   59394: result <= 12'b110001110001;
   59395: result <= 12'b110001110001;
   59396: result <= 12'b110001110001;
   59397: result <= 12'b110001110000;
   59398: result <= 12'b110001110000;
   59399: result <= 12'b110001110000;
   59400: result <= 12'b110001110000;
   59401: result <= 12'b110001110000;
   59402: result <= 12'b110001110000;
   59403: result <= 12'b110001110000;
   59404: result <= 12'b110001101111;
   59405: result <= 12'b110001101111;
   59406: result <= 12'b110001101111;
   59407: result <= 12'b110001101111;
   59408: result <= 12'b110001101111;
   59409: result <= 12'b110001101111;
   59410: result <= 12'b110001101110;
   59411: result <= 12'b110001101110;
   59412: result <= 12'b110001101110;
   59413: result <= 12'b110001101110;
   59414: result <= 12'b110001101110;
   59415: result <= 12'b110001101110;
   59416: result <= 12'b110001101101;
   59417: result <= 12'b110001101101;
   59418: result <= 12'b110001101101;
   59419: result <= 12'b110001101101;
   59420: result <= 12'b110001101101;
   59421: result <= 12'b110001101101;
   59422: result <= 12'b110001101100;
   59423: result <= 12'b110001101100;
   59424: result <= 12'b110001101100;
   59425: result <= 12'b110001101100;
   59426: result <= 12'b110001101100;
   59427: result <= 12'b110001101100;
   59428: result <= 12'b110001101011;
   59429: result <= 12'b110001101011;
   59430: result <= 12'b110001101011;
   59431: result <= 12'b110001101011;
   59432: result <= 12'b110001101011;
   59433: result <= 12'b110001101011;
   59434: result <= 12'b110001101010;
   59435: result <= 12'b110001101010;
   59436: result <= 12'b110001101010;
   59437: result <= 12'b110001101010;
   59438: result <= 12'b110001101010;
   59439: result <= 12'b110001101010;
   59440: result <= 12'b110001101001;
   59441: result <= 12'b110001101001;
   59442: result <= 12'b110001101001;
   59443: result <= 12'b110001101001;
   59444: result <= 12'b110001101001;
   59445: result <= 12'b110001101001;
   59446: result <= 12'b110001101000;
   59447: result <= 12'b110001101000;
   59448: result <= 12'b110001101000;
   59449: result <= 12'b110001101000;
   59450: result <= 12'b110001101000;
   59451: result <= 12'b110001101000;
   59452: result <= 12'b110001100111;
   59453: result <= 12'b110001100111;
   59454: result <= 12'b110001100111;
   59455: result <= 12'b110001100111;
   59456: result <= 12'b110001100111;
   59457: result <= 12'b110001100111;
   59458: result <= 12'b110001100111;
   59459: result <= 12'b110001100110;
   59460: result <= 12'b110001100110;
   59461: result <= 12'b110001100110;
   59462: result <= 12'b110001100110;
   59463: result <= 12'b110001100110;
   59464: result <= 12'b110001100110;
   59465: result <= 12'b110001100101;
   59466: result <= 12'b110001100101;
   59467: result <= 12'b110001100101;
   59468: result <= 12'b110001100101;
   59469: result <= 12'b110001100101;
   59470: result <= 12'b110001100101;
   59471: result <= 12'b110001100100;
   59472: result <= 12'b110001100100;
   59473: result <= 12'b110001100100;
   59474: result <= 12'b110001100100;
   59475: result <= 12'b110001100100;
   59476: result <= 12'b110001100100;
   59477: result <= 12'b110001100011;
   59478: result <= 12'b110001100011;
   59479: result <= 12'b110001100011;
   59480: result <= 12'b110001100011;
   59481: result <= 12'b110001100011;
   59482: result <= 12'b110001100011;
   59483: result <= 12'b110001100010;
   59484: result <= 12'b110001100010;
   59485: result <= 12'b110001100010;
   59486: result <= 12'b110001100010;
   59487: result <= 12'b110001100010;
   59488: result <= 12'b110001100010;
   59489: result <= 12'b110001100001;
   59490: result <= 12'b110001100001;
   59491: result <= 12'b110001100001;
   59492: result <= 12'b110001100001;
   59493: result <= 12'b110001100001;
   59494: result <= 12'b110001100001;
   59495: result <= 12'b110001100000;
   59496: result <= 12'b110001100000;
   59497: result <= 12'b110001100000;
   59498: result <= 12'b110001100000;
   59499: result <= 12'b110001100000;
   59500: result <= 12'b110001100000;
   59501: result <= 12'b110001011111;
   59502: result <= 12'b110001011111;
   59503: result <= 12'b110001011111;
   59504: result <= 12'b110001011111;
   59505: result <= 12'b110001011111;
   59506: result <= 12'b110001011111;
   59507: result <= 12'b110001011110;
   59508: result <= 12'b110001011110;
   59509: result <= 12'b110001011110;
   59510: result <= 12'b110001011110;
   59511: result <= 12'b110001011110;
   59512: result <= 12'b110001011110;
   59513: result <= 12'b110001011101;
   59514: result <= 12'b110001011101;
   59515: result <= 12'b110001011101;
   59516: result <= 12'b110001011101;
   59517: result <= 12'b110001011101;
   59518: result <= 12'b110001011101;
   59519: result <= 12'b110001011100;
   59520: result <= 12'b110001011100;
   59521: result <= 12'b110001011100;
   59522: result <= 12'b110001011100;
   59523: result <= 12'b110001011100;
   59524: result <= 12'b110001011100;
   59525: result <= 12'b110001011100;
   59526: result <= 12'b110001011011;
   59527: result <= 12'b110001011011;
   59528: result <= 12'b110001011011;
   59529: result <= 12'b110001011011;
   59530: result <= 12'b110001011011;
   59531: result <= 12'b110001011011;
   59532: result <= 12'b110001011010;
   59533: result <= 12'b110001011010;
   59534: result <= 12'b110001011010;
   59535: result <= 12'b110001011010;
   59536: result <= 12'b110001011010;
   59537: result <= 12'b110001011010;
   59538: result <= 12'b110001011001;
   59539: result <= 12'b110001011001;
   59540: result <= 12'b110001011001;
   59541: result <= 12'b110001011001;
   59542: result <= 12'b110001011001;
   59543: result <= 12'b110001011001;
   59544: result <= 12'b110001011000;
   59545: result <= 12'b110001011000;
   59546: result <= 12'b110001011000;
   59547: result <= 12'b110001011000;
   59548: result <= 12'b110001011000;
   59549: result <= 12'b110001011000;
   59550: result <= 12'b110001010111;
   59551: result <= 12'b110001010111;
   59552: result <= 12'b110001010111;
   59553: result <= 12'b110001010111;
   59554: result <= 12'b110001010111;
   59555: result <= 12'b110001010111;
   59556: result <= 12'b110001010110;
   59557: result <= 12'b110001010110;
   59558: result <= 12'b110001010110;
   59559: result <= 12'b110001010110;
   59560: result <= 12'b110001010110;
   59561: result <= 12'b110001010110;
   59562: result <= 12'b110001010101;
   59563: result <= 12'b110001010101;
   59564: result <= 12'b110001010101;
   59565: result <= 12'b110001010101;
   59566: result <= 12'b110001010101;
   59567: result <= 12'b110001010101;
   59568: result <= 12'b110001010100;
   59569: result <= 12'b110001010100;
   59570: result <= 12'b110001010100;
   59571: result <= 12'b110001010100;
   59572: result <= 12'b110001010100;
   59573: result <= 12'b110001010100;
   59574: result <= 12'b110001010011;
   59575: result <= 12'b110001010011;
   59576: result <= 12'b110001010011;
   59577: result <= 12'b110001010011;
   59578: result <= 12'b110001010011;
   59579: result <= 12'b110001010011;
   59580: result <= 12'b110001010010;
   59581: result <= 12'b110001010010;
   59582: result <= 12'b110001010010;
   59583: result <= 12'b110001010010;
   59584: result <= 12'b110001010010;
   59585: result <= 12'b110001010010;
   59586: result <= 12'b110001010001;
   59587: result <= 12'b110001010001;
   59588: result <= 12'b110001010001;
   59589: result <= 12'b110001010001;
   59590: result <= 12'b110001010001;
   59591: result <= 12'b110001010001;
   59592: result <= 12'b110001010000;
   59593: result <= 12'b110001010000;
   59594: result <= 12'b110001010000;
   59595: result <= 12'b110001010000;
   59596: result <= 12'b110001010000;
   59597: result <= 12'b110001010000;
   59598: result <= 12'b110001001111;
   59599: result <= 12'b110001001111;
   59600: result <= 12'b110001001111;
   59601: result <= 12'b110001001111;
   59602: result <= 12'b110001001111;
   59603: result <= 12'b110001001111;
   59604: result <= 12'b110001001110;
   59605: result <= 12'b110001001110;
   59606: result <= 12'b110001001110;
   59607: result <= 12'b110001001110;
   59608: result <= 12'b110001001110;
   59609: result <= 12'b110001001110;
   59610: result <= 12'b110001001101;
   59611: result <= 12'b110001001101;
   59612: result <= 12'b110001001101;
   59613: result <= 12'b110001001101;
   59614: result <= 12'b110001001101;
   59615: result <= 12'b110001001101;
   59616: result <= 12'b110001001100;
   59617: result <= 12'b110001001100;
   59618: result <= 12'b110001001100;
   59619: result <= 12'b110001001100;
   59620: result <= 12'b110001001100;
   59621: result <= 12'b110001001100;
   59622: result <= 12'b110001001011;
   59623: result <= 12'b110001001011;
   59624: result <= 12'b110001001011;
   59625: result <= 12'b110001001011;
   59626: result <= 12'b110001001011;
   59627: result <= 12'b110001001011;
   59628: result <= 12'b110001001010;
   59629: result <= 12'b110001001010;
   59630: result <= 12'b110001001010;
   59631: result <= 12'b110001001010;
   59632: result <= 12'b110001001010;
   59633: result <= 12'b110001001010;
   59634: result <= 12'b110001001001;
   59635: result <= 12'b110001001001;
   59636: result <= 12'b110001001001;
   59637: result <= 12'b110001001001;
   59638: result <= 12'b110001001001;
   59639: result <= 12'b110001001001;
   59640: result <= 12'b110001001001;
   59641: result <= 12'b110001001000;
   59642: result <= 12'b110001001000;
   59643: result <= 12'b110001001000;
   59644: result <= 12'b110001001000;
   59645: result <= 12'b110001001000;
   59646: result <= 12'b110001001000;
   59647: result <= 12'b110001000111;
   59648: result <= 12'b110001000111;
   59649: result <= 12'b110001000111;
   59650: result <= 12'b110001000111;
   59651: result <= 12'b110001000111;
   59652: result <= 12'b110001000111;
   59653: result <= 12'b110001000110;
   59654: result <= 12'b110001000110;
   59655: result <= 12'b110001000110;
   59656: result <= 12'b110001000110;
   59657: result <= 12'b110001000110;
   59658: result <= 12'b110001000110;
   59659: result <= 12'b110001000101;
   59660: result <= 12'b110001000101;
   59661: result <= 12'b110001000101;
   59662: result <= 12'b110001000101;
   59663: result <= 12'b110001000101;
   59664: result <= 12'b110001000101;
   59665: result <= 12'b110001000100;
   59666: result <= 12'b110001000100;
   59667: result <= 12'b110001000100;
   59668: result <= 12'b110001000100;
   59669: result <= 12'b110001000100;
   59670: result <= 12'b110001000100;
   59671: result <= 12'b110001000011;
   59672: result <= 12'b110001000011;
   59673: result <= 12'b110001000011;
   59674: result <= 12'b110001000011;
   59675: result <= 12'b110001000011;
   59676: result <= 12'b110001000011;
   59677: result <= 12'b110001000010;
   59678: result <= 12'b110001000010;
   59679: result <= 12'b110001000010;
   59680: result <= 12'b110001000010;
   59681: result <= 12'b110001000010;
   59682: result <= 12'b110001000010;
   59683: result <= 12'b110001000001;
   59684: result <= 12'b110001000001;
   59685: result <= 12'b110001000001;
   59686: result <= 12'b110001000001;
   59687: result <= 12'b110001000001;
   59688: result <= 12'b110001000001;
   59689: result <= 12'b110001000000;
   59690: result <= 12'b110001000000;
   59691: result <= 12'b110001000000;
   59692: result <= 12'b110001000000;
   59693: result <= 12'b110001000000;
   59694: result <= 12'b110001000000;
   59695: result <= 12'b110000111111;
   59696: result <= 12'b110000111111;
   59697: result <= 12'b110000111111;
   59698: result <= 12'b110000111111;
   59699: result <= 12'b110000111111;
   59700: result <= 12'b110000111111;
   59701: result <= 12'b110000111110;
   59702: result <= 12'b110000111110;
   59703: result <= 12'b110000111110;
   59704: result <= 12'b110000111110;
   59705: result <= 12'b110000111110;
   59706: result <= 12'b110000111110;
   59707: result <= 12'b110000111101;
   59708: result <= 12'b110000111101;
   59709: result <= 12'b110000111101;
   59710: result <= 12'b110000111101;
   59711: result <= 12'b110000111101;
   59712: result <= 12'b110000111101;
   59713: result <= 12'b110000111100;
   59714: result <= 12'b110000111100;
   59715: result <= 12'b110000111100;
   59716: result <= 12'b110000111100;
   59717: result <= 12'b110000111100;
   59718: result <= 12'b110000111100;
   59719: result <= 12'b110000111011;
   59720: result <= 12'b110000111011;
   59721: result <= 12'b110000111011;
   59722: result <= 12'b110000111011;
   59723: result <= 12'b110000111011;
   59724: result <= 12'b110000111011;
   59725: result <= 12'b110000111010;
   59726: result <= 12'b110000111010;
   59727: result <= 12'b110000111010;
   59728: result <= 12'b110000111010;
   59729: result <= 12'b110000111010;
   59730: result <= 12'b110000111010;
   59731: result <= 12'b110000111001;
   59732: result <= 12'b110000111001;
   59733: result <= 12'b110000111001;
   59734: result <= 12'b110000111001;
   59735: result <= 12'b110000111001;
   59736: result <= 12'b110000111001;
   59737: result <= 12'b110000111000;
   59738: result <= 12'b110000111000;
   59739: result <= 12'b110000111000;
   59740: result <= 12'b110000111000;
   59741: result <= 12'b110000111000;
   59742: result <= 12'b110000111000;
   59743: result <= 12'b110000110111;
   59744: result <= 12'b110000110111;
   59745: result <= 12'b110000110111;
   59746: result <= 12'b110000110111;
   59747: result <= 12'b110000110111;
   59748: result <= 12'b110000110111;
   59749: result <= 12'b110000110110;
   59750: result <= 12'b110000110110;
   59751: result <= 12'b110000110110;
   59752: result <= 12'b110000110110;
   59753: result <= 12'b110000110110;
   59754: result <= 12'b110000110110;
   59755: result <= 12'b110000110101;
   59756: result <= 12'b110000110101;
   59757: result <= 12'b110000110101;
   59758: result <= 12'b110000110101;
   59759: result <= 12'b110000110101;
   59760: result <= 12'b110000110101;
   59761: result <= 12'b110000110100;
   59762: result <= 12'b110000110100;
   59763: result <= 12'b110000110100;
   59764: result <= 12'b110000110100;
   59765: result <= 12'b110000110100;
   59766: result <= 12'b110000110100;
   59767: result <= 12'b110000110011;
   59768: result <= 12'b110000110011;
   59769: result <= 12'b110000110011;
   59770: result <= 12'b110000110011;
   59771: result <= 12'b110000110011;
   59772: result <= 12'b110000110011;
   59773: result <= 12'b110000110010;
   59774: result <= 12'b110000110010;
   59775: result <= 12'b110000110010;
   59776: result <= 12'b110000110010;
   59777: result <= 12'b110000110010;
   59778: result <= 12'b110000110010;
   59779: result <= 12'b110000110001;
   59780: result <= 12'b110000110001;
   59781: result <= 12'b110000110001;
   59782: result <= 12'b110000110001;
   59783: result <= 12'b110000110001;
   59784: result <= 12'b110000110001;
   59785: result <= 12'b110000110000;
   59786: result <= 12'b110000110000;
   59787: result <= 12'b110000110000;
   59788: result <= 12'b110000110000;
   59789: result <= 12'b110000110000;
   59790: result <= 12'b110000110000;
   59791: result <= 12'b110000101111;
   59792: result <= 12'b110000101111;
   59793: result <= 12'b110000101111;
   59794: result <= 12'b110000101111;
   59795: result <= 12'b110000101111;
   59796: result <= 12'b110000101111;
   59797: result <= 12'b110000101110;
   59798: result <= 12'b110000101110;
   59799: result <= 12'b110000101110;
   59800: result <= 12'b110000101110;
   59801: result <= 12'b110000101110;
   59802: result <= 12'b110000101110;
   59803: result <= 12'b110000101101;
   59804: result <= 12'b110000101101;
   59805: result <= 12'b110000101101;
   59806: result <= 12'b110000101101;
   59807: result <= 12'b110000101101;
   59808: result <= 12'b110000101101;
   59809: result <= 12'b110000101100;
   59810: result <= 12'b110000101100;
   59811: result <= 12'b110000101100;
   59812: result <= 12'b110000101100;
   59813: result <= 12'b110000101100;
   59814: result <= 12'b110000101100;
   59815: result <= 12'b110000101011;
   59816: result <= 12'b110000101011;
   59817: result <= 12'b110000101011;
   59818: result <= 12'b110000101011;
   59819: result <= 12'b110000101011;
   59820: result <= 12'b110000101010;
   59821: result <= 12'b110000101010;
   59822: result <= 12'b110000101010;
   59823: result <= 12'b110000101010;
   59824: result <= 12'b110000101010;
   59825: result <= 12'b110000101010;
   59826: result <= 12'b110000101001;
   59827: result <= 12'b110000101001;
   59828: result <= 12'b110000101001;
   59829: result <= 12'b110000101001;
   59830: result <= 12'b110000101001;
   59831: result <= 12'b110000101001;
   59832: result <= 12'b110000101000;
   59833: result <= 12'b110000101000;
   59834: result <= 12'b110000101000;
   59835: result <= 12'b110000101000;
   59836: result <= 12'b110000101000;
   59837: result <= 12'b110000101000;
   59838: result <= 12'b110000100111;
   59839: result <= 12'b110000100111;
   59840: result <= 12'b110000100111;
   59841: result <= 12'b110000100111;
   59842: result <= 12'b110000100111;
   59843: result <= 12'b110000100111;
   59844: result <= 12'b110000100110;
   59845: result <= 12'b110000100110;
   59846: result <= 12'b110000100110;
   59847: result <= 12'b110000100110;
   59848: result <= 12'b110000100110;
   59849: result <= 12'b110000100110;
   59850: result <= 12'b110000100101;
   59851: result <= 12'b110000100101;
   59852: result <= 12'b110000100101;
   59853: result <= 12'b110000100101;
   59854: result <= 12'b110000100101;
   59855: result <= 12'b110000100101;
   59856: result <= 12'b110000100100;
   59857: result <= 12'b110000100100;
   59858: result <= 12'b110000100100;
   59859: result <= 12'b110000100100;
   59860: result <= 12'b110000100100;
   59861: result <= 12'b110000100100;
   59862: result <= 12'b110000100011;
   59863: result <= 12'b110000100011;
   59864: result <= 12'b110000100011;
   59865: result <= 12'b110000100011;
   59866: result <= 12'b110000100011;
   59867: result <= 12'b110000100011;
   59868: result <= 12'b110000100010;
   59869: result <= 12'b110000100010;
   59870: result <= 12'b110000100010;
   59871: result <= 12'b110000100010;
   59872: result <= 12'b110000100010;
   59873: result <= 12'b110000100010;
   59874: result <= 12'b110000100001;
   59875: result <= 12'b110000100001;
   59876: result <= 12'b110000100001;
   59877: result <= 12'b110000100001;
   59878: result <= 12'b110000100001;
   59879: result <= 12'b110000100001;
   59880: result <= 12'b110000100000;
   59881: result <= 12'b110000100000;
   59882: result <= 12'b110000100000;
   59883: result <= 12'b110000100000;
   59884: result <= 12'b110000100000;
   59885: result <= 12'b110000100000;
   59886: result <= 12'b110000011111;
   59887: result <= 12'b110000011111;
   59888: result <= 12'b110000011111;
   59889: result <= 12'b110000011111;
   59890: result <= 12'b110000011111;
   59891: result <= 12'b110000011111;
   59892: result <= 12'b110000011110;
   59893: result <= 12'b110000011110;
   59894: result <= 12'b110000011110;
   59895: result <= 12'b110000011110;
   59896: result <= 12'b110000011110;
   59897: result <= 12'b110000011110;
   59898: result <= 12'b110000011101;
   59899: result <= 12'b110000011101;
   59900: result <= 12'b110000011101;
   59901: result <= 12'b110000011101;
   59902: result <= 12'b110000011101;
   59903: result <= 12'b110000011101;
   59904: result <= 12'b110000011100;
   59905: result <= 12'b110000011100;
   59906: result <= 12'b110000011100;
   59907: result <= 12'b110000011100;
   59908: result <= 12'b110000011100;
   59909: result <= 12'b110000011100;
   59910: result <= 12'b110000011011;
   59911: result <= 12'b110000011011;
   59912: result <= 12'b110000011011;
   59913: result <= 12'b110000011011;
   59914: result <= 12'b110000011011;
   59915: result <= 12'b110000011011;
   59916: result <= 12'b110000011010;
   59917: result <= 12'b110000011010;
   59918: result <= 12'b110000011010;
   59919: result <= 12'b110000011010;
   59920: result <= 12'b110000011010;
   59921: result <= 12'b110000011010;
   59922: result <= 12'b110000011001;
   59923: result <= 12'b110000011001;
   59924: result <= 12'b110000011001;
   59925: result <= 12'b110000011001;
   59926: result <= 12'b110000011001;
   59927: result <= 12'b110000011001;
   59928: result <= 12'b110000011000;
   59929: result <= 12'b110000011000;
   59930: result <= 12'b110000011000;
   59931: result <= 12'b110000011000;
   59932: result <= 12'b110000011000;
   59933: result <= 12'b110000010111;
   59934: result <= 12'b110000010111;
   59935: result <= 12'b110000010111;
   59936: result <= 12'b110000010111;
   59937: result <= 12'b110000010111;
   59938: result <= 12'b110000010111;
   59939: result <= 12'b110000010110;
   59940: result <= 12'b110000010110;
   59941: result <= 12'b110000010110;
   59942: result <= 12'b110000010110;
   59943: result <= 12'b110000010110;
   59944: result <= 12'b110000010110;
   59945: result <= 12'b110000010101;
   59946: result <= 12'b110000010101;
   59947: result <= 12'b110000010101;
   59948: result <= 12'b110000010101;
   59949: result <= 12'b110000010101;
   59950: result <= 12'b110000010101;
   59951: result <= 12'b110000010100;
   59952: result <= 12'b110000010100;
   59953: result <= 12'b110000010100;
   59954: result <= 12'b110000010100;
   59955: result <= 12'b110000010100;
   59956: result <= 12'b110000010100;
   59957: result <= 12'b110000010011;
   59958: result <= 12'b110000010011;
   59959: result <= 12'b110000010011;
   59960: result <= 12'b110000010011;
   59961: result <= 12'b110000010011;
   59962: result <= 12'b110000010011;
   59963: result <= 12'b110000010010;
   59964: result <= 12'b110000010010;
   59965: result <= 12'b110000010010;
   59966: result <= 12'b110000010010;
   59967: result <= 12'b110000010010;
   59968: result <= 12'b110000010010;
   59969: result <= 12'b110000010001;
   59970: result <= 12'b110000010001;
   59971: result <= 12'b110000010001;
   59972: result <= 12'b110000010001;
   59973: result <= 12'b110000010001;
   59974: result <= 12'b110000010001;
   59975: result <= 12'b110000010000;
   59976: result <= 12'b110000010000;
   59977: result <= 12'b110000010000;
   59978: result <= 12'b110000010000;
   59979: result <= 12'b110000010000;
   59980: result <= 12'b110000010000;
   59981: result <= 12'b110000001111;
   59982: result <= 12'b110000001111;
   59983: result <= 12'b110000001111;
   59984: result <= 12'b110000001111;
   59985: result <= 12'b110000001111;
   59986: result <= 12'b110000001111;
   59987: result <= 12'b110000001110;
   59988: result <= 12'b110000001110;
   59989: result <= 12'b110000001110;
   59990: result <= 12'b110000001110;
   59991: result <= 12'b110000001110;
   59992: result <= 12'b110000001110;
   59993: result <= 12'b110000001101;
   59994: result <= 12'b110000001101;
   59995: result <= 12'b110000001101;
   59996: result <= 12'b110000001101;
   59997: result <= 12'b110000001101;
   59998: result <= 12'b110000001101;
   59999: result <= 12'b110000001100;
   60000: result <= 12'b110000001100;
   60001: result <= 12'b110000001100;
   60002: result <= 12'b110000001100;
   60003: result <= 12'b110000001100;
   60004: result <= 12'b110000001011;
   60005: result <= 12'b110000001011;
   60006: result <= 12'b110000001011;
   60007: result <= 12'b110000001011;
   60008: result <= 12'b110000001011;
   60009: result <= 12'b110000001011;
   60010: result <= 12'b110000001010;
   60011: result <= 12'b110000001010;
   60012: result <= 12'b110000001010;
   60013: result <= 12'b110000001010;
   60014: result <= 12'b110000001010;
   60015: result <= 12'b110000001010;
   60016: result <= 12'b110000001001;
   60017: result <= 12'b110000001001;
   60018: result <= 12'b110000001001;
   60019: result <= 12'b110000001001;
   60020: result <= 12'b110000001001;
   60021: result <= 12'b110000001001;
   60022: result <= 12'b110000001000;
   60023: result <= 12'b110000001000;
   60024: result <= 12'b110000001000;
   60025: result <= 12'b110000001000;
   60026: result <= 12'b110000001000;
   60027: result <= 12'b110000001000;
   60028: result <= 12'b110000000111;
   60029: result <= 12'b110000000111;
   60030: result <= 12'b110000000111;
   60031: result <= 12'b110000000111;
   60032: result <= 12'b110000000111;
   60033: result <= 12'b110000000111;
   60034: result <= 12'b110000000110;
   60035: result <= 12'b110000000110;
   60036: result <= 12'b110000000110;
   60037: result <= 12'b110000000110;
   60038: result <= 12'b110000000110;
   60039: result <= 12'b110000000110;
   60040: result <= 12'b110000000101;
   60041: result <= 12'b110000000101;
   60042: result <= 12'b110000000101;
   60043: result <= 12'b110000000101;
   60044: result <= 12'b110000000101;
   60045: result <= 12'b110000000101;
   60046: result <= 12'b110000000100;
   60047: result <= 12'b110000000100;
   60048: result <= 12'b110000000100;
   60049: result <= 12'b110000000100;
   60050: result <= 12'b110000000100;
   60051: result <= 12'b110000000100;
   60052: result <= 12'b110000000011;
   60053: result <= 12'b110000000011;
   60054: result <= 12'b110000000011;
   60055: result <= 12'b110000000011;
   60056: result <= 12'b110000000011;
   60057: result <= 12'b110000000011;
   60058: result <= 12'b110000000010;
   60059: result <= 12'b110000000010;
   60060: result <= 12'b110000000010;
   60061: result <= 12'b110000000010;
   60062: result <= 12'b110000000010;
   60063: result <= 12'b110000000001;
   60064: result <= 12'b110000000001;
   60065: result <= 12'b110000000001;
   60066: result <= 12'b110000000001;
   60067: result <= 12'b110000000001;
   60068: result <= 12'b110000000001;
   60069: result <= 12'b110000000000;
   60070: result <= 12'b110000000000;
   60071: result <= 12'b110000000000;
   60072: result <= 12'b110000000000;
   60073: result <= 12'b110000000000;
   60074: result <= 12'b110000000000;
   60075: result <= 12'b111111111111;
   60076: result <= 12'b111111111111;
   60077: result <= 12'b111111111111;
   60078: result <= 12'b111111111111;
   60079: result <= 12'b111111111111;
   60080: result <= 12'b111111111111;
   60081: result <= 12'b111111111110;
   60082: result <= 12'b111111111110;
   60083: result <= 12'b111111111110;
   60084: result <= 12'b111111111110;
   60085: result <= 12'b111111111110;
   60086: result <= 12'b111111111110;
   60087: result <= 12'b111111111101;
   60088: result <= 12'b111111111101;
   60089: result <= 12'b111111111101;
   60090: result <= 12'b111111111101;
   60091: result <= 12'b111111111101;
   60092: result <= 12'b111111111101;
   60093: result <= 12'b111111111100;
   60094: result <= 12'b111111111100;
   60095: result <= 12'b111111111100;
   60096: result <= 12'b111111111100;
   60097: result <= 12'b111111111100;
   60098: result <= 12'b111111111100;
   60099: result <= 12'b111111111011;
   60100: result <= 12'b111111111011;
   60101: result <= 12'b111111111011;
   60102: result <= 12'b111111111011;
   60103: result <= 12'b111111111011;
   60104: result <= 12'b111111111011;
   60105: result <= 12'b111111111010;
   60106: result <= 12'b111111111010;
   60107: result <= 12'b111111111010;
   60108: result <= 12'b111111111010;
   60109: result <= 12'b111111111010;
   60110: result <= 12'b111111111001;
   60111: result <= 12'b111111111001;
   60112: result <= 12'b111111111001;
   60113: result <= 12'b111111111001;
   60114: result <= 12'b111111111001;
   60115: result <= 12'b111111111001;
   60116: result <= 12'b111111111000;
   60117: result <= 12'b111111111000;
   60118: result <= 12'b111111111000;
   60119: result <= 12'b111111111000;
   60120: result <= 12'b111111111000;
   60121: result <= 12'b111111111000;
   60122: result <= 12'b111111110111;
   60123: result <= 12'b111111110111;
   60124: result <= 12'b111111110111;
   60125: result <= 12'b111111110111;
   60126: result <= 12'b111111110111;
   60127: result <= 12'b111111110111;
   60128: result <= 12'b111111110110;
   60129: result <= 12'b111111110110;
   60130: result <= 12'b111111110110;
   60131: result <= 12'b111111110110;
   60132: result <= 12'b111111110110;
   60133: result <= 12'b111111110110;
   60134: result <= 12'b111111110101;
   60135: result <= 12'b111111110101;
   60136: result <= 12'b111111110101;
   60137: result <= 12'b111111110101;
   60138: result <= 12'b111111110101;
   60139: result <= 12'b111111110101;
   60140: result <= 12'b111111110100;
   60141: result <= 12'b111111110100;
   60142: result <= 12'b111111110100;
   60143: result <= 12'b111111110100;
   60144: result <= 12'b111111110100;
   60145: result <= 12'b111111110100;
   60146: result <= 12'b111111110011;
   60147: result <= 12'b111111110011;
   60148: result <= 12'b111111110011;
   60149: result <= 12'b111111110011;
   60150: result <= 12'b111111110011;
   60151: result <= 12'b111111110010;
   60152: result <= 12'b111111110010;
   60153: result <= 12'b111111110010;
   60154: result <= 12'b111111110010;
   60155: result <= 12'b111111110010;
   60156: result <= 12'b111111110010;
   60157: result <= 12'b111111110001;
   60158: result <= 12'b111111110001;
   60159: result <= 12'b111111110001;
   60160: result <= 12'b111111110001;
   60161: result <= 12'b111111110001;
   60162: result <= 12'b111111110001;
   60163: result <= 12'b111111110000;
   60164: result <= 12'b111111110000;
   60165: result <= 12'b111111110000;
   60166: result <= 12'b111111110000;
   60167: result <= 12'b111111110000;
   60168: result <= 12'b111111110000;
   60169: result <= 12'b111111101111;
   60170: result <= 12'b111111101111;
   60171: result <= 12'b111111101111;
   60172: result <= 12'b111111101111;
   60173: result <= 12'b111111101111;
   60174: result <= 12'b111111101111;
   60175: result <= 12'b111111101110;
   60176: result <= 12'b111111101110;
   60177: result <= 12'b111111101110;
   60178: result <= 12'b111111101110;
   60179: result <= 12'b111111101110;
   60180: result <= 12'b111111101110;
   60181: result <= 12'b111111101101;
   60182: result <= 12'b111111101101;
   60183: result <= 12'b111111101101;
   60184: result <= 12'b111111101101;
   60185: result <= 12'b111111101101;
   60186: result <= 12'b111111101101;
   60187: result <= 12'b111111101100;
   60188: result <= 12'b111111101100;
   60189: result <= 12'b111111101100;
   60190: result <= 12'b111111101100;
   60191: result <= 12'b111111101100;
   60192: result <= 12'b111111101011;
   60193: result <= 12'b111111101011;
   60194: result <= 12'b111111101011;
   60195: result <= 12'b111111101011;
   60196: result <= 12'b111111101011;
   60197: result <= 12'b111111101011;
   60198: result <= 12'b111111101010;
   60199: result <= 12'b111111101010;
   60200: result <= 12'b111111101010;
   60201: result <= 12'b111111101010;
   60202: result <= 12'b111111101010;
   60203: result <= 12'b111111101010;
   60204: result <= 12'b111111101001;
   60205: result <= 12'b111111101001;
   60206: result <= 12'b111111101001;
   60207: result <= 12'b111111101001;
   60208: result <= 12'b111111101001;
   60209: result <= 12'b111111101001;
   60210: result <= 12'b111111101000;
   60211: result <= 12'b111111101000;
   60212: result <= 12'b111111101000;
   60213: result <= 12'b111111101000;
   60214: result <= 12'b111111101000;
   60215: result <= 12'b111111101000;
   60216: result <= 12'b111111100111;
   60217: result <= 12'b111111100111;
   60218: result <= 12'b111111100111;
   60219: result <= 12'b111111100111;
   60220: result <= 12'b111111100111;
   60221: result <= 12'b111111100111;
   60222: result <= 12'b111111100110;
   60223: result <= 12'b111111100110;
   60224: result <= 12'b111111100110;
   60225: result <= 12'b111111100110;
   60226: result <= 12'b111111100110;
   60227: result <= 12'b111111100101;
   60228: result <= 12'b111111100101;
   60229: result <= 12'b111111100101;
   60230: result <= 12'b111111100101;
   60231: result <= 12'b111111100101;
   60232: result <= 12'b111111100101;
   60233: result <= 12'b111111100100;
   60234: result <= 12'b111111100100;
   60235: result <= 12'b111111100100;
   60236: result <= 12'b111111100100;
   60237: result <= 12'b111111100100;
   60238: result <= 12'b111111100100;
   60239: result <= 12'b111111100011;
   60240: result <= 12'b111111100011;
   60241: result <= 12'b111111100011;
   60242: result <= 12'b111111100011;
   60243: result <= 12'b111111100011;
   60244: result <= 12'b111111100011;
   60245: result <= 12'b111111100010;
   60246: result <= 12'b111111100010;
   60247: result <= 12'b111111100010;
   60248: result <= 12'b111111100010;
   60249: result <= 12'b111111100010;
   60250: result <= 12'b111111100010;
   60251: result <= 12'b111111100001;
   60252: result <= 12'b111111100001;
   60253: result <= 12'b111111100001;
   60254: result <= 12'b111111100001;
   60255: result <= 12'b111111100001;
   60256: result <= 12'b111111100001;
   60257: result <= 12'b111111100000;
   60258: result <= 12'b111111100000;
   60259: result <= 12'b111111100000;
   60260: result <= 12'b111111100000;
   60261: result <= 12'b111111100000;
   60262: result <= 12'b111111011111;
   60263: result <= 12'b111111011111;
   60264: result <= 12'b111111011111;
   60265: result <= 12'b111111011111;
   60266: result <= 12'b111111011111;
   60267: result <= 12'b111111011111;
   60268: result <= 12'b111111011110;
   60269: result <= 12'b111111011110;
   60270: result <= 12'b111111011110;
   60271: result <= 12'b111111011110;
   60272: result <= 12'b111111011110;
   60273: result <= 12'b111111011110;
   60274: result <= 12'b111111011101;
   60275: result <= 12'b111111011101;
   60276: result <= 12'b111111011101;
   60277: result <= 12'b111111011101;
   60278: result <= 12'b111111011101;
   60279: result <= 12'b111111011101;
   60280: result <= 12'b111111011100;
   60281: result <= 12'b111111011100;
   60282: result <= 12'b111111011100;
   60283: result <= 12'b111111011100;
   60284: result <= 12'b111111011100;
   60285: result <= 12'b111111011100;
   60286: result <= 12'b111111011011;
   60287: result <= 12'b111111011011;
   60288: result <= 12'b111111011011;
   60289: result <= 12'b111111011011;
   60290: result <= 12'b111111011011;
   60291: result <= 12'b111111011010;
   60292: result <= 12'b111111011010;
   60293: result <= 12'b111111011010;
   60294: result <= 12'b111111011010;
   60295: result <= 12'b111111011010;
   60296: result <= 12'b111111011010;
   60297: result <= 12'b111111011001;
   60298: result <= 12'b111111011001;
   60299: result <= 12'b111111011001;
   60300: result <= 12'b111111011001;
   60301: result <= 12'b111111011001;
   60302: result <= 12'b111111011001;
   60303: result <= 12'b111111011000;
   60304: result <= 12'b111111011000;
   60305: result <= 12'b111111011000;
   60306: result <= 12'b111111011000;
   60307: result <= 12'b111111011000;
   60308: result <= 12'b111111011000;
   60309: result <= 12'b111111010111;
   60310: result <= 12'b111111010111;
   60311: result <= 12'b111111010111;
   60312: result <= 12'b111111010111;
   60313: result <= 12'b111111010111;
   60314: result <= 12'b111111010111;
   60315: result <= 12'b111111010110;
   60316: result <= 12'b111111010110;
   60317: result <= 12'b111111010110;
   60318: result <= 12'b111111010110;
   60319: result <= 12'b111111010110;
   60320: result <= 12'b111111010110;
   60321: result <= 12'b111111010101;
   60322: result <= 12'b111111010101;
   60323: result <= 12'b111111010101;
   60324: result <= 12'b111111010101;
   60325: result <= 12'b111111010101;
   60326: result <= 12'b111111010100;
   60327: result <= 12'b111111010100;
   60328: result <= 12'b111111010100;
   60329: result <= 12'b111111010100;
   60330: result <= 12'b111111010100;
   60331: result <= 12'b111111010100;
   60332: result <= 12'b111111010011;
   60333: result <= 12'b111111010011;
   60334: result <= 12'b111111010011;
   60335: result <= 12'b111111010011;
   60336: result <= 12'b111111010011;
   60337: result <= 12'b111111010011;
   60338: result <= 12'b111111010010;
   60339: result <= 12'b111111010010;
   60340: result <= 12'b111111010010;
   60341: result <= 12'b111111010010;
   60342: result <= 12'b111111010010;
   60343: result <= 12'b111111010010;
   60344: result <= 12'b111111010001;
   60345: result <= 12'b111111010001;
   60346: result <= 12'b111111010001;
   60347: result <= 12'b111111010001;
   60348: result <= 12'b111111010001;
   60349: result <= 12'b111111010001;
   60350: result <= 12'b111111010000;
   60351: result <= 12'b111111010000;
   60352: result <= 12'b111111010000;
   60353: result <= 12'b111111010000;
   60354: result <= 12'b111111010000;
   60355: result <= 12'b111111001111;
   60356: result <= 12'b111111001111;
   60357: result <= 12'b111111001111;
   60358: result <= 12'b111111001111;
   60359: result <= 12'b111111001111;
   60360: result <= 12'b111111001111;
   60361: result <= 12'b111111001110;
   60362: result <= 12'b111111001110;
   60363: result <= 12'b111111001110;
   60364: result <= 12'b111111001110;
   60365: result <= 12'b111111001110;
   60366: result <= 12'b111111001110;
   60367: result <= 12'b111111001101;
   60368: result <= 12'b111111001101;
   60369: result <= 12'b111111001101;
   60370: result <= 12'b111111001101;
   60371: result <= 12'b111111001101;
   60372: result <= 12'b111111001101;
   60373: result <= 12'b111111001100;
   60374: result <= 12'b111111001100;
   60375: result <= 12'b111111001100;
   60376: result <= 12'b111111001100;
   60377: result <= 12'b111111001100;
   60378: result <= 12'b111111001011;
   60379: result <= 12'b111111001011;
   60380: result <= 12'b111111001011;
   60381: result <= 12'b111111001011;
   60382: result <= 12'b111111001011;
   60383: result <= 12'b111111001011;
   60384: result <= 12'b111111001010;
   60385: result <= 12'b111111001010;
   60386: result <= 12'b111111001010;
   60387: result <= 12'b111111001010;
   60388: result <= 12'b111111001010;
   60389: result <= 12'b111111001010;
   60390: result <= 12'b111111001001;
   60391: result <= 12'b111111001001;
   60392: result <= 12'b111111001001;
   60393: result <= 12'b111111001001;
   60394: result <= 12'b111111001001;
   60395: result <= 12'b111111001001;
   60396: result <= 12'b111111001000;
   60397: result <= 12'b111111001000;
   60398: result <= 12'b111111001000;
   60399: result <= 12'b111111001000;
   60400: result <= 12'b111111001000;
   60401: result <= 12'b111111001000;
   60402: result <= 12'b111111000111;
   60403: result <= 12'b111111000111;
   60404: result <= 12'b111111000111;
   60405: result <= 12'b111111000111;
   60406: result <= 12'b111111000111;
   60407: result <= 12'b111111000110;
   60408: result <= 12'b111111000110;
   60409: result <= 12'b111111000110;
   60410: result <= 12'b111111000110;
   60411: result <= 12'b111111000110;
   60412: result <= 12'b111111000110;
   60413: result <= 12'b111111000101;
   60414: result <= 12'b111111000101;
   60415: result <= 12'b111111000101;
   60416: result <= 12'b111111000101;
   60417: result <= 12'b111111000101;
   60418: result <= 12'b111111000101;
   60419: result <= 12'b111111000100;
   60420: result <= 12'b111111000100;
   60421: result <= 12'b111111000100;
   60422: result <= 12'b111111000100;
   60423: result <= 12'b111111000100;
   60424: result <= 12'b111111000100;
   60425: result <= 12'b111111000011;
   60426: result <= 12'b111111000011;
   60427: result <= 12'b111111000011;
   60428: result <= 12'b111111000011;
   60429: result <= 12'b111111000011;
   60430: result <= 12'b111111000010;
   60431: result <= 12'b111111000010;
   60432: result <= 12'b111111000010;
   60433: result <= 12'b111111000010;
   60434: result <= 12'b111111000010;
   60435: result <= 12'b111111000010;
   60436: result <= 12'b111111000001;
   60437: result <= 12'b111111000001;
   60438: result <= 12'b111111000001;
   60439: result <= 12'b111111000001;
   60440: result <= 12'b111111000001;
   60441: result <= 12'b111111000001;
   60442: result <= 12'b111111000000;
   60443: result <= 12'b111111000000;
   60444: result <= 12'b111111000000;
   60445: result <= 12'b111111000000;
   60446: result <= 12'b111111000000;
   60447: result <= 12'b111111000000;
   60448: result <= 12'b111110111111;
   60449: result <= 12'b111110111111;
   60450: result <= 12'b111110111111;
   60451: result <= 12'b111110111111;
   60452: result <= 12'b111110111111;
   60453: result <= 12'b111110111111;
   60454: result <= 12'b111110111110;
   60455: result <= 12'b111110111110;
   60456: result <= 12'b111110111110;
   60457: result <= 12'b111110111110;
   60458: result <= 12'b111110111110;
   60459: result <= 12'b111110111101;
   60460: result <= 12'b111110111101;
   60461: result <= 12'b111110111101;
   60462: result <= 12'b111110111101;
   60463: result <= 12'b111110111101;
   60464: result <= 12'b111110111101;
   60465: result <= 12'b111110111100;
   60466: result <= 12'b111110111100;
   60467: result <= 12'b111110111100;
   60468: result <= 12'b111110111100;
   60469: result <= 12'b111110111100;
   60470: result <= 12'b111110111100;
   60471: result <= 12'b111110111011;
   60472: result <= 12'b111110111011;
   60473: result <= 12'b111110111011;
   60474: result <= 12'b111110111011;
   60475: result <= 12'b111110111011;
   60476: result <= 12'b111110111011;
   60477: result <= 12'b111110111010;
   60478: result <= 12'b111110111010;
   60479: result <= 12'b111110111010;
   60480: result <= 12'b111110111010;
   60481: result <= 12'b111110111010;
   60482: result <= 12'b111110111001;
   60483: result <= 12'b111110111001;
   60484: result <= 12'b111110111001;
   60485: result <= 12'b111110111001;
   60486: result <= 12'b111110111001;
   60487: result <= 12'b111110111001;
   60488: result <= 12'b111110111000;
   60489: result <= 12'b111110111000;
   60490: result <= 12'b111110111000;
   60491: result <= 12'b111110111000;
   60492: result <= 12'b111110111000;
   60493: result <= 12'b111110111000;
   60494: result <= 12'b111110110111;
   60495: result <= 12'b111110110111;
   60496: result <= 12'b111110110111;
   60497: result <= 12'b111110110111;
   60498: result <= 12'b111110110111;
   60499: result <= 12'b111110110111;
   60500: result <= 12'b111110110110;
   60501: result <= 12'b111110110110;
   60502: result <= 12'b111110110110;
   60503: result <= 12'b111110110110;
   60504: result <= 12'b111110110110;
   60505: result <= 12'b111110110101;
   60506: result <= 12'b111110110101;
   60507: result <= 12'b111110110101;
   60508: result <= 12'b111110110101;
   60509: result <= 12'b111110110101;
   60510: result <= 12'b111110110101;
   60511: result <= 12'b111110110100;
   60512: result <= 12'b111110110100;
   60513: result <= 12'b111110110100;
   60514: result <= 12'b111110110100;
   60515: result <= 12'b111110110100;
   60516: result <= 12'b111110110100;
   60517: result <= 12'b111110110011;
   60518: result <= 12'b111110110011;
   60519: result <= 12'b111110110011;
   60520: result <= 12'b111110110011;
   60521: result <= 12'b111110110011;
   60522: result <= 12'b111110110011;
   60523: result <= 12'b111110110010;
   60524: result <= 12'b111110110010;
   60525: result <= 12'b111110110010;
   60526: result <= 12'b111110110010;
   60527: result <= 12'b111110110010;
   60528: result <= 12'b111110110001;
   60529: result <= 12'b111110110001;
   60530: result <= 12'b111110110001;
   60531: result <= 12'b111110110001;
   60532: result <= 12'b111110110001;
   60533: result <= 12'b111110110001;
   60534: result <= 12'b111110110000;
   60535: result <= 12'b111110110000;
   60536: result <= 12'b111110110000;
   60537: result <= 12'b111110110000;
   60538: result <= 12'b111110110000;
   60539: result <= 12'b111110110000;
   60540: result <= 12'b111110101111;
   60541: result <= 12'b111110101111;
   60542: result <= 12'b111110101111;
   60543: result <= 12'b111110101111;
   60544: result <= 12'b111110101111;
   60545: result <= 12'b111110101111;
   60546: result <= 12'b111110101110;
   60547: result <= 12'b111110101110;
   60548: result <= 12'b111110101110;
   60549: result <= 12'b111110101110;
   60550: result <= 12'b111110101110;
   60551: result <= 12'b111110101101;
   60552: result <= 12'b111110101101;
   60553: result <= 12'b111110101101;
   60554: result <= 12'b111110101101;
   60555: result <= 12'b111110101101;
   60556: result <= 12'b111110101101;
   60557: result <= 12'b111110101100;
   60558: result <= 12'b111110101100;
   60559: result <= 12'b111110101100;
   60560: result <= 12'b111110101100;
   60561: result <= 12'b111110101100;
   60562: result <= 12'b111110101100;
   60563: result <= 12'b111110101011;
   60564: result <= 12'b111110101011;
   60565: result <= 12'b111110101011;
   60566: result <= 12'b111110101011;
   60567: result <= 12'b111110101011;
   60568: result <= 12'b111110101010;
   60569: result <= 12'b111110101010;
   60570: result <= 12'b111110101010;
   60571: result <= 12'b111110101010;
   60572: result <= 12'b111110101010;
   60573: result <= 12'b111110101010;
   60574: result <= 12'b111110101001;
   60575: result <= 12'b111110101001;
   60576: result <= 12'b111110101001;
   60577: result <= 12'b111110101001;
   60578: result <= 12'b111110101001;
   60579: result <= 12'b111110101001;
   60580: result <= 12'b111110101000;
   60581: result <= 12'b111110101000;
   60582: result <= 12'b111110101000;
   60583: result <= 12'b111110101000;
   60584: result <= 12'b111110101000;
   60585: result <= 12'b111110101000;
   60586: result <= 12'b111110100111;
   60587: result <= 12'b111110100111;
   60588: result <= 12'b111110100111;
   60589: result <= 12'b111110100111;
   60590: result <= 12'b111110100111;
   60591: result <= 12'b111110100110;
   60592: result <= 12'b111110100110;
   60593: result <= 12'b111110100110;
   60594: result <= 12'b111110100110;
   60595: result <= 12'b111110100110;
   60596: result <= 12'b111110100110;
   60597: result <= 12'b111110100101;
   60598: result <= 12'b111110100101;
   60599: result <= 12'b111110100101;
   60600: result <= 12'b111110100101;
   60601: result <= 12'b111110100101;
   60602: result <= 12'b111110100101;
   60603: result <= 12'b111110100100;
   60604: result <= 12'b111110100100;
   60605: result <= 12'b111110100100;
   60606: result <= 12'b111110100100;
   60607: result <= 12'b111110100100;
   60608: result <= 12'b111110100100;
   60609: result <= 12'b111110100011;
   60610: result <= 12'b111110100011;
   60611: result <= 12'b111110100011;
   60612: result <= 12'b111110100011;
   60613: result <= 12'b111110100011;
   60614: result <= 12'b111110100010;
   60615: result <= 12'b111110100010;
   60616: result <= 12'b111110100010;
   60617: result <= 12'b111110100010;
   60618: result <= 12'b111110100010;
   60619: result <= 12'b111110100010;
   60620: result <= 12'b111110100001;
   60621: result <= 12'b111110100001;
   60622: result <= 12'b111110100001;
   60623: result <= 12'b111110100001;
   60624: result <= 12'b111110100001;
   60625: result <= 12'b111110100001;
   60626: result <= 12'b111110100000;
   60627: result <= 12'b111110100000;
   60628: result <= 12'b111110100000;
   60629: result <= 12'b111110100000;
   60630: result <= 12'b111110100000;
   60631: result <= 12'b111110011111;
   60632: result <= 12'b111110011111;
   60633: result <= 12'b111110011111;
   60634: result <= 12'b111110011111;
   60635: result <= 12'b111110011111;
   60636: result <= 12'b111110011111;
   60637: result <= 12'b111110011110;
   60638: result <= 12'b111110011110;
   60639: result <= 12'b111110011110;
   60640: result <= 12'b111110011110;
   60641: result <= 12'b111110011110;
   60642: result <= 12'b111110011110;
   60643: result <= 12'b111110011101;
   60644: result <= 12'b111110011101;
   60645: result <= 12'b111110011101;
   60646: result <= 12'b111110011101;
   60647: result <= 12'b111110011101;
   60648: result <= 12'b111110011101;
   60649: result <= 12'b111110011100;
   60650: result <= 12'b111110011100;
   60651: result <= 12'b111110011100;
   60652: result <= 12'b111110011100;
   60653: result <= 12'b111110011100;
   60654: result <= 12'b111110011011;
   60655: result <= 12'b111110011011;
   60656: result <= 12'b111110011011;
   60657: result <= 12'b111110011011;
   60658: result <= 12'b111110011011;
   60659: result <= 12'b111110011011;
   60660: result <= 12'b111110011010;
   60661: result <= 12'b111110011010;
   60662: result <= 12'b111110011010;
   60663: result <= 12'b111110011010;
   60664: result <= 12'b111110011010;
   60665: result <= 12'b111110011010;
   60666: result <= 12'b111110011001;
   60667: result <= 12'b111110011001;
   60668: result <= 12'b111110011001;
   60669: result <= 12'b111110011001;
   60670: result <= 12'b111110011001;
   60671: result <= 12'b111110011000;
   60672: result <= 12'b111110011000;
   60673: result <= 12'b111110011000;
   60674: result <= 12'b111110011000;
   60675: result <= 12'b111110011000;
   60676: result <= 12'b111110011000;
   60677: result <= 12'b111110010111;
   60678: result <= 12'b111110010111;
   60679: result <= 12'b111110010111;
   60680: result <= 12'b111110010111;
   60681: result <= 12'b111110010111;
   60682: result <= 12'b111110010111;
   60683: result <= 12'b111110010110;
   60684: result <= 12'b111110010110;
   60685: result <= 12'b111110010110;
   60686: result <= 12'b111110010110;
   60687: result <= 12'b111110010110;
   60688: result <= 12'b111110010101;
   60689: result <= 12'b111110010101;
   60690: result <= 12'b111110010101;
   60691: result <= 12'b111110010101;
   60692: result <= 12'b111110010101;
   60693: result <= 12'b111110010101;
   60694: result <= 12'b111110010100;
   60695: result <= 12'b111110010100;
   60696: result <= 12'b111110010100;
   60697: result <= 12'b111110010100;
   60698: result <= 12'b111110010100;
   60699: result <= 12'b111110010100;
   60700: result <= 12'b111110010011;
   60701: result <= 12'b111110010011;
   60702: result <= 12'b111110010011;
   60703: result <= 12'b111110010011;
   60704: result <= 12'b111110010011;
   60705: result <= 12'b111110010011;
   60706: result <= 12'b111110010010;
   60707: result <= 12'b111110010010;
   60708: result <= 12'b111110010010;
   60709: result <= 12'b111110010010;
   60710: result <= 12'b111110010010;
   60711: result <= 12'b111110010001;
   60712: result <= 12'b111110010001;
   60713: result <= 12'b111110010001;
   60714: result <= 12'b111110010001;
   60715: result <= 12'b111110010001;
   60716: result <= 12'b111110010001;
   60717: result <= 12'b111110010000;
   60718: result <= 12'b111110010000;
   60719: result <= 12'b111110010000;
   60720: result <= 12'b111110010000;
   60721: result <= 12'b111110010000;
   60722: result <= 12'b111110010000;
   60723: result <= 12'b111110001111;
   60724: result <= 12'b111110001111;
   60725: result <= 12'b111110001111;
   60726: result <= 12'b111110001111;
   60727: result <= 12'b111110001111;
   60728: result <= 12'b111110001110;
   60729: result <= 12'b111110001110;
   60730: result <= 12'b111110001110;
   60731: result <= 12'b111110001110;
   60732: result <= 12'b111110001110;
   60733: result <= 12'b111110001110;
   60734: result <= 12'b111110001101;
   60735: result <= 12'b111110001101;
   60736: result <= 12'b111110001101;
   60737: result <= 12'b111110001101;
   60738: result <= 12'b111110001101;
   60739: result <= 12'b111110001101;
   60740: result <= 12'b111110001100;
   60741: result <= 12'b111110001100;
   60742: result <= 12'b111110001100;
   60743: result <= 12'b111110001100;
   60744: result <= 12'b111110001100;
   60745: result <= 12'b111110001011;
   60746: result <= 12'b111110001011;
   60747: result <= 12'b111110001011;
   60748: result <= 12'b111110001011;
   60749: result <= 12'b111110001011;
   60750: result <= 12'b111110001011;
   60751: result <= 12'b111110001010;
   60752: result <= 12'b111110001010;
   60753: result <= 12'b111110001010;
   60754: result <= 12'b111110001010;
   60755: result <= 12'b111110001010;
   60756: result <= 12'b111110001010;
   60757: result <= 12'b111110001001;
   60758: result <= 12'b111110001001;
   60759: result <= 12'b111110001001;
   60760: result <= 12'b111110001001;
   60761: result <= 12'b111110001001;
   60762: result <= 12'b111110001000;
   60763: result <= 12'b111110001000;
   60764: result <= 12'b111110001000;
   60765: result <= 12'b111110001000;
   60766: result <= 12'b111110001000;
   60767: result <= 12'b111110001000;
   60768: result <= 12'b111110000111;
   60769: result <= 12'b111110000111;
   60770: result <= 12'b111110000111;
   60771: result <= 12'b111110000111;
   60772: result <= 12'b111110000111;
   60773: result <= 12'b111110000111;
   60774: result <= 12'b111110000110;
   60775: result <= 12'b111110000110;
   60776: result <= 12'b111110000110;
   60777: result <= 12'b111110000110;
   60778: result <= 12'b111110000110;
   60779: result <= 12'b111110000101;
   60780: result <= 12'b111110000101;
   60781: result <= 12'b111110000101;
   60782: result <= 12'b111110000101;
   60783: result <= 12'b111110000101;
   60784: result <= 12'b111110000101;
   60785: result <= 12'b111110000100;
   60786: result <= 12'b111110000100;
   60787: result <= 12'b111110000100;
   60788: result <= 12'b111110000100;
   60789: result <= 12'b111110000100;
   60790: result <= 12'b111110000100;
   60791: result <= 12'b111110000011;
   60792: result <= 12'b111110000011;
   60793: result <= 12'b111110000011;
   60794: result <= 12'b111110000011;
   60795: result <= 12'b111110000011;
   60796: result <= 12'b111110000010;
   60797: result <= 12'b111110000010;
   60798: result <= 12'b111110000010;
   60799: result <= 12'b111110000010;
   60800: result <= 12'b111110000010;
   60801: result <= 12'b111110000010;
   60802: result <= 12'b111110000001;
   60803: result <= 12'b111110000001;
   60804: result <= 12'b111110000001;
   60805: result <= 12'b111110000001;
   60806: result <= 12'b111110000001;
   60807: result <= 12'b111110000001;
   60808: result <= 12'b111110000000;
   60809: result <= 12'b111110000000;
   60810: result <= 12'b111110000000;
   60811: result <= 12'b111110000000;
   60812: result <= 12'b111110000000;
   60813: result <= 12'b111101111111;
   60814: result <= 12'b111101111111;
   60815: result <= 12'b111101111111;
   60816: result <= 12'b111101111111;
   60817: result <= 12'b111101111111;
   60818: result <= 12'b111101111111;
   60819: result <= 12'b111101111110;
   60820: result <= 12'b111101111110;
   60821: result <= 12'b111101111110;
   60822: result <= 12'b111101111110;
   60823: result <= 12'b111101111110;
   60824: result <= 12'b111101111110;
   60825: result <= 12'b111101111101;
   60826: result <= 12'b111101111101;
   60827: result <= 12'b111101111101;
   60828: result <= 12'b111101111101;
   60829: result <= 12'b111101111101;
   60830: result <= 12'b111101111100;
   60831: result <= 12'b111101111100;
   60832: result <= 12'b111101111100;
   60833: result <= 12'b111101111100;
   60834: result <= 12'b111101111100;
   60835: result <= 12'b111101111100;
   60836: result <= 12'b111101111011;
   60837: result <= 12'b111101111011;
   60838: result <= 12'b111101111011;
   60839: result <= 12'b111101111011;
   60840: result <= 12'b111101111011;
   60841: result <= 12'b111101111011;
   60842: result <= 12'b111101111010;
   60843: result <= 12'b111101111010;
   60844: result <= 12'b111101111010;
   60845: result <= 12'b111101111010;
   60846: result <= 12'b111101111010;
   60847: result <= 12'b111101111001;
   60848: result <= 12'b111101111001;
   60849: result <= 12'b111101111001;
   60850: result <= 12'b111101111001;
   60851: result <= 12'b111101111001;
   60852: result <= 12'b111101111001;
   60853: result <= 12'b111101111000;
   60854: result <= 12'b111101111000;
   60855: result <= 12'b111101111000;
   60856: result <= 12'b111101111000;
   60857: result <= 12'b111101111000;
   60858: result <= 12'b111101111000;
   60859: result <= 12'b111101110111;
   60860: result <= 12'b111101110111;
   60861: result <= 12'b111101110111;
   60862: result <= 12'b111101110111;
   60863: result <= 12'b111101110111;
   60864: result <= 12'b111101110110;
   60865: result <= 12'b111101110110;
   60866: result <= 12'b111101110110;
   60867: result <= 12'b111101110110;
   60868: result <= 12'b111101110110;
   60869: result <= 12'b111101110110;
   60870: result <= 12'b111101110101;
   60871: result <= 12'b111101110101;
   60872: result <= 12'b111101110101;
   60873: result <= 12'b111101110101;
   60874: result <= 12'b111101110101;
   60875: result <= 12'b111101110101;
   60876: result <= 12'b111101110100;
   60877: result <= 12'b111101110100;
   60878: result <= 12'b111101110100;
   60879: result <= 12'b111101110100;
   60880: result <= 12'b111101110100;
   60881: result <= 12'b111101110011;
   60882: result <= 12'b111101110011;
   60883: result <= 12'b111101110011;
   60884: result <= 12'b111101110011;
   60885: result <= 12'b111101110011;
   60886: result <= 12'b111101110011;
   60887: result <= 12'b111101110010;
   60888: result <= 12'b111101110010;
   60889: result <= 12'b111101110010;
   60890: result <= 12'b111101110010;
   60891: result <= 12'b111101110010;
   60892: result <= 12'b111101110010;
   60893: result <= 12'b111101110001;
   60894: result <= 12'b111101110001;
   60895: result <= 12'b111101110001;
   60896: result <= 12'b111101110001;
   60897: result <= 12'b111101110001;
   60898: result <= 12'b111101110000;
   60899: result <= 12'b111101110000;
   60900: result <= 12'b111101110000;
   60901: result <= 12'b111101110000;
   60902: result <= 12'b111101110000;
   60903: result <= 12'b111101110000;
   60904: result <= 12'b111101101111;
   60905: result <= 12'b111101101111;
   60906: result <= 12'b111101101111;
   60907: result <= 12'b111101101111;
   60908: result <= 12'b111101101111;
   60909: result <= 12'b111101101111;
   60910: result <= 12'b111101101110;
   60911: result <= 12'b111101101110;
   60912: result <= 12'b111101101110;
   60913: result <= 12'b111101101110;
   60914: result <= 12'b111101101110;
   60915: result <= 12'b111101101101;
   60916: result <= 12'b111101101101;
   60917: result <= 12'b111101101101;
   60918: result <= 12'b111101101101;
   60919: result <= 12'b111101101101;
   60920: result <= 12'b111101101101;
   60921: result <= 12'b111101101100;
   60922: result <= 12'b111101101100;
   60923: result <= 12'b111101101100;
   60924: result <= 12'b111101101100;
   60925: result <= 12'b111101101100;
   60926: result <= 12'b111101101011;
   60927: result <= 12'b111101101011;
   60928: result <= 12'b111101101011;
   60929: result <= 12'b111101101011;
   60930: result <= 12'b111101101011;
   60931: result <= 12'b111101101011;
   60932: result <= 12'b111101101010;
   60933: result <= 12'b111101101010;
   60934: result <= 12'b111101101010;
   60935: result <= 12'b111101101010;
   60936: result <= 12'b111101101010;
   60937: result <= 12'b111101101010;
   60938: result <= 12'b111101101001;
   60939: result <= 12'b111101101001;
   60940: result <= 12'b111101101001;
   60941: result <= 12'b111101101001;
   60942: result <= 12'b111101101001;
   60943: result <= 12'b111101101000;
   60944: result <= 12'b111101101000;
   60945: result <= 12'b111101101000;
   60946: result <= 12'b111101101000;
   60947: result <= 12'b111101101000;
   60948: result <= 12'b111101101000;
   60949: result <= 12'b111101100111;
   60950: result <= 12'b111101100111;
   60951: result <= 12'b111101100111;
   60952: result <= 12'b111101100111;
   60953: result <= 12'b111101100111;
   60954: result <= 12'b111101100111;
   60955: result <= 12'b111101100110;
   60956: result <= 12'b111101100110;
   60957: result <= 12'b111101100110;
   60958: result <= 12'b111101100110;
   60959: result <= 12'b111101100110;
   60960: result <= 12'b111101100101;
   60961: result <= 12'b111101100101;
   60962: result <= 12'b111101100101;
   60963: result <= 12'b111101100101;
   60964: result <= 12'b111101100101;
   60965: result <= 12'b111101100101;
   60966: result <= 12'b111101100100;
   60967: result <= 12'b111101100100;
   60968: result <= 12'b111101100100;
   60969: result <= 12'b111101100100;
   60970: result <= 12'b111101100100;
   60971: result <= 12'b111101100011;
   60972: result <= 12'b111101100011;
   60973: result <= 12'b111101100011;
   60974: result <= 12'b111101100011;
   60975: result <= 12'b111101100011;
   60976: result <= 12'b111101100011;
   60977: result <= 12'b111101100010;
   60978: result <= 12'b111101100010;
   60979: result <= 12'b111101100010;
   60980: result <= 12'b111101100010;
   60981: result <= 12'b111101100010;
   60982: result <= 12'b111101100010;
   60983: result <= 12'b111101100001;
   60984: result <= 12'b111101100001;
   60985: result <= 12'b111101100001;
   60986: result <= 12'b111101100001;
   60987: result <= 12'b111101100001;
   60988: result <= 12'b111101100000;
   60989: result <= 12'b111101100000;
   60990: result <= 12'b111101100000;
   60991: result <= 12'b111101100000;
   60992: result <= 12'b111101100000;
   60993: result <= 12'b111101100000;
   60994: result <= 12'b111101011111;
   60995: result <= 12'b111101011111;
   60996: result <= 12'b111101011111;
   60997: result <= 12'b111101011111;
   60998: result <= 12'b111101011111;
   60999: result <= 12'b111101011111;
   61000: result <= 12'b111101011110;
   61001: result <= 12'b111101011110;
   61002: result <= 12'b111101011110;
   61003: result <= 12'b111101011110;
   61004: result <= 12'b111101011110;
   61005: result <= 12'b111101011101;
   61006: result <= 12'b111101011101;
   61007: result <= 12'b111101011101;
   61008: result <= 12'b111101011101;
   61009: result <= 12'b111101011101;
   61010: result <= 12'b111101011101;
   61011: result <= 12'b111101011100;
   61012: result <= 12'b111101011100;
   61013: result <= 12'b111101011100;
   61014: result <= 12'b111101011100;
   61015: result <= 12'b111101011100;
   61016: result <= 12'b111101011011;
   61017: result <= 12'b111101011011;
   61018: result <= 12'b111101011011;
   61019: result <= 12'b111101011011;
   61020: result <= 12'b111101011011;
   61021: result <= 12'b111101011011;
   61022: result <= 12'b111101011010;
   61023: result <= 12'b111101011010;
   61024: result <= 12'b111101011010;
   61025: result <= 12'b111101011010;
   61026: result <= 12'b111101011010;
   61027: result <= 12'b111101011010;
   61028: result <= 12'b111101011001;
   61029: result <= 12'b111101011001;
   61030: result <= 12'b111101011001;
   61031: result <= 12'b111101011001;
   61032: result <= 12'b111101011001;
   61033: result <= 12'b111101011000;
   61034: result <= 12'b111101011000;
   61035: result <= 12'b111101011000;
   61036: result <= 12'b111101011000;
   61037: result <= 12'b111101011000;
   61038: result <= 12'b111101011000;
   61039: result <= 12'b111101010111;
   61040: result <= 12'b111101010111;
   61041: result <= 12'b111101010111;
   61042: result <= 12'b111101010111;
   61043: result <= 12'b111101010111;
   61044: result <= 12'b111101010110;
   61045: result <= 12'b111101010110;
   61046: result <= 12'b111101010110;
   61047: result <= 12'b111101010110;
   61048: result <= 12'b111101010110;
   61049: result <= 12'b111101010110;
   61050: result <= 12'b111101010101;
   61051: result <= 12'b111101010101;
   61052: result <= 12'b111101010101;
   61053: result <= 12'b111101010101;
   61054: result <= 12'b111101010101;
   61055: result <= 12'b111101010101;
   61056: result <= 12'b111101010100;
   61057: result <= 12'b111101010100;
   61058: result <= 12'b111101010100;
   61059: result <= 12'b111101010100;
   61060: result <= 12'b111101010100;
   61061: result <= 12'b111101010011;
   61062: result <= 12'b111101010011;
   61063: result <= 12'b111101010011;
   61064: result <= 12'b111101010011;
   61065: result <= 12'b111101010011;
   61066: result <= 12'b111101010011;
   61067: result <= 12'b111101010010;
   61068: result <= 12'b111101010010;
   61069: result <= 12'b111101010010;
   61070: result <= 12'b111101010010;
   61071: result <= 12'b111101010010;
   61072: result <= 12'b111101010001;
   61073: result <= 12'b111101010001;
   61074: result <= 12'b111101010001;
   61075: result <= 12'b111101010001;
   61076: result <= 12'b111101010001;
   61077: result <= 12'b111101010001;
   61078: result <= 12'b111101010000;
   61079: result <= 12'b111101010000;
   61080: result <= 12'b111101010000;
   61081: result <= 12'b111101010000;
   61082: result <= 12'b111101010000;
   61083: result <= 12'b111101010000;
   61084: result <= 12'b111101001111;
   61085: result <= 12'b111101001111;
   61086: result <= 12'b111101001111;
   61087: result <= 12'b111101001111;
   61088: result <= 12'b111101001111;
   61089: result <= 12'b111101001110;
   61090: result <= 12'b111101001110;
   61091: result <= 12'b111101001110;
   61092: result <= 12'b111101001110;
   61093: result <= 12'b111101001110;
   61094: result <= 12'b111101001110;
   61095: result <= 12'b111101001101;
   61096: result <= 12'b111101001101;
   61097: result <= 12'b111101001101;
   61098: result <= 12'b111101001101;
   61099: result <= 12'b111101001101;
   61100: result <= 12'b111101001100;
   61101: result <= 12'b111101001100;
   61102: result <= 12'b111101001100;
   61103: result <= 12'b111101001100;
   61104: result <= 12'b111101001100;
   61105: result <= 12'b111101001100;
   61106: result <= 12'b111101001011;
   61107: result <= 12'b111101001011;
   61108: result <= 12'b111101001011;
   61109: result <= 12'b111101001011;
   61110: result <= 12'b111101001011;
   61111: result <= 12'b111101001011;
   61112: result <= 12'b111101001010;
   61113: result <= 12'b111101001010;
   61114: result <= 12'b111101001010;
   61115: result <= 12'b111101001010;
   61116: result <= 12'b111101001010;
   61117: result <= 12'b111101001001;
   61118: result <= 12'b111101001001;
   61119: result <= 12'b111101001001;
   61120: result <= 12'b111101001001;
   61121: result <= 12'b111101001001;
   61122: result <= 12'b111101001001;
   61123: result <= 12'b111101001000;
   61124: result <= 12'b111101001000;
   61125: result <= 12'b111101001000;
   61126: result <= 12'b111101001000;
   61127: result <= 12'b111101001000;
   61128: result <= 12'b111101000111;
   61129: result <= 12'b111101000111;
   61130: result <= 12'b111101000111;
   61131: result <= 12'b111101000111;
   61132: result <= 12'b111101000111;
   61133: result <= 12'b111101000111;
   61134: result <= 12'b111101000110;
   61135: result <= 12'b111101000110;
   61136: result <= 12'b111101000110;
   61137: result <= 12'b111101000110;
   61138: result <= 12'b111101000110;
   61139: result <= 12'b111101000110;
   61140: result <= 12'b111101000101;
   61141: result <= 12'b111101000101;
   61142: result <= 12'b111101000101;
   61143: result <= 12'b111101000101;
   61144: result <= 12'b111101000101;
   61145: result <= 12'b111101000100;
   61146: result <= 12'b111101000100;
   61147: result <= 12'b111101000100;
   61148: result <= 12'b111101000100;
   61149: result <= 12'b111101000100;
   61150: result <= 12'b111101000100;
   61151: result <= 12'b111101000011;
   61152: result <= 12'b111101000011;
   61153: result <= 12'b111101000011;
   61154: result <= 12'b111101000011;
   61155: result <= 12'b111101000011;
   61156: result <= 12'b111101000010;
   61157: result <= 12'b111101000010;
   61158: result <= 12'b111101000010;
   61159: result <= 12'b111101000010;
   61160: result <= 12'b111101000010;
   61161: result <= 12'b111101000010;
   61162: result <= 12'b111101000001;
   61163: result <= 12'b111101000001;
   61164: result <= 12'b111101000001;
   61165: result <= 12'b111101000001;
   61166: result <= 12'b111101000001;
   61167: result <= 12'b111101000000;
   61168: result <= 12'b111101000000;
   61169: result <= 12'b111101000000;
   61170: result <= 12'b111101000000;
   61171: result <= 12'b111101000000;
   61172: result <= 12'b111101000000;
   61173: result <= 12'b111100111111;
   61174: result <= 12'b111100111111;
   61175: result <= 12'b111100111111;
   61176: result <= 12'b111100111111;
   61177: result <= 12'b111100111111;
   61178: result <= 12'b111100111111;
   61179: result <= 12'b111100111110;
   61180: result <= 12'b111100111110;
   61181: result <= 12'b111100111110;
   61182: result <= 12'b111100111110;
   61183: result <= 12'b111100111110;
   61184: result <= 12'b111100111101;
   61185: result <= 12'b111100111101;
   61186: result <= 12'b111100111101;
   61187: result <= 12'b111100111101;
   61188: result <= 12'b111100111101;
   61189: result <= 12'b111100111101;
   61190: result <= 12'b111100111100;
   61191: result <= 12'b111100111100;
   61192: result <= 12'b111100111100;
   61193: result <= 12'b111100111100;
   61194: result <= 12'b111100111100;
   61195: result <= 12'b111100111011;
   61196: result <= 12'b111100111011;
   61197: result <= 12'b111100111011;
   61198: result <= 12'b111100111011;
   61199: result <= 12'b111100111011;
   61200: result <= 12'b111100111011;
   61201: result <= 12'b111100111010;
   61202: result <= 12'b111100111010;
   61203: result <= 12'b111100111010;
   61204: result <= 12'b111100111010;
   61205: result <= 12'b111100111010;
   61206: result <= 12'b111100111001;
   61207: result <= 12'b111100111001;
   61208: result <= 12'b111100111001;
   61209: result <= 12'b111100111001;
   61210: result <= 12'b111100111001;
   61211: result <= 12'b111100111001;
   61212: result <= 12'b111100111000;
   61213: result <= 12'b111100111000;
   61214: result <= 12'b111100111000;
   61215: result <= 12'b111100111000;
   61216: result <= 12'b111100111000;
   61217: result <= 12'b111100111000;
   61218: result <= 12'b111100110111;
   61219: result <= 12'b111100110111;
   61220: result <= 12'b111100110111;
   61221: result <= 12'b111100110111;
   61222: result <= 12'b111100110111;
   61223: result <= 12'b111100110110;
   61224: result <= 12'b111100110110;
   61225: result <= 12'b111100110110;
   61226: result <= 12'b111100110110;
   61227: result <= 12'b111100110110;
   61228: result <= 12'b111100110110;
   61229: result <= 12'b111100110101;
   61230: result <= 12'b111100110101;
   61231: result <= 12'b111100110101;
   61232: result <= 12'b111100110101;
   61233: result <= 12'b111100110101;
   61234: result <= 12'b111100110100;
   61235: result <= 12'b111100110100;
   61236: result <= 12'b111100110100;
   61237: result <= 12'b111100110100;
   61238: result <= 12'b111100110100;
   61239: result <= 12'b111100110100;
   61240: result <= 12'b111100110011;
   61241: result <= 12'b111100110011;
   61242: result <= 12'b111100110011;
   61243: result <= 12'b111100110011;
   61244: result <= 12'b111100110011;
   61245: result <= 12'b111100110010;
   61246: result <= 12'b111100110010;
   61247: result <= 12'b111100110010;
   61248: result <= 12'b111100110010;
   61249: result <= 12'b111100110010;
   61250: result <= 12'b111100110010;
   61251: result <= 12'b111100110001;
   61252: result <= 12'b111100110001;
   61253: result <= 12'b111100110001;
   61254: result <= 12'b111100110001;
   61255: result <= 12'b111100110001;
   61256: result <= 12'b111100110000;
   61257: result <= 12'b111100110000;
   61258: result <= 12'b111100110000;
   61259: result <= 12'b111100110000;
   61260: result <= 12'b111100110000;
   61261: result <= 12'b111100110000;
   61262: result <= 12'b111100101111;
   61263: result <= 12'b111100101111;
   61264: result <= 12'b111100101111;
   61265: result <= 12'b111100101111;
   61266: result <= 12'b111100101111;
   61267: result <= 12'b111100101111;
   61268: result <= 12'b111100101110;
   61269: result <= 12'b111100101110;
   61270: result <= 12'b111100101110;
   61271: result <= 12'b111100101110;
   61272: result <= 12'b111100101110;
   61273: result <= 12'b111100101101;
   61274: result <= 12'b111100101101;
   61275: result <= 12'b111100101101;
   61276: result <= 12'b111100101101;
   61277: result <= 12'b111100101101;
   61278: result <= 12'b111100101101;
   61279: result <= 12'b111100101100;
   61280: result <= 12'b111100101100;
   61281: result <= 12'b111100101100;
   61282: result <= 12'b111100101100;
   61283: result <= 12'b111100101100;
   61284: result <= 12'b111100101011;
   61285: result <= 12'b111100101011;
   61286: result <= 12'b111100101011;
   61287: result <= 12'b111100101011;
   61288: result <= 12'b111100101011;
   61289: result <= 12'b111100101011;
   61290: result <= 12'b111100101010;
   61291: result <= 12'b111100101010;
   61292: result <= 12'b111100101010;
   61293: result <= 12'b111100101010;
   61294: result <= 12'b111100101010;
   61295: result <= 12'b111100101001;
   61296: result <= 12'b111100101001;
   61297: result <= 12'b111100101001;
   61298: result <= 12'b111100101001;
   61299: result <= 12'b111100101001;
   61300: result <= 12'b111100101001;
   61301: result <= 12'b111100101000;
   61302: result <= 12'b111100101000;
   61303: result <= 12'b111100101000;
   61304: result <= 12'b111100101000;
   61305: result <= 12'b111100101000;
   61306: result <= 12'b111100100111;
   61307: result <= 12'b111100100111;
   61308: result <= 12'b111100100111;
   61309: result <= 12'b111100100111;
   61310: result <= 12'b111100100111;
   61311: result <= 12'b111100100111;
   61312: result <= 12'b111100100110;
   61313: result <= 12'b111100100110;
   61314: result <= 12'b111100100110;
   61315: result <= 12'b111100100110;
   61316: result <= 12'b111100100110;
   61317: result <= 12'b111100100101;
   61318: result <= 12'b111100100101;
   61319: result <= 12'b111100100101;
   61320: result <= 12'b111100100101;
   61321: result <= 12'b111100100101;
   61322: result <= 12'b111100100101;
   61323: result <= 12'b111100100100;
   61324: result <= 12'b111100100100;
   61325: result <= 12'b111100100100;
   61326: result <= 12'b111100100100;
   61327: result <= 12'b111100100100;
   61328: result <= 12'b111100100100;
   61329: result <= 12'b111100100011;
   61330: result <= 12'b111100100011;
   61331: result <= 12'b111100100011;
   61332: result <= 12'b111100100011;
   61333: result <= 12'b111100100011;
   61334: result <= 12'b111100100010;
   61335: result <= 12'b111100100010;
   61336: result <= 12'b111100100010;
   61337: result <= 12'b111100100010;
   61338: result <= 12'b111100100010;
   61339: result <= 12'b111100100010;
   61340: result <= 12'b111100100001;
   61341: result <= 12'b111100100001;
   61342: result <= 12'b111100100001;
   61343: result <= 12'b111100100001;
   61344: result <= 12'b111100100001;
   61345: result <= 12'b111100100000;
   61346: result <= 12'b111100100000;
   61347: result <= 12'b111100100000;
   61348: result <= 12'b111100100000;
   61349: result <= 12'b111100100000;
   61350: result <= 12'b111100100000;
   61351: result <= 12'b111100011111;
   61352: result <= 12'b111100011111;
   61353: result <= 12'b111100011111;
   61354: result <= 12'b111100011111;
   61355: result <= 12'b111100011111;
   61356: result <= 12'b111100011110;
   61357: result <= 12'b111100011110;
   61358: result <= 12'b111100011110;
   61359: result <= 12'b111100011110;
   61360: result <= 12'b111100011110;
   61361: result <= 12'b111100011110;
   61362: result <= 12'b111100011101;
   61363: result <= 12'b111100011101;
   61364: result <= 12'b111100011101;
   61365: result <= 12'b111100011101;
   61366: result <= 12'b111100011101;
   61367: result <= 12'b111100011100;
   61368: result <= 12'b111100011100;
   61369: result <= 12'b111100011100;
   61370: result <= 12'b111100011100;
   61371: result <= 12'b111100011100;
   61372: result <= 12'b111100011100;
   61373: result <= 12'b111100011011;
   61374: result <= 12'b111100011011;
   61375: result <= 12'b111100011011;
   61376: result <= 12'b111100011011;
   61377: result <= 12'b111100011011;
   61378: result <= 12'b111100011010;
   61379: result <= 12'b111100011010;
   61380: result <= 12'b111100011010;
   61381: result <= 12'b111100011010;
   61382: result <= 12'b111100011010;
   61383: result <= 12'b111100011010;
   61384: result <= 12'b111100011001;
   61385: result <= 12'b111100011001;
   61386: result <= 12'b111100011001;
   61387: result <= 12'b111100011001;
   61388: result <= 12'b111100011001;
   61389: result <= 12'b111100011000;
   61390: result <= 12'b111100011000;
   61391: result <= 12'b111100011000;
   61392: result <= 12'b111100011000;
   61393: result <= 12'b111100011000;
   61394: result <= 12'b111100011000;
   61395: result <= 12'b111100010111;
   61396: result <= 12'b111100010111;
   61397: result <= 12'b111100010111;
   61398: result <= 12'b111100010111;
   61399: result <= 12'b111100010111;
   61400: result <= 12'b111100010110;
   61401: result <= 12'b111100010110;
   61402: result <= 12'b111100010110;
   61403: result <= 12'b111100010110;
   61404: result <= 12'b111100010110;
   61405: result <= 12'b111100010110;
   61406: result <= 12'b111100010101;
   61407: result <= 12'b111100010101;
   61408: result <= 12'b111100010101;
   61409: result <= 12'b111100010101;
   61410: result <= 12'b111100010101;
   61411: result <= 12'b111100010100;
   61412: result <= 12'b111100010100;
   61413: result <= 12'b111100010100;
   61414: result <= 12'b111100010100;
   61415: result <= 12'b111100010100;
   61416: result <= 12'b111100010100;
   61417: result <= 12'b111100010011;
   61418: result <= 12'b111100010011;
   61419: result <= 12'b111100010011;
   61420: result <= 12'b111100010011;
   61421: result <= 12'b111100010011;
   61422: result <= 12'b111100010010;
   61423: result <= 12'b111100010010;
   61424: result <= 12'b111100010010;
   61425: result <= 12'b111100010010;
   61426: result <= 12'b111100010010;
   61427: result <= 12'b111100010010;
   61428: result <= 12'b111100010001;
   61429: result <= 12'b111100010001;
   61430: result <= 12'b111100010001;
   61431: result <= 12'b111100010001;
   61432: result <= 12'b111100010001;
   61433: result <= 12'b111100010001;
   61434: result <= 12'b111100010000;
   61435: result <= 12'b111100010000;
   61436: result <= 12'b111100010000;
   61437: result <= 12'b111100010000;
   61438: result <= 12'b111100010000;
   61439: result <= 12'b111100001111;
   61440: result <= 12'b111100001111;
   61441: result <= 12'b111100001111;
   61442: result <= 12'b111100001111;
   61443: result <= 12'b111100001111;
   61444: result <= 12'b111100001111;
   61445: result <= 12'b111100001110;
   61446: result <= 12'b111100001110;
   61447: result <= 12'b111100001110;
   61448: result <= 12'b111100001110;
   61449: result <= 12'b111100001110;
   61450: result <= 12'b111100001101;
   61451: result <= 12'b111100001101;
   61452: result <= 12'b111100001101;
   61453: result <= 12'b111100001101;
   61454: result <= 12'b111100001101;
   61455: result <= 12'b111100001101;
   61456: result <= 12'b111100001100;
   61457: result <= 12'b111100001100;
   61458: result <= 12'b111100001100;
   61459: result <= 12'b111100001100;
   61460: result <= 12'b111100001100;
   61461: result <= 12'b111100001011;
   61462: result <= 12'b111100001011;
   61463: result <= 12'b111100001011;
   61464: result <= 12'b111100001011;
   61465: result <= 12'b111100001011;
   61466: result <= 12'b111100001011;
   61467: result <= 12'b111100001010;
   61468: result <= 12'b111100001010;
   61469: result <= 12'b111100001010;
   61470: result <= 12'b111100001010;
   61471: result <= 12'b111100001010;
   61472: result <= 12'b111100001001;
   61473: result <= 12'b111100001001;
   61474: result <= 12'b111100001001;
   61475: result <= 12'b111100001001;
   61476: result <= 12'b111100001001;
   61477: result <= 12'b111100001001;
   61478: result <= 12'b111100001000;
   61479: result <= 12'b111100001000;
   61480: result <= 12'b111100001000;
   61481: result <= 12'b111100001000;
   61482: result <= 12'b111100001000;
   61483: result <= 12'b111100000111;
   61484: result <= 12'b111100000111;
   61485: result <= 12'b111100000111;
   61486: result <= 12'b111100000111;
   61487: result <= 12'b111100000111;
   61488: result <= 12'b111100000111;
   61489: result <= 12'b111100000110;
   61490: result <= 12'b111100000110;
   61491: result <= 12'b111100000110;
   61492: result <= 12'b111100000110;
   61493: result <= 12'b111100000110;
   61494: result <= 12'b111100000101;
   61495: result <= 12'b111100000101;
   61496: result <= 12'b111100000101;
   61497: result <= 12'b111100000101;
   61498: result <= 12'b111100000101;
   61499: result <= 12'b111100000101;
   61500: result <= 12'b111100000100;
   61501: result <= 12'b111100000100;
   61502: result <= 12'b111100000100;
   61503: result <= 12'b111100000100;
   61504: result <= 12'b111100000100;
   61505: result <= 12'b111100000011;
   61506: result <= 12'b111100000011;
   61507: result <= 12'b111100000011;
   61508: result <= 12'b111100000011;
   61509: result <= 12'b111100000011;
   61510: result <= 12'b111100000011;
   61511: result <= 12'b111100000010;
   61512: result <= 12'b111100000010;
   61513: result <= 12'b111100000010;
   61514: result <= 12'b111100000010;
   61515: result <= 12'b111100000010;
   61516: result <= 12'b111100000001;
   61517: result <= 12'b111100000001;
   61518: result <= 12'b111100000001;
   61519: result <= 12'b111100000001;
   61520: result <= 12'b111100000001;
   61521: result <= 12'b111100000001;
   61522: result <= 12'b111100000000;
   61523: result <= 12'b111100000000;
   61524: result <= 12'b111100000000;
   61525: result <= 12'b111100000000;
   61526: result <= 12'b111100000000;
   61527: result <= 12'b111011111111;
   61528: result <= 12'b111011111111;
   61529: result <= 12'b111011111111;
   61530: result <= 12'b111011111111;
   61531: result <= 12'b111011111111;
   61532: result <= 12'b111011111111;
   61533: result <= 12'b111011111110;
   61534: result <= 12'b111011111110;
   61535: result <= 12'b111011111110;
   61536: result <= 12'b111011111110;
   61537: result <= 12'b111011111110;
   61538: result <= 12'b111011111101;
   61539: result <= 12'b111011111101;
   61540: result <= 12'b111011111101;
   61541: result <= 12'b111011111101;
   61542: result <= 12'b111011111101;
   61543: result <= 12'b111011111101;
   61544: result <= 12'b111011111100;
   61545: result <= 12'b111011111100;
   61546: result <= 12'b111011111100;
   61547: result <= 12'b111011111100;
   61548: result <= 12'b111011111100;
   61549: result <= 12'b111011111011;
   61550: result <= 12'b111011111011;
   61551: result <= 12'b111011111011;
   61552: result <= 12'b111011111011;
   61553: result <= 12'b111011111011;
   61554: result <= 12'b111011111011;
   61555: result <= 12'b111011111010;
   61556: result <= 12'b111011111010;
   61557: result <= 12'b111011111010;
   61558: result <= 12'b111011111010;
   61559: result <= 12'b111011111010;
   61560: result <= 12'b111011111001;
   61561: result <= 12'b111011111001;
   61562: result <= 12'b111011111001;
   61563: result <= 12'b111011111001;
   61564: result <= 12'b111011111001;
   61565: result <= 12'b111011111001;
   61566: result <= 12'b111011111000;
   61567: result <= 12'b111011111000;
   61568: result <= 12'b111011111000;
   61569: result <= 12'b111011111000;
   61570: result <= 12'b111011111000;
   61571: result <= 12'b111011110111;
   61572: result <= 12'b111011110111;
   61573: result <= 12'b111011110111;
   61574: result <= 12'b111011110111;
   61575: result <= 12'b111011110111;
   61576: result <= 12'b111011110110;
   61577: result <= 12'b111011110110;
   61578: result <= 12'b111011110110;
   61579: result <= 12'b111011110110;
   61580: result <= 12'b111011110110;
   61581: result <= 12'b111011110110;
   61582: result <= 12'b111011110101;
   61583: result <= 12'b111011110101;
   61584: result <= 12'b111011110101;
   61585: result <= 12'b111011110101;
   61586: result <= 12'b111011110101;
   61587: result <= 12'b111011110100;
   61588: result <= 12'b111011110100;
   61589: result <= 12'b111011110100;
   61590: result <= 12'b111011110100;
   61591: result <= 12'b111011110100;
   61592: result <= 12'b111011110100;
   61593: result <= 12'b111011110011;
   61594: result <= 12'b111011110011;
   61595: result <= 12'b111011110011;
   61596: result <= 12'b111011110011;
   61597: result <= 12'b111011110011;
   61598: result <= 12'b111011110010;
   61599: result <= 12'b111011110010;
   61600: result <= 12'b111011110010;
   61601: result <= 12'b111011110010;
   61602: result <= 12'b111011110010;
   61603: result <= 12'b111011110010;
   61604: result <= 12'b111011110001;
   61605: result <= 12'b111011110001;
   61606: result <= 12'b111011110001;
   61607: result <= 12'b111011110001;
   61608: result <= 12'b111011110001;
   61609: result <= 12'b111011110000;
   61610: result <= 12'b111011110000;
   61611: result <= 12'b111011110000;
   61612: result <= 12'b111011110000;
   61613: result <= 12'b111011110000;
   61614: result <= 12'b111011110000;
   61615: result <= 12'b111011101111;
   61616: result <= 12'b111011101111;
   61617: result <= 12'b111011101111;
   61618: result <= 12'b111011101111;
   61619: result <= 12'b111011101111;
   61620: result <= 12'b111011101110;
   61621: result <= 12'b111011101110;
   61622: result <= 12'b111011101110;
   61623: result <= 12'b111011101110;
   61624: result <= 12'b111011101110;
   61625: result <= 12'b111011101110;
   61626: result <= 12'b111011101101;
   61627: result <= 12'b111011101101;
   61628: result <= 12'b111011101101;
   61629: result <= 12'b111011101101;
   61630: result <= 12'b111011101101;
   61631: result <= 12'b111011101100;
   61632: result <= 12'b111011101100;
   61633: result <= 12'b111011101100;
   61634: result <= 12'b111011101100;
   61635: result <= 12'b111011101100;
   61636: result <= 12'b111011101100;
   61637: result <= 12'b111011101011;
   61638: result <= 12'b111011101011;
   61639: result <= 12'b111011101011;
   61640: result <= 12'b111011101011;
   61641: result <= 12'b111011101011;
   61642: result <= 12'b111011101010;
   61643: result <= 12'b111011101010;
   61644: result <= 12'b111011101010;
   61645: result <= 12'b111011101010;
   61646: result <= 12'b111011101010;
   61647: result <= 12'b111011101010;
   61648: result <= 12'b111011101001;
   61649: result <= 12'b111011101001;
   61650: result <= 12'b111011101001;
   61651: result <= 12'b111011101001;
   61652: result <= 12'b111011101001;
   61653: result <= 12'b111011101000;
   61654: result <= 12'b111011101000;
   61655: result <= 12'b111011101000;
   61656: result <= 12'b111011101000;
   61657: result <= 12'b111011101000;
   61658: result <= 12'b111011101000;
   61659: result <= 12'b111011100111;
   61660: result <= 12'b111011100111;
   61661: result <= 12'b111011100111;
   61662: result <= 12'b111011100111;
   61663: result <= 12'b111011100111;
   61664: result <= 12'b111011100110;
   61665: result <= 12'b111011100110;
   61666: result <= 12'b111011100110;
   61667: result <= 12'b111011100110;
   61668: result <= 12'b111011100110;
   61669: result <= 12'b111011100110;
   61670: result <= 12'b111011100101;
   61671: result <= 12'b111011100101;
   61672: result <= 12'b111011100101;
   61673: result <= 12'b111011100101;
   61674: result <= 12'b111011100101;
   61675: result <= 12'b111011100100;
   61676: result <= 12'b111011100100;
   61677: result <= 12'b111011100100;
   61678: result <= 12'b111011100100;
   61679: result <= 12'b111011100100;
   61680: result <= 12'b111011100011;
   61681: result <= 12'b111011100011;
   61682: result <= 12'b111011100011;
   61683: result <= 12'b111011100011;
   61684: result <= 12'b111011100011;
   61685: result <= 12'b111011100011;
   61686: result <= 12'b111011100010;
   61687: result <= 12'b111011100010;
   61688: result <= 12'b111011100010;
   61689: result <= 12'b111011100010;
   61690: result <= 12'b111011100010;
   61691: result <= 12'b111011100001;
   61692: result <= 12'b111011100001;
   61693: result <= 12'b111011100001;
   61694: result <= 12'b111011100001;
   61695: result <= 12'b111011100001;
   61696: result <= 12'b111011100001;
   61697: result <= 12'b111011100000;
   61698: result <= 12'b111011100000;
   61699: result <= 12'b111011100000;
   61700: result <= 12'b111011100000;
   61701: result <= 12'b111011100000;
   61702: result <= 12'b111011011111;
   61703: result <= 12'b111011011111;
   61704: result <= 12'b111011011111;
   61705: result <= 12'b111011011111;
   61706: result <= 12'b111011011111;
   61707: result <= 12'b111011011111;
   61708: result <= 12'b111011011110;
   61709: result <= 12'b111011011110;
   61710: result <= 12'b111011011110;
   61711: result <= 12'b111011011110;
   61712: result <= 12'b111011011110;
   61713: result <= 12'b111011011101;
   61714: result <= 12'b111011011101;
   61715: result <= 12'b111011011101;
   61716: result <= 12'b111011011101;
   61717: result <= 12'b111011011101;
   61718: result <= 12'b111011011101;
   61719: result <= 12'b111011011100;
   61720: result <= 12'b111011011100;
   61721: result <= 12'b111011011100;
   61722: result <= 12'b111011011100;
   61723: result <= 12'b111011011100;
   61724: result <= 12'b111011011011;
   61725: result <= 12'b111011011011;
   61726: result <= 12'b111011011011;
   61727: result <= 12'b111011011011;
   61728: result <= 12'b111011011011;
   61729: result <= 12'b111011011011;
   61730: result <= 12'b111011011010;
   61731: result <= 12'b111011011010;
   61732: result <= 12'b111011011010;
   61733: result <= 12'b111011011010;
   61734: result <= 12'b111011011010;
   61735: result <= 12'b111011011001;
   61736: result <= 12'b111011011001;
   61737: result <= 12'b111011011001;
   61738: result <= 12'b111011011001;
   61739: result <= 12'b111011011001;
   61740: result <= 12'b111011011000;
   61741: result <= 12'b111011011000;
   61742: result <= 12'b111011011000;
   61743: result <= 12'b111011011000;
   61744: result <= 12'b111011011000;
   61745: result <= 12'b111011011000;
   61746: result <= 12'b111011010111;
   61747: result <= 12'b111011010111;
   61748: result <= 12'b111011010111;
   61749: result <= 12'b111011010111;
   61750: result <= 12'b111011010111;
   61751: result <= 12'b111011010110;
   61752: result <= 12'b111011010110;
   61753: result <= 12'b111011010110;
   61754: result <= 12'b111011010110;
   61755: result <= 12'b111011010110;
   61756: result <= 12'b111011010110;
   61757: result <= 12'b111011010101;
   61758: result <= 12'b111011010101;
   61759: result <= 12'b111011010101;
   61760: result <= 12'b111011010101;
   61761: result <= 12'b111011010101;
   61762: result <= 12'b111011010100;
   61763: result <= 12'b111011010100;
   61764: result <= 12'b111011010100;
   61765: result <= 12'b111011010100;
   61766: result <= 12'b111011010100;
   61767: result <= 12'b111011010100;
   61768: result <= 12'b111011010011;
   61769: result <= 12'b111011010011;
   61770: result <= 12'b111011010011;
   61771: result <= 12'b111011010011;
   61772: result <= 12'b111011010011;
   61773: result <= 12'b111011010010;
   61774: result <= 12'b111011010010;
   61775: result <= 12'b111011010010;
   61776: result <= 12'b111011010010;
   61777: result <= 12'b111011010010;
   61778: result <= 12'b111011010010;
   61779: result <= 12'b111011010001;
   61780: result <= 12'b111011010001;
   61781: result <= 12'b111011010001;
   61782: result <= 12'b111011010001;
   61783: result <= 12'b111011010001;
   61784: result <= 12'b111011010000;
   61785: result <= 12'b111011010000;
   61786: result <= 12'b111011010000;
   61787: result <= 12'b111011010000;
   61788: result <= 12'b111011010000;
   61789: result <= 12'b111011001111;
   61790: result <= 12'b111011001111;
   61791: result <= 12'b111011001111;
   61792: result <= 12'b111011001111;
   61793: result <= 12'b111011001111;
   61794: result <= 12'b111011001111;
   61795: result <= 12'b111011001110;
   61796: result <= 12'b111011001110;
   61797: result <= 12'b111011001110;
   61798: result <= 12'b111011001110;
   61799: result <= 12'b111011001110;
   61800: result <= 12'b111011001101;
   61801: result <= 12'b111011001101;
   61802: result <= 12'b111011001101;
   61803: result <= 12'b111011001101;
   61804: result <= 12'b111011001101;
   61805: result <= 12'b111011001101;
   61806: result <= 12'b111011001100;
   61807: result <= 12'b111011001100;
   61808: result <= 12'b111011001100;
   61809: result <= 12'b111011001100;
   61810: result <= 12'b111011001100;
   61811: result <= 12'b111011001011;
   61812: result <= 12'b111011001011;
   61813: result <= 12'b111011001011;
   61814: result <= 12'b111011001011;
   61815: result <= 12'b111011001011;
   61816: result <= 12'b111011001011;
   61817: result <= 12'b111011001010;
   61818: result <= 12'b111011001010;
   61819: result <= 12'b111011001010;
   61820: result <= 12'b111011001010;
   61821: result <= 12'b111011001010;
   61822: result <= 12'b111011001001;
   61823: result <= 12'b111011001001;
   61824: result <= 12'b111011001001;
   61825: result <= 12'b111011001001;
   61826: result <= 12'b111011001001;
   61827: result <= 12'b111011001001;
   61828: result <= 12'b111011001000;
   61829: result <= 12'b111011001000;
   61830: result <= 12'b111011001000;
   61831: result <= 12'b111011001000;
   61832: result <= 12'b111011001000;
   61833: result <= 12'b111011000111;
   61834: result <= 12'b111011000111;
   61835: result <= 12'b111011000111;
   61836: result <= 12'b111011000111;
   61837: result <= 12'b111011000111;
   61838: result <= 12'b111011000110;
   61839: result <= 12'b111011000110;
   61840: result <= 12'b111011000110;
   61841: result <= 12'b111011000110;
   61842: result <= 12'b111011000110;
   61843: result <= 12'b111011000110;
   61844: result <= 12'b111011000101;
   61845: result <= 12'b111011000101;
   61846: result <= 12'b111011000101;
   61847: result <= 12'b111011000101;
   61848: result <= 12'b111011000101;
   61849: result <= 12'b111011000100;
   61850: result <= 12'b111011000100;
   61851: result <= 12'b111011000100;
   61852: result <= 12'b111011000100;
   61853: result <= 12'b111011000100;
   61854: result <= 12'b111011000100;
   61855: result <= 12'b111011000011;
   61856: result <= 12'b111011000011;
   61857: result <= 12'b111011000011;
   61858: result <= 12'b111011000011;
   61859: result <= 12'b111011000011;
   61860: result <= 12'b111011000010;
   61861: result <= 12'b111011000010;
   61862: result <= 12'b111011000010;
   61863: result <= 12'b111011000010;
   61864: result <= 12'b111011000010;
   61865: result <= 12'b111011000010;
   61866: result <= 12'b111011000001;
   61867: result <= 12'b111011000001;
   61868: result <= 12'b111011000001;
   61869: result <= 12'b111011000001;
   61870: result <= 12'b111011000001;
   61871: result <= 12'b111011000000;
   61872: result <= 12'b111011000000;
   61873: result <= 12'b111011000000;
   61874: result <= 12'b111011000000;
   61875: result <= 12'b111011000000;
   61876: result <= 12'b111010111111;
   61877: result <= 12'b111010111111;
   61878: result <= 12'b111010111111;
   61879: result <= 12'b111010111111;
   61880: result <= 12'b111010111111;
   61881: result <= 12'b111010111111;
   61882: result <= 12'b111010111110;
   61883: result <= 12'b111010111110;
   61884: result <= 12'b111010111110;
   61885: result <= 12'b111010111110;
   61886: result <= 12'b111010111110;
   61887: result <= 12'b111010111101;
   61888: result <= 12'b111010111101;
   61889: result <= 12'b111010111101;
   61890: result <= 12'b111010111101;
   61891: result <= 12'b111010111101;
   61892: result <= 12'b111010111101;
   61893: result <= 12'b111010111100;
   61894: result <= 12'b111010111100;
   61895: result <= 12'b111010111100;
   61896: result <= 12'b111010111100;
   61897: result <= 12'b111010111100;
   61898: result <= 12'b111010111011;
   61899: result <= 12'b111010111011;
   61900: result <= 12'b111010111011;
   61901: result <= 12'b111010111011;
   61902: result <= 12'b111010111011;
   61903: result <= 12'b111010111011;
   61904: result <= 12'b111010111010;
   61905: result <= 12'b111010111010;
   61906: result <= 12'b111010111010;
   61907: result <= 12'b111010111010;
   61908: result <= 12'b111010111010;
   61909: result <= 12'b111010111001;
   61910: result <= 12'b111010111001;
   61911: result <= 12'b111010111001;
   61912: result <= 12'b111010111001;
   61913: result <= 12'b111010111001;
   61914: result <= 12'b111010111000;
   61915: result <= 12'b111010111000;
   61916: result <= 12'b111010111000;
   61917: result <= 12'b111010111000;
   61918: result <= 12'b111010111000;
   61919: result <= 12'b111010111000;
   61920: result <= 12'b111010110111;
   61921: result <= 12'b111010110111;
   61922: result <= 12'b111010110111;
   61923: result <= 12'b111010110111;
   61924: result <= 12'b111010110111;
   61925: result <= 12'b111010110110;
   61926: result <= 12'b111010110110;
   61927: result <= 12'b111010110110;
   61928: result <= 12'b111010110110;
   61929: result <= 12'b111010110110;
   61930: result <= 12'b111010110110;
   61931: result <= 12'b111010110101;
   61932: result <= 12'b111010110101;
   61933: result <= 12'b111010110101;
   61934: result <= 12'b111010110101;
   61935: result <= 12'b111010110101;
   61936: result <= 12'b111010110100;
   61937: result <= 12'b111010110100;
   61938: result <= 12'b111010110100;
   61939: result <= 12'b111010110100;
   61940: result <= 12'b111010110100;
   61941: result <= 12'b111010110011;
   61942: result <= 12'b111010110011;
   61943: result <= 12'b111010110011;
   61944: result <= 12'b111010110011;
   61945: result <= 12'b111010110011;
   61946: result <= 12'b111010110011;
   61947: result <= 12'b111010110010;
   61948: result <= 12'b111010110010;
   61949: result <= 12'b111010110010;
   61950: result <= 12'b111010110010;
   61951: result <= 12'b111010110010;
   61952: result <= 12'b111010110001;
   61953: result <= 12'b111010110001;
   61954: result <= 12'b111010110001;
   61955: result <= 12'b111010110001;
   61956: result <= 12'b111010110001;
   61957: result <= 12'b111010110001;
   61958: result <= 12'b111010110000;
   61959: result <= 12'b111010110000;
   61960: result <= 12'b111010110000;
   61961: result <= 12'b111010110000;
   61962: result <= 12'b111010110000;
   61963: result <= 12'b111010101111;
   61964: result <= 12'b111010101111;
   61965: result <= 12'b111010101111;
   61966: result <= 12'b111010101111;
   61967: result <= 12'b111010101111;
   61968: result <= 12'b111010101110;
   61969: result <= 12'b111010101110;
   61970: result <= 12'b111010101110;
   61971: result <= 12'b111010101110;
   61972: result <= 12'b111010101110;
   61973: result <= 12'b111010101110;
   61974: result <= 12'b111010101101;
   61975: result <= 12'b111010101101;
   61976: result <= 12'b111010101101;
   61977: result <= 12'b111010101101;
   61978: result <= 12'b111010101101;
   61979: result <= 12'b111010101100;
   61980: result <= 12'b111010101100;
   61981: result <= 12'b111010101100;
   61982: result <= 12'b111010101100;
   61983: result <= 12'b111010101100;
   61984: result <= 12'b111010101100;
   61985: result <= 12'b111010101011;
   61986: result <= 12'b111010101011;
   61987: result <= 12'b111010101011;
   61988: result <= 12'b111010101011;
   61989: result <= 12'b111010101011;
   61990: result <= 12'b111010101010;
   61991: result <= 12'b111010101010;
   61992: result <= 12'b111010101010;
   61993: result <= 12'b111010101010;
   61994: result <= 12'b111010101010;
   61995: result <= 12'b111010101001;
   61996: result <= 12'b111010101001;
   61997: result <= 12'b111010101001;
   61998: result <= 12'b111010101001;
   61999: result <= 12'b111010101001;
   62000: result <= 12'b111010101001;
   62001: result <= 12'b111010101000;
   62002: result <= 12'b111010101000;
   62003: result <= 12'b111010101000;
   62004: result <= 12'b111010101000;
   62005: result <= 12'b111010101000;
   62006: result <= 12'b111010100111;
   62007: result <= 12'b111010100111;
   62008: result <= 12'b111010100111;
   62009: result <= 12'b111010100111;
   62010: result <= 12'b111010100111;
   62011: result <= 12'b111010100111;
   62012: result <= 12'b111010100110;
   62013: result <= 12'b111010100110;
   62014: result <= 12'b111010100110;
   62015: result <= 12'b111010100110;
   62016: result <= 12'b111010100110;
   62017: result <= 12'b111010100101;
   62018: result <= 12'b111010100101;
   62019: result <= 12'b111010100101;
   62020: result <= 12'b111010100101;
   62021: result <= 12'b111010100101;
   62022: result <= 12'b111010100100;
   62023: result <= 12'b111010100100;
   62024: result <= 12'b111010100100;
   62025: result <= 12'b111010100100;
   62026: result <= 12'b111010100100;
   62027: result <= 12'b111010100100;
   62028: result <= 12'b111010100011;
   62029: result <= 12'b111010100011;
   62030: result <= 12'b111010100011;
   62031: result <= 12'b111010100011;
   62032: result <= 12'b111010100011;
   62033: result <= 12'b111010100010;
   62034: result <= 12'b111010100010;
   62035: result <= 12'b111010100010;
   62036: result <= 12'b111010100010;
   62037: result <= 12'b111010100010;
   62038: result <= 12'b111010100010;
   62039: result <= 12'b111010100001;
   62040: result <= 12'b111010100001;
   62041: result <= 12'b111010100001;
   62042: result <= 12'b111010100001;
   62043: result <= 12'b111010100001;
   62044: result <= 12'b111010100000;
   62045: result <= 12'b111010100000;
   62046: result <= 12'b111010100000;
   62047: result <= 12'b111010100000;
   62048: result <= 12'b111010100000;
   62049: result <= 12'b111010011111;
   62050: result <= 12'b111010011111;
   62051: result <= 12'b111010011111;
   62052: result <= 12'b111010011111;
   62053: result <= 12'b111010011111;
   62054: result <= 12'b111010011111;
   62055: result <= 12'b111010011110;
   62056: result <= 12'b111010011110;
   62057: result <= 12'b111010011110;
   62058: result <= 12'b111010011110;
   62059: result <= 12'b111010011110;
   62060: result <= 12'b111010011101;
   62061: result <= 12'b111010011101;
   62062: result <= 12'b111010011101;
   62063: result <= 12'b111010011101;
   62064: result <= 12'b111010011101;
   62065: result <= 12'b111010011101;
   62066: result <= 12'b111010011100;
   62067: result <= 12'b111010011100;
   62068: result <= 12'b111010011100;
   62069: result <= 12'b111010011100;
   62070: result <= 12'b111010011100;
   62071: result <= 12'b111010011011;
   62072: result <= 12'b111010011011;
   62073: result <= 12'b111010011011;
   62074: result <= 12'b111010011011;
   62075: result <= 12'b111010011011;
   62076: result <= 12'b111010011010;
   62077: result <= 12'b111010011010;
   62078: result <= 12'b111010011010;
   62079: result <= 12'b111010011010;
   62080: result <= 12'b111010011010;
   62081: result <= 12'b111010011010;
   62082: result <= 12'b111010011001;
   62083: result <= 12'b111010011001;
   62084: result <= 12'b111010011001;
   62085: result <= 12'b111010011001;
   62086: result <= 12'b111010011001;
   62087: result <= 12'b111010011000;
   62088: result <= 12'b111010011000;
   62089: result <= 12'b111010011000;
   62090: result <= 12'b111010011000;
   62091: result <= 12'b111010011000;
   62092: result <= 12'b111010011000;
   62093: result <= 12'b111010010111;
   62094: result <= 12'b111010010111;
   62095: result <= 12'b111010010111;
   62096: result <= 12'b111010010111;
   62097: result <= 12'b111010010111;
   62098: result <= 12'b111010010110;
   62099: result <= 12'b111010010110;
   62100: result <= 12'b111010010110;
   62101: result <= 12'b111010010110;
   62102: result <= 12'b111010010110;
   62103: result <= 12'b111010010101;
   62104: result <= 12'b111010010101;
   62105: result <= 12'b111010010101;
   62106: result <= 12'b111010010101;
   62107: result <= 12'b111010010101;
   62108: result <= 12'b111010010101;
   62109: result <= 12'b111010010100;
   62110: result <= 12'b111010010100;
   62111: result <= 12'b111010010100;
   62112: result <= 12'b111010010100;
   62113: result <= 12'b111010010100;
   62114: result <= 12'b111010010011;
   62115: result <= 12'b111010010011;
   62116: result <= 12'b111010010011;
   62117: result <= 12'b111010010011;
   62118: result <= 12'b111010010011;
   62119: result <= 12'b111010010010;
   62120: result <= 12'b111010010010;
   62121: result <= 12'b111010010010;
   62122: result <= 12'b111010010010;
   62123: result <= 12'b111010010010;
   62124: result <= 12'b111010010010;
   62125: result <= 12'b111010010001;
   62126: result <= 12'b111010010001;
   62127: result <= 12'b111010010001;
   62128: result <= 12'b111010010001;
   62129: result <= 12'b111010010001;
   62130: result <= 12'b111010010000;
   62131: result <= 12'b111010010000;
   62132: result <= 12'b111010010000;
   62133: result <= 12'b111010010000;
   62134: result <= 12'b111010010000;
   62135: result <= 12'b111010010000;
   62136: result <= 12'b111010001111;
   62137: result <= 12'b111010001111;
   62138: result <= 12'b111010001111;
   62139: result <= 12'b111010001111;
   62140: result <= 12'b111010001111;
   62141: result <= 12'b111010001110;
   62142: result <= 12'b111010001110;
   62143: result <= 12'b111010001110;
   62144: result <= 12'b111010001110;
   62145: result <= 12'b111010001110;
   62146: result <= 12'b111010001101;
   62147: result <= 12'b111010001101;
   62148: result <= 12'b111010001101;
   62149: result <= 12'b111010001101;
   62150: result <= 12'b111010001101;
   62151: result <= 12'b111010001101;
   62152: result <= 12'b111010001100;
   62153: result <= 12'b111010001100;
   62154: result <= 12'b111010001100;
   62155: result <= 12'b111010001100;
   62156: result <= 12'b111010001100;
   62157: result <= 12'b111010001011;
   62158: result <= 12'b111010001011;
   62159: result <= 12'b111010001011;
   62160: result <= 12'b111010001011;
   62161: result <= 12'b111010001011;
   62162: result <= 12'b111010001010;
   62163: result <= 12'b111010001010;
   62164: result <= 12'b111010001010;
   62165: result <= 12'b111010001010;
   62166: result <= 12'b111010001010;
   62167: result <= 12'b111010001010;
   62168: result <= 12'b111010001001;
   62169: result <= 12'b111010001001;
   62170: result <= 12'b111010001001;
   62171: result <= 12'b111010001001;
   62172: result <= 12'b111010001001;
   62173: result <= 12'b111010001000;
   62174: result <= 12'b111010001000;
   62175: result <= 12'b111010001000;
   62176: result <= 12'b111010001000;
   62177: result <= 12'b111010001000;
   62178: result <= 12'b111010001000;
   62179: result <= 12'b111010000111;
   62180: result <= 12'b111010000111;
   62181: result <= 12'b111010000111;
   62182: result <= 12'b111010000111;
   62183: result <= 12'b111010000111;
   62184: result <= 12'b111010000110;
   62185: result <= 12'b111010000110;
   62186: result <= 12'b111010000110;
   62187: result <= 12'b111010000110;
   62188: result <= 12'b111010000110;
   62189: result <= 12'b111010000101;
   62190: result <= 12'b111010000101;
   62191: result <= 12'b111010000101;
   62192: result <= 12'b111010000101;
   62193: result <= 12'b111010000101;
   62194: result <= 12'b111010000101;
   62195: result <= 12'b111010000100;
   62196: result <= 12'b111010000100;
   62197: result <= 12'b111010000100;
   62198: result <= 12'b111010000100;
   62199: result <= 12'b111010000100;
   62200: result <= 12'b111010000011;
   62201: result <= 12'b111010000011;
   62202: result <= 12'b111010000011;
   62203: result <= 12'b111010000011;
   62204: result <= 12'b111010000011;
   62205: result <= 12'b111010000010;
   62206: result <= 12'b111010000010;
   62207: result <= 12'b111010000010;
   62208: result <= 12'b111010000010;
   62209: result <= 12'b111010000010;
   62210: result <= 12'b111010000010;
   62211: result <= 12'b111010000001;
   62212: result <= 12'b111010000001;
   62213: result <= 12'b111010000001;
   62214: result <= 12'b111010000001;
   62215: result <= 12'b111010000001;
   62216: result <= 12'b111010000000;
   62217: result <= 12'b111010000000;
   62218: result <= 12'b111010000000;
   62219: result <= 12'b111010000000;
   62220: result <= 12'b111010000000;
   62221: result <= 12'b111001111111;
   62222: result <= 12'b111001111111;
   62223: result <= 12'b111001111111;
   62224: result <= 12'b111001111111;
   62225: result <= 12'b111001111111;
   62226: result <= 12'b111001111111;
   62227: result <= 12'b111001111110;
   62228: result <= 12'b111001111110;
   62229: result <= 12'b111001111110;
   62230: result <= 12'b111001111110;
   62231: result <= 12'b111001111110;
   62232: result <= 12'b111001111101;
   62233: result <= 12'b111001111101;
   62234: result <= 12'b111001111101;
   62235: result <= 12'b111001111101;
   62236: result <= 12'b111001111101;
   62237: result <= 12'b111001111101;
   62238: result <= 12'b111001111100;
   62239: result <= 12'b111001111100;
   62240: result <= 12'b111001111100;
   62241: result <= 12'b111001111100;
   62242: result <= 12'b111001111100;
   62243: result <= 12'b111001111011;
   62244: result <= 12'b111001111011;
   62245: result <= 12'b111001111011;
   62246: result <= 12'b111001111011;
   62247: result <= 12'b111001111011;
   62248: result <= 12'b111001111010;
   62249: result <= 12'b111001111010;
   62250: result <= 12'b111001111010;
   62251: result <= 12'b111001111010;
   62252: result <= 12'b111001111010;
   62253: result <= 12'b111001111010;
   62254: result <= 12'b111001111001;
   62255: result <= 12'b111001111001;
   62256: result <= 12'b111001111001;
   62257: result <= 12'b111001111001;
   62258: result <= 12'b111001111001;
   62259: result <= 12'b111001111000;
   62260: result <= 12'b111001111000;
   62261: result <= 12'b111001111000;
   62262: result <= 12'b111001111000;
   62263: result <= 12'b111001111000;
   62264: result <= 12'b111001110111;
   62265: result <= 12'b111001110111;
   62266: result <= 12'b111001110111;
   62267: result <= 12'b111001110111;
   62268: result <= 12'b111001110111;
   62269: result <= 12'b111001110111;
   62270: result <= 12'b111001110110;
   62271: result <= 12'b111001110110;
   62272: result <= 12'b111001110110;
   62273: result <= 12'b111001110110;
   62274: result <= 12'b111001110110;
   62275: result <= 12'b111001110101;
   62276: result <= 12'b111001110101;
   62277: result <= 12'b111001110101;
   62278: result <= 12'b111001110101;
   62279: result <= 12'b111001110101;
   62280: result <= 12'b111001110100;
   62281: result <= 12'b111001110100;
   62282: result <= 12'b111001110100;
   62283: result <= 12'b111001110100;
   62284: result <= 12'b111001110100;
   62285: result <= 12'b111001110100;
   62286: result <= 12'b111001110011;
   62287: result <= 12'b111001110011;
   62288: result <= 12'b111001110011;
   62289: result <= 12'b111001110011;
   62290: result <= 12'b111001110011;
   62291: result <= 12'b111001110010;
   62292: result <= 12'b111001110010;
   62293: result <= 12'b111001110010;
   62294: result <= 12'b111001110010;
   62295: result <= 12'b111001110010;
   62296: result <= 12'b111001110001;
   62297: result <= 12'b111001110001;
   62298: result <= 12'b111001110001;
   62299: result <= 12'b111001110001;
   62300: result <= 12'b111001110001;
   62301: result <= 12'b111001110001;
   62302: result <= 12'b111001110000;
   62303: result <= 12'b111001110000;
   62304: result <= 12'b111001110000;
   62305: result <= 12'b111001110000;
   62306: result <= 12'b111001110000;
   62307: result <= 12'b111001101111;
   62308: result <= 12'b111001101111;
   62309: result <= 12'b111001101111;
   62310: result <= 12'b111001101111;
   62311: result <= 12'b111001101111;
   62312: result <= 12'b111001101110;
   62313: result <= 12'b111001101110;
   62314: result <= 12'b111001101110;
   62315: result <= 12'b111001101110;
   62316: result <= 12'b111001101110;
   62317: result <= 12'b111001101110;
   62318: result <= 12'b111001101101;
   62319: result <= 12'b111001101101;
   62320: result <= 12'b111001101101;
   62321: result <= 12'b111001101101;
   62322: result <= 12'b111001101101;
   62323: result <= 12'b111001101100;
   62324: result <= 12'b111001101100;
   62325: result <= 12'b111001101100;
   62326: result <= 12'b111001101100;
   62327: result <= 12'b111001101100;
   62328: result <= 12'b111001101100;
   62329: result <= 12'b111001101011;
   62330: result <= 12'b111001101011;
   62331: result <= 12'b111001101011;
   62332: result <= 12'b111001101011;
   62333: result <= 12'b111001101011;
   62334: result <= 12'b111001101010;
   62335: result <= 12'b111001101010;
   62336: result <= 12'b111001101010;
   62337: result <= 12'b111001101010;
   62338: result <= 12'b111001101010;
   62339: result <= 12'b111001101001;
   62340: result <= 12'b111001101001;
   62341: result <= 12'b111001101001;
   62342: result <= 12'b111001101001;
   62343: result <= 12'b111001101001;
   62344: result <= 12'b111001101001;
   62345: result <= 12'b111001101000;
   62346: result <= 12'b111001101000;
   62347: result <= 12'b111001101000;
   62348: result <= 12'b111001101000;
   62349: result <= 12'b111001101000;
   62350: result <= 12'b111001100111;
   62351: result <= 12'b111001100111;
   62352: result <= 12'b111001100111;
   62353: result <= 12'b111001100111;
   62354: result <= 12'b111001100111;
   62355: result <= 12'b111001100110;
   62356: result <= 12'b111001100110;
   62357: result <= 12'b111001100110;
   62358: result <= 12'b111001100110;
   62359: result <= 12'b111001100110;
   62360: result <= 12'b111001100110;
   62361: result <= 12'b111001100101;
   62362: result <= 12'b111001100101;
   62363: result <= 12'b111001100101;
   62364: result <= 12'b111001100101;
   62365: result <= 12'b111001100101;
   62366: result <= 12'b111001100100;
   62367: result <= 12'b111001100100;
   62368: result <= 12'b111001100100;
   62369: result <= 12'b111001100100;
   62370: result <= 12'b111001100100;
   62371: result <= 12'b111001100011;
   62372: result <= 12'b111001100011;
   62373: result <= 12'b111001100011;
   62374: result <= 12'b111001100011;
   62375: result <= 12'b111001100011;
   62376: result <= 12'b111001100011;
   62377: result <= 12'b111001100010;
   62378: result <= 12'b111001100010;
   62379: result <= 12'b111001100010;
   62380: result <= 12'b111001100010;
   62381: result <= 12'b111001100010;
   62382: result <= 12'b111001100001;
   62383: result <= 12'b111001100001;
   62384: result <= 12'b111001100001;
   62385: result <= 12'b111001100001;
   62386: result <= 12'b111001100001;
   62387: result <= 12'b111001100000;
   62388: result <= 12'b111001100000;
   62389: result <= 12'b111001100000;
   62390: result <= 12'b111001100000;
   62391: result <= 12'b111001100000;
   62392: result <= 12'b111001100000;
   62393: result <= 12'b111001011111;
   62394: result <= 12'b111001011111;
   62395: result <= 12'b111001011111;
   62396: result <= 12'b111001011111;
   62397: result <= 12'b111001011111;
   62398: result <= 12'b111001011110;
   62399: result <= 12'b111001011110;
   62400: result <= 12'b111001011110;
   62401: result <= 12'b111001011110;
   62402: result <= 12'b111001011110;
   62403: result <= 12'b111001011101;
   62404: result <= 12'b111001011101;
   62405: result <= 12'b111001011101;
   62406: result <= 12'b111001011101;
   62407: result <= 12'b111001011101;
   62408: result <= 12'b111001011101;
   62409: result <= 12'b111001011100;
   62410: result <= 12'b111001011100;
   62411: result <= 12'b111001011100;
   62412: result <= 12'b111001011100;
   62413: result <= 12'b111001011100;
   62414: result <= 12'b111001011011;
   62415: result <= 12'b111001011011;
   62416: result <= 12'b111001011011;
   62417: result <= 12'b111001011011;
   62418: result <= 12'b111001011011;
   62419: result <= 12'b111001011010;
   62420: result <= 12'b111001011010;
   62421: result <= 12'b111001011010;
   62422: result <= 12'b111001011010;
   62423: result <= 12'b111001011010;
   62424: result <= 12'b111001011010;
   62425: result <= 12'b111001011001;
   62426: result <= 12'b111001011001;
   62427: result <= 12'b111001011001;
   62428: result <= 12'b111001011001;
   62429: result <= 12'b111001011001;
   62430: result <= 12'b111001011000;
   62431: result <= 12'b111001011000;
   62432: result <= 12'b111001011000;
   62433: result <= 12'b111001011000;
   62434: result <= 12'b111001011000;
   62435: result <= 12'b111001010111;
   62436: result <= 12'b111001010111;
   62437: result <= 12'b111001010111;
   62438: result <= 12'b111001010111;
   62439: result <= 12'b111001010111;
   62440: result <= 12'b111001010111;
   62441: result <= 12'b111001010110;
   62442: result <= 12'b111001010110;
   62443: result <= 12'b111001010110;
   62444: result <= 12'b111001010110;
   62445: result <= 12'b111001010110;
   62446: result <= 12'b111001010101;
   62447: result <= 12'b111001010101;
   62448: result <= 12'b111001010101;
   62449: result <= 12'b111001010101;
   62450: result <= 12'b111001010101;
   62451: result <= 12'b111001010100;
   62452: result <= 12'b111001010100;
   62453: result <= 12'b111001010100;
   62454: result <= 12'b111001010100;
   62455: result <= 12'b111001010100;
   62456: result <= 12'b111001010100;
   62457: result <= 12'b111001010011;
   62458: result <= 12'b111001010011;
   62459: result <= 12'b111001010011;
   62460: result <= 12'b111001010011;
   62461: result <= 12'b111001010011;
   62462: result <= 12'b111001010010;
   62463: result <= 12'b111001010010;
   62464: result <= 12'b111001010010;
   62465: result <= 12'b111001010010;
   62466: result <= 12'b111001010010;
   62467: result <= 12'b111001010001;
   62468: result <= 12'b111001010001;
   62469: result <= 12'b111001010001;
   62470: result <= 12'b111001010001;
   62471: result <= 12'b111001010001;
   62472: result <= 12'b111001010000;
   62473: result <= 12'b111001010000;
   62474: result <= 12'b111001010000;
   62475: result <= 12'b111001010000;
   62476: result <= 12'b111001010000;
   62477: result <= 12'b111001010000;
   62478: result <= 12'b111001001111;
   62479: result <= 12'b111001001111;
   62480: result <= 12'b111001001111;
   62481: result <= 12'b111001001111;
   62482: result <= 12'b111001001111;
   62483: result <= 12'b111001001110;
   62484: result <= 12'b111001001110;
   62485: result <= 12'b111001001110;
   62486: result <= 12'b111001001110;
   62487: result <= 12'b111001001110;
   62488: result <= 12'b111001001101;
   62489: result <= 12'b111001001101;
   62490: result <= 12'b111001001101;
   62491: result <= 12'b111001001101;
   62492: result <= 12'b111001001101;
   62493: result <= 12'b111001001101;
   62494: result <= 12'b111001001100;
   62495: result <= 12'b111001001100;
   62496: result <= 12'b111001001100;
   62497: result <= 12'b111001001100;
   62498: result <= 12'b111001001100;
   62499: result <= 12'b111001001011;
   62500: result <= 12'b111001001011;
   62501: result <= 12'b111001001011;
   62502: result <= 12'b111001001011;
   62503: result <= 12'b111001001011;
   62504: result <= 12'b111001001010;
   62505: result <= 12'b111001001010;
   62506: result <= 12'b111001001010;
   62507: result <= 12'b111001001010;
   62508: result <= 12'b111001001010;
   62509: result <= 12'b111001001010;
   62510: result <= 12'b111001001001;
   62511: result <= 12'b111001001001;
   62512: result <= 12'b111001001001;
   62513: result <= 12'b111001001001;
   62514: result <= 12'b111001001001;
   62515: result <= 12'b111001001000;
   62516: result <= 12'b111001001000;
   62517: result <= 12'b111001001000;
   62518: result <= 12'b111001001000;
   62519: result <= 12'b111001001000;
   62520: result <= 12'b111001000111;
   62521: result <= 12'b111001000111;
   62522: result <= 12'b111001000111;
   62523: result <= 12'b111001000111;
   62524: result <= 12'b111001000111;
   62525: result <= 12'b111001000111;
   62526: result <= 12'b111001000110;
   62527: result <= 12'b111001000110;
   62528: result <= 12'b111001000110;
   62529: result <= 12'b111001000110;
   62530: result <= 12'b111001000110;
   62531: result <= 12'b111001000101;
   62532: result <= 12'b111001000101;
   62533: result <= 12'b111001000101;
   62534: result <= 12'b111001000101;
   62535: result <= 12'b111001000101;
   62536: result <= 12'b111001000100;
   62537: result <= 12'b111001000100;
   62538: result <= 12'b111001000100;
   62539: result <= 12'b111001000100;
   62540: result <= 12'b111001000100;
   62541: result <= 12'b111001000100;
   62542: result <= 12'b111001000011;
   62543: result <= 12'b111001000011;
   62544: result <= 12'b111001000011;
   62545: result <= 12'b111001000011;
   62546: result <= 12'b111001000011;
   62547: result <= 12'b111001000010;
   62548: result <= 12'b111001000010;
   62549: result <= 12'b111001000010;
   62550: result <= 12'b111001000010;
   62551: result <= 12'b111001000010;
   62552: result <= 12'b111001000001;
   62553: result <= 12'b111001000001;
   62554: result <= 12'b111001000001;
   62555: result <= 12'b111001000001;
   62556: result <= 12'b111001000001;
   62557: result <= 12'b111001000001;
   62558: result <= 12'b111001000000;
   62559: result <= 12'b111001000000;
   62560: result <= 12'b111001000000;
   62561: result <= 12'b111001000000;
   62562: result <= 12'b111001000000;
   62563: result <= 12'b111000111111;
   62564: result <= 12'b111000111111;
   62565: result <= 12'b111000111111;
   62566: result <= 12'b111000111111;
   62567: result <= 12'b111000111111;
   62568: result <= 12'b111000111110;
   62569: result <= 12'b111000111110;
   62570: result <= 12'b111000111110;
   62571: result <= 12'b111000111110;
   62572: result <= 12'b111000111110;
   62573: result <= 12'b111000111101;
   62574: result <= 12'b111000111101;
   62575: result <= 12'b111000111101;
   62576: result <= 12'b111000111101;
   62577: result <= 12'b111000111101;
   62578: result <= 12'b111000111101;
   62579: result <= 12'b111000111100;
   62580: result <= 12'b111000111100;
   62581: result <= 12'b111000111100;
   62582: result <= 12'b111000111100;
   62583: result <= 12'b111000111100;
   62584: result <= 12'b111000111011;
   62585: result <= 12'b111000111011;
   62586: result <= 12'b111000111011;
   62587: result <= 12'b111000111011;
   62588: result <= 12'b111000111011;
   62589: result <= 12'b111000111010;
   62590: result <= 12'b111000111010;
   62591: result <= 12'b111000111010;
   62592: result <= 12'b111000111010;
   62593: result <= 12'b111000111010;
   62594: result <= 12'b111000111010;
   62595: result <= 12'b111000111001;
   62596: result <= 12'b111000111001;
   62597: result <= 12'b111000111001;
   62598: result <= 12'b111000111001;
   62599: result <= 12'b111000111001;
   62600: result <= 12'b111000111000;
   62601: result <= 12'b111000111000;
   62602: result <= 12'b111000111000;
   62603: result <= 12'b111000111000;
   62604: result <= 12'b111000111000;
   62605: result <= 12'b111000110111;
   62606: result <= 12'b111000110111;
   62607: result <= 12'b111000110111;
   62608: result <= 12'b111000110111;
   62609: result <= 12'b111000110111;
   62610: result <= 12'b111000110111;
   62611: result <= 12'b111000110110;
   62612: result <= 12'b111000110110;
   62613: result <= 12'b111000110110;
   62614: result <= 12'b111000110110;
   62615: result <= 12'b111000110110;
   62616: result <= 12'b111000110101;
   62617: result <= 12'b111000110101;
   62618: result <= 12'b111000110101;
   62619: result <= 12'b111000110101;
   62620: result <= 12'b111000110101;
   62621: result <= 12'b111000110100;
   62622: result <= 12'b111000110100;
   62623: result <= 12'b111000110100;
   62624: result <= 12'b111000110100;
   62625: result <= 12'b111000110100;
   62626: result <= 12'b111000110011;
   62627: result <= 12'b111000110011;
   62628: result <= 12'b111000110011;
   62629: result <= 12'b111000110011;
   62630: result <= 12'b111000110011;
   62631: result <= 12'b111000110011;
   62632: result <= 12'b111000110010;
   62633: result <= 12'b111000110010;
   62634: result <= 12'b111000110010;
   62635: result <= 12'b111000110010;
   62636: result <= 12'b111000110010;
   62637: result <= 12'b111000110001;
   62638: result <= 12'b111000110001;
   62639: result <= 12'b111000110001;
   62640: result <= 12'b111000110001;
   62641: result <= 12'b111000110001;
   62642: result <= 12'b111000110000;
   62643: result <= 12'b111000110000;
   62644: result <= 12'b111000110000;
   62645: result <= 12'b111000110000;
   62646: result <= 12'b111000110000;
   62647: result <= 12'b111000110000;
   62648: result <= 12'b111000101111;
   62649: result <= 12'b111000101111;
   62650: result <= 12'b111000101111;
   62651: result <= 12'b111000101111;
   62652: result <= 12'b111000101111;
   62653: result <= 12'b111000101110;
   62654: result <= 12'b111000101110;
   62655: result <= 12'b111000101110;
   62656: result <= 12'b111000101110;
   62657: result <= 12'b111000101110;
   62658: result <= 12'b111000101101;
   62659: result <= 12'b111000101101;
   62660: result <= 12'b111000101101;
   62661: result <= 12'b111000101101;
   62662: result <= 12'b111000101101;
   62663: result <= 12'b111000101101;
   62664: result <= 12'b111000101100;
   62665: result <= 12'b111000101100;
   62666: result <= 12'b111000101100;
   62667: result <= 12'b111000101100;
   62668: result <= 12'b111000101100;
   62669: result <= 12'b111000101011;
   62670: result <= 12'b111000101011;
   62671: result <= 12'b111000101011;
   62672: result <= 12'b111000101011;
   62673: result <= 12'b111000101011;
   62674: result <= 12'b111000101010;
   62675: result <= 12'b111000101010;
   62676: result <= 12'b111000101010;
   62677: result <= 12'b111000101010;
   62678: result <= 12'b111000101010;
   62679: result <= 12'b111000101001;
   62680: result <= 12'b111000101001;
   62681: result <= 12'b111000101001;
   62682: result <= 12'b111000101001;
   62683: result <= 12'b111000101001;
   62684: result <= 12'b111000101001;
   62685: result <= 12'b111000101000;
   62686: result <= 12'b111000101000;
   62687: result <= 12'b111000101000;
   62688: result <= 12'b111000101000;
   62689: result <= 12'b111000101000;
   62690: result <= 12'b111000100111;
   62691: result <= 12'b111000100111;
   62692: result <= 12'b111000100111;
   62693: result <= 12'b111000100111;
   62694: result <= 12'b111000100111;
   62695: result <= 12'b111000100110;
   62696: result <= 12'b111000100110;
   62697: result <= 12'b111000100110;
   62698: result <= 12'b111000100110;
   62699: result <= 12'b111000100110;
   62700: result <= 12'b111000100110;
   62701: result <= 12'b111000100101;
   62702: result <= 12'b111000100101;
   62703: result <= 12'b111000100101;
   62704: result <= 12'b111000100101;
   62705: result <= 12'b111000100101;
   62706: result <= 12'b111000100100;
   62707: result <= 12'b111000100100;
   62708: result <= 12'b111000100100;
   62709: result <= 12'b111000100100;
   62710: result <= 12'b111000100100;
   62711: result <= 12'b111000100011;
   62712: result <= 12'b111000100011;
   62713: result <= 12'b111000100011;
   62714: result <= 12'b111000100011;
   62715: result <= 12'b111000100011;
   62716: result <= 12'b111000100010;
   62717: result <= 12'b111000100010;
   62718: result <= 12'b111000100010;
   62719: result <= 12'b111000100010;
   62720: result <= 12'b111000100010;
   62721: result <= 12'b111000100010;
   62722: result <= 12'b111000100001;
   62723: result <= 12'b111000100001;
   62724: result <= 12'b111000100001;
   62725: result <= 12'b111000100001;
   62726: result <= 12'b111000100001;
   62727: result <= 12'b111000100000;
   62728: result <= 12'b111000100000;
   62729: result <= 12'b111000100000;
   62730: result <= 12'b111000100000;
   62731: result <= 12'b111000100000;
   62732: result <= 12'b111000011111;
   62733: result <= 12'b111000011111;
   62734: result <= 12'b111000011111;
   62735: result <= 12'b111000011111;
   62736: result <= 12'b111000011111;
   62737: result <= 12'b111000011111;
   62738: result <= 12'b111000011110;
   62739: result <= 12'b111000011110;
   62740: result <= 12'b111000011110;
   62741: result <= 12'b111000011110;
   62742: result <= 12'b111000011110;
   62743: result <= 12'b111000011101;
   62744: result <= 12'b111000011101;
   62745: result <= 12'b111000011101;
   62746: result <= 12'b111000011101;
   62747: result <= 12'b111000011101;
   62748: result <= 12'b111000011100;
   62749: result <= 12'b111000011100;
   62750: result <= 12'b111000011100;
   62751: result <= 12'b111000011100;
   62752: result <= 12'b111000011100;
   62753: result <= 12'b111000011011;
   62754: result <= 12'b111000011011;
   62755: result <= 12'b111000011011;
   62756: result <= 12'b111000011011;
   62757: result <= 12'b111000011011;
   62758: result <= 12'b111000011011;
   62759: result <= 12'b111000011010;
   62760: result <= 12'b111000011010;
   62761: result <= 12'b111000011010;
   62762: result <= 12'b111000011010;
   62763: result <= 12'b111000011010;
   62764: result <= 12'b111000011001;
   62765: result <= 12'b111000011001;
   62766: result <= 12'b111000011001;
   62767: result <= 12'b111000011001;
   62768: result <= 12'b111000011001;
   62769: result <= 12'b111000011000;
   62770: result <= 12'b111000011000;
   62771: result <= 12'b111000011000;
   62772: result <= 12'b111000011000;
   62773: result <= 12'b111000011000;
   62774: result <= 12'b111000011000;
   62775: result <= 12'b111000010111;
   62776: result <= 12'b111000010111;
   62777: result <= 12'b111000010111;
   62778: result <= 12'b111000010111;
   62779: result <= 12'b111000010111;
   62780: result <= 12'b111000010110;
   62781: result <= 12'b111000010110;
   62782: result <= 12'b111000010110;
   62783: result <= 12'b111000010110;
   62784: result <= 12'b111000010110;
   62785: result <= 12'b111000010101;
   62786: result <= 12'b111000010101;
   62787: result <= 12'b111000010101;
   62788: result <= 12'b111000010101;
   62789: result <= 12'b111000010101;
   62790: result <= 12'b111000010100;
   62791: result <= 12'b111000010100;
   62792: result <= 12'b111000010100;
   62793: result <= 12'b111000010100;
   62794: result <= 12'b111000010100;
   62795: result <= 12'b111000010100;
   62796: result <= 12'b111000010011;
   62797: result <= 12'b111000010011;
   62798: result <= 12'b111000010011;
   62799: result <= 12'b111000010011;
   62800: result <= 12'b111000010011;
   62801: result <= 12'b111000010010;
   62802: result <= 12'b111000010010;
   62803: result <= 12'b111000010010;
   62804: result <= 12'b111000010010;
   62805: result <= 12'b111000010010;
   62806: result <= 12'b111000010001;
   62807: result <= 12'b111000010001;
   62808: result <= 12'b111000010001;
   62809: result <= 12'b111000010001;
   62810: result <= 12'b111000010001;
   62811: result <= 12'b111000010000;
   62812: result <= 12'b111000010000;
   62813: result <= 12'b111000010000;
   62814: result <= 12'b111000010000;
   62815: result <= 12'b111000010000;
   62816: result <= 12'b111000010000;
   62817: result <= 12'b111000001111;
   62818: result <= 12'b111000001111;
   62819: result <= 12'b111000001111;
   62820: result <= 12'b111000001111;
   62821: result <= 12'b111000001111;
   62822: result <= 12'b111000001110;
   62823: result <= 12'b111000001110;
   62824: result <= 12'b111000001110;
   62825: result <= 12'b111000001110;
   62826: result <= 12'b111000001110;
   62827: result <= 12'b111000001101;
   62828: result <= 12'b111000001101;
   62829: result <= 12'b111000001101;
   62830: result <= 12'b111000001101;
   62831: result <= 12'b111000001101;
   62832: result <= 12'b111000001101;
   62833: result <= 12'b111000001100;
   62834: result <= 12'b111000001100;
   62835: result <= 12'b111000001100;
   62836: result <= 12'b111000001100;
   62837: result <= 12'b111000001100;
   62838: result <= 12'b111000001011;
   62839: result <= 12'b111000001011;
   62840: result <= 12'b111000001011;
   62841: result <= 12'b111000001011;
   62842: result <= 12'b111000001011;
   62843: result <= 12'b111000001010;
   62844: result <= 12'b111000001010;
   62845: result <= 12'b111000001010;
   62846: result <= 12'b111000001010;
   62847: result <= 12'b111000001010;
   62848: result <= 12'b111000001001;
   62849: result <= 12'b111000001001;
   62850: result <= 12'b111000001001;
   62851: result <= 12'b111000001001;
   62852: result <= 12'b111000001001;
   62853: result <= 12'b111000001001;
   62854: result <= 12'b111000001000;
   62855: result <= 12'b111000001000;
   62856: result <= 12'b111000001000;
   62857: result <= 12'b111000001000;
   62858: result <= 12'b111000001000;
   62859: result <= 12'b111000000111;
   62860: result <= 12'b111000000111;
   62861: result <= 12'b111000000111;
   62862: result <= 12'b111000000111;
   62863: result <= 12'b111000000111;
   62864: result <= 12'b111000000110;
   62865: result <= 12'b111000000110;
   62866: result <= 12'b111000000110;
   62867: result <= 12'b111000000110;
   62868: result <= 12'b111000000110;
   62869: result <= 12'b111000000101;
   62870: result <= 12'b111000000101;
   62871: result <= 12'b111000000101;
   62872: result <= 12'b111000000101;
   62873: result <= 12'b111000000101;
   62874: result <= 12'b111000000101;
   62875: result <= 12'b111000000100;
   62876: result <= 12'b111000000100;
   62877: result <= 12'b111000000100;
   62878: result <= 12'b111000000100;
   62879: result <= 12'b111000000100;
   62880: result <= 12'b111000000011;
   62881: result <= 12'b111000000011;
   62882: result <= 12'b111000000011;
   62883: result <= 12'b111000000011;
   62884: result <= 12'b111000000011;
   62885: result <= 12'b111000000010;
   62886: result <= 12'b111000000010;
   62887: result <= 12'b111000000010;
   62888: result <= 12'b111000000010;
   62889: result <= 12'b111000000010;
   62890: result <= 12'b111000000001;
   62891: result <= 12'b111000000001;
   62892: result <= 12'b111000000001;
   62893: result <= 12'b111000000001;
   62894: result <= 12'b111000000001;
   62895: result <= 12'b111000000001;
   62896: result <= 12'b111000000000;
   62897: result <= 12'b111000000000;
   62898: result <= 12'b111000000000;
   62899: result <= 12'b111000000000;
   62900: result <= 12'b111000000000;
   62901: result <= 12'b111111111111;
   62902: result <= 12'b111111111111;
   62903: result <= 12'b111111111111;
   62904: result <= 12'b111111111111;
   62905: result <= 12'b111111111111;
   62906: result <= 12'b111111111110;
   62907: result <= 12'b111111111110;
   62908: result <= 12'b111111111110;
   62909: result <= 12'b111111111110;
   62910: result <= 12'b111111111110;
   62911: result <= 12'b111111111101;
   62912: result <= 12'b111111111101;
   62913: result <= 12'b111111111101;
   62914: result <= 12'b111111111101;
   62915: result <= 12'b111111111101;
   62916: result <= 12'b111111111101;
   62917: result <= 12'b111111111100;
   62918: result <= 12'b111111111100;
   62919: result <= 12'b111111111100;
   62920: result <= 12'b111111111100;
   62921: result <= 12'b111111111100;
   62922: result <= 12'b111111111011;
   62923: result <= 12'b111111111011;
   62924: result <= 12'b111111111011;
   62925: result <= 12'b111111111011;
   62926: result <= 12'b111111111011;
   62927: result <= 12'b111111111010;
   62928: result <= 12'b111111111010;
   62929: result <= 12'b111111111010;
   62930: result <= 12'b111111111010;
   62931: result <= 12'b111111111010;
   62932: result <= 12'b111111111001;
   62933: result <= 12'b111111111001;
   62934: result <= 12'b111111111001;
   62935: result <= 12'b111111111001;
   62936: result <= 12'b111111111001;
   62937: result <= 12'b111111111001;
   62938: result <= 12'b111111111000;
   62939: result <= 12'b111111111000;
   62940: result <= 12'b111111111000;
   62941: result <= 12'b111111111000;
   62942: result <= 12'b111111111000;
   62943: result <= 12'b111111110111;
   62944: result <= 12'b111111110111;
   62945: result <= 12'b111111110111;
   62946: result <= 12'b111111110111;
   62947: result <= 12'b111111110111;
   62948: result <= 12'b111111110110;
   62949: result <= 12'b111111110110;
   62950: result <= 12'b111111110110;
   62951: result <= 12'b111111110110;
   62952: result <= 12'b111111110110;
   62953: result <= 12'b111111110110;
   62954: result <= 12'b111111110101;
   62955: result <= 12'b111111110101;
   62956: result <= 12'b111111110101;
   62957: result <= 12'b111111110101;
   62958: result <= 12'b111111110101;
   62959: result <= 12'b111111110100;
   62960: result <= 12'b111111110100;
   62961: result <= 12'b111111110100;
   62962: result <= 12'b111111110100;
   62963: result <= 12'b111111110100;
   62964: result <= 12'b111111110011;
   62965: result <= 12'b111111110011;
   62966: result <= 12'b111111110011;
   62967: result <= 12'b111111110011;
   62968: result <= 12'b111111110011;
   62969: result <= 12'b111111110010;
   62970: result <= 12'b111111110010;
   62971: result <= 12'b111111110010;
   62972: result <= 12'b111111110010;
   62973: result <= 12'b111111110010;
   62974: result <= 12'b111111110010;
   62975: result <= 12'b111111110001;
   62976: result <= 12'b111111110001;
   62977: result <= 12'b111111110001;
   62978: result <= 12'b111111110001;
   62979: result <= 12'b111111110001;
   62980: result <= 12'b111111110000;
   62981: result <= 12'b111111110000;
   62982: result <= 12'b111111110000;
   62983: result <= 12'b111111110000;
   62984: result <= 12'b111111110000;
   62985: result <= 12'b111111101111;
   62986: result <= 12'b111111101111;
   62987: result <= 12'b111111101111;
   62988: result <= 12'b111111101111;
   62989: result <= 12'b111111101111;
   62990: result <= 12'b111111101110;
   62991: result <= 12'b111111101110;
   62992: result <= 12'b111111101110;
   62993: result <= 12'b111111101110;
   62994: result <= 12'b111111101110;
   62995: result <= 12'b111111101110;
   62996: result <= 12'b111111101101;
   62997: result <= 12'b111111101101;
   62998: result <= 12'b111111101101;
   62999: result <= 12'b111111101101;
   63000: result <= 12'b111111101101;
   63001: result <= 12'b111111101100;
   63002: result <= 12'b111111101100;
   63003: result <= 12'b111111101100;
   63004: result <= 12'b111111101100;
   63005: result <= 12'b111111101100;
   63006: result <= 12'b111111101011;
   63007: result <= 12'b111111101011;
   63008: result <= 12'b111111101011;
   63009: result <= 12'b111111101011;
   63010: result <= 12'b111111101011;
   63011: result <= 12'b111111101010;
   63012: result <= 12'b111111101010;
   63013: result <= 12'b111111101010;
   63014: result <= 12'b111111101010;
   63015: result <= 12'b111111101010;
   63016: result <= 12'b111111101010;
   63017: result <= 12'b111111101001;
   63018: result <= 12'b111111101001;
   63019: result <= 12'b111111101001;
   63020: result <= 12'b111111101001;
   63021: result <= 12'b111111101001;
   63022: result <= 12'b111111101000;
   63023: result <= 12'b111111101000;
   63024: result <= 12'b111111101000;
   63025: result <= 12'b111111101000;
   63026: result <= 12'b111111101000;
   63027: result <= 12'b111111100111;
   63028: result <= 12'b111111100111;
   63029: result <= 12'b111111100111;
   63030: result <= 12'b111111100111;
   63031: result <= 12'b111111100111;
   63032: result <= 12'b111111100110;
   63033: result <= 12'b111111100110;
   63034: result <= 12'b111111100110;
   63035: result <= 12'b111111100110;
   63036: result <= 12'b111111100110;
   63037: result <= 12'b111111100101;
   63038: result <= 12'b111111100101;
   63039: result <= 12'b111111100101;
   63040: result <= 12'b111111100101;
   63041: result <= 12'b111111100101;
   63042: result <= 12'b111111100101;
   63043: result <= 12'b111111100100;
   63044: result <= 12'b111111100100;
   63045: result <= 12'b111111100100;
   63046: result <= 12'b111111100100;
   63047: result <= 12'b111111100100;
   63048: result <= 12'b111111100011;
   63049: result <= 12'b111111100011;
   63050: result <= 12'b111111100011;
   63051: result <= 12'b111111100011;
   63052: result <= 12'b111111100011;
   63053: result <= 12'b111111100010;
   63054: result <= 12'b111111100010;
   63055: result <= 12'b111111100010;
   63056: result <= 12'b111111100010;
   63057: result <= 12'b111111100010;
   63058: result <= 12'b111111100001;
   63059: result <= 12'b111111100001;
   63060: result <= 12'b111111100001;
   63061: result <= 12'b111111100001;
   63062: result <= 12'b111111100001;
   63063: result <= 12'b111111100001;
   63064: result <= 12'b111111100000;
   63065: result <= 12'b111111100000;
   63066: result <= 12'b111111100000;
   63067: result <= 12'b111111100000;
   63068: result <= 12'b111111100000;
   63069: result <= 12'b111111011111;
   63070: result <= 12'b111111011111;
   63071: result <= 12'b111111011111;
   63072: result <= 12'b111111011111;
   63073: result <= 12'b111111011111;
   63074: result <= 12'b111111011110;
   63075: result <= 12'b111111011110;
   63076: result <= 12'b111111011110;
   63077: result <= 12'b111111011110;
   63078: result <= 12'b111111011110;
   63079: result <= 12'b111111011101;
   63080: result <= 12'b111111011101;
   63081: result <= 12'b111111011101;
   63082: result <= 12'b111111011101;
   63083: result <= 12'b111111011101;
   63084: result <= 12'b111111011101;
   63085: result <= 12'b111111011100;
   63086: result <= 12'b111111011100;
   63087: result <= 12'b111111011100;
   63088: result <= 12'b111111011100;
   63089: result <= 12'b111111011100;
   63090: result <= 12'b111111011011;
   63091: result <= 12'b111111011011;
   63092: result <= 12'b111111011011;
   63093: result <= 12'b111111011011;
   63094: result <= 12'b111111011011;
   63095: result <= 12'b111111011010;
   63096: result <= 12'b111111011010;
   63097: result <= 12'b111111011010;
   63098: result <= 12'b111111011010;
   63099: result <= 12'b111111011010;
   63100: result <= 12'b111111011001;
   63101: result <= 12'b111111011001;
   63102: result <= 12'b111111011001;
   63103: result <= 12'b111111011001;
   63104: result <= 12'b111111011001;
   63105: result <= 12'b111111011001;
   63106: result <= 12'b111111011000;
   63107: result <= 12'b111111011000;
   63108: result <= 12'b111111011000;
   63109: result <= 12'b111111011000;
   63110: result <= 12'b111111011000;
   63111: result <= 12'b111111010111;
   63112: result <= 12'b111111010111;
   63113: result <= 12'b111111010111;
   63114: result <= 12'b111111010111;
   63115: result <= 12'b111111010111;
   63116: result <= 12'b111111010110;
   63117: result <= 12'b111111010110;
   63118: result <= 12'b111111010110;
   63119: result <= 12'b111111010110;
   63120: result <= 12'b111111010110;
   63121: result <= 12'b111111010101;
   63122: result <= 12'b111111010101;
   63123: result <= 12'b111111010101;
   63124: result <= 12'b111111010101;
   63125: result <= 12'b111111010101;
   63126: result <= 12'b111111010101;
   63127: result <= 12'b111111010100;
   63128: result <= 12'b111111010100;
   63129: result <= 12'b111111010100;
   63130: result <= 12'b111111010100;
   63131: result <= 12'b111111010100;
   63132: result <= 12'b111111010011;
   63133: result <= 12'b111111010011;
   63134: result <= 12'b111111010011;
   63135: result <= 12'b111111010011;
   63136: result <= 12'b111111010011;
   63137: result <= 12'b111111010010;
   63138: result <= 12'b111111010010;
   63139: result <= 12'b111111010010;
   63140: result <= 12'b111111010010;
   63141: result <= 12'b111111010010;
   63142: result <= 12'b111111010001;
   63143: result <= 12'b111111010001;
   63144: result <= 12'b111111010001;
   63145: result <= 12'b111111010001;
   63146: result <= 12'b111111010001;
   63147: result <= 12'b111111010000;
   63148: result <= 12'b111111010000;
   63149: result <= 12'b111111010000;
   63150: result <= 12'b111111010000;
   63151: result <= 12'b111111010000;
   63152: result <= 12'b111111010000;
   63153: result <= 12'b111111001111;
   63154: result <= 12'b111111001111;
   63155: result <= 12'b111111001111;
   63156: result <= 12'b111111001111;
   63157: result <= 12'b111111001111;
   63158: result <= 12'b111111001110;
   63159: result <= 12'b111111001110;
   63160: result <= 12'b111111001110;
   63161: result <= 12'b111111001110;
   63162: result <= 12'b111111001110;
   63163: result <= 12'b111111001101;
   63164: result <= 12'b111111001101;
   63165: result <= 12'b111111001101;
   63166: result <= 12'b111111001101;
   63167: result <= 12'b111111001101;
   63168: result <= 12'b111111001100;
   63169: result <= 12'b111111001100;
   63170: result <= 12'b111111001100;
   63171: result <= 12'b111111001100;
   63172: result <= 12'b111111001100;
   63173: result <= 12'b111111001100;
   63174: result <= 12'b111111001011;
   63175: result <= 12'b111111001011;
   63176: result <= 12'b111111001011;
   63177: result <= 12'b111111001011;
   63178: result <= 12'b111111001011;
   63179: result <= 12'b111111001010;
   63180: result <= 12'b111111001010;
   63181: result <= 12'b111111001010;
   63182: result <= 12'b111111001010;
   63183: result <= 12'b111111001010;
   63184: result <= 12'b111111001001;
   63185: result <= 12'b111111001001;
   63186: result <= 12'b111111001001;
   63187: result <= 12'b111111001001;
   63188: result <= 12'b111111001001;
   63189: result <= 12'b111111001000;
   63190: result <= 12'b111111001000;
   63191: result <= 12'b111111001000;
   63192: result <= 12'b111111001000;
   63193: result <= 12'b111111001000;
   63194: result <= 12'b111111000111;
   63195: result <= 12'b111111000111;
   63196: result <= 12'b111111000111;
   63197: result <= 12'b111111000111;
   63198: result <= 12'b111111000111;
   63199: result <= 12'b111111000111;
   63200: result <= 12'b111111000110;
   63201: result <= 12'b111111000110;
   63202: result <= 12'b111111000110;
   63203: result <= 12'b111111000110;
   63204: result <= 12'b111111000110;
   63205: result <= 12'b111111000101;
   63206: result <= 12'b111111000101;
   63207: result <= 12'b111111000101;
   63208: result <= 12'b111111000101;
   63209: result <= 12'b111111000101;
   63210: result <= 12'b111111000100;
   63211: result <= 12'b111111000100;
   63212: result <= 12'b111111000100;
   63213: result <= 12'b111111000100;
   63214: result <= 12'b111111000100;
   63215: result <= 12'b111111000011;
   63216: result <= 12'b111111000011;
   63217: result <= 12'b111111000011;
   63218: result <= 12'b111111000011;
   63219: result <= 12'b111111000011;
   63220: result <= 12'b111111000011;
   63221: result <= 12'b111111000010;
   63222: result <= 12'b111111000010;
   63223: result <= 12'b111111000010;
   63224: result <= 12'b111111000010;
   63225: result <= 12'b111111000010;
   63226: result <= 12'b111111000001;
   63227: result <= 12'b111111000001;
   63228: result <= 12'b111111000001;
   63229: result <= 12'b111111000001;
   63230: result <= 12'b111111000001;
   63231: result <= 12'b111111000000;
   63232: result <= 12'b111111000000;
   63233: result <= 12'b111111000000;
   63234: result <= 12'b111111000000;
   63235: result <= 12'b111111000000;
   63236: result <= 12'b111110111111;
   63237: result <= 12'b111110111111;
   63238: result <= 12'b111110111111;
   63239: result <= 12'b111110111111;
   63240: result <= 12'b111110111111;
   63241: result <= 12'b111110111110;
   63242: result <= 12'b111110111110;
   63243: result <= 12'b111110111110;
   63244: result <= 12'b111110111110;
   63245: result <= 12'b111110111110;
   63246: result <= 12'b111110111110;
   63247: result <= 12'b111110111101;
   63248: result <= 12'b111110111101;
   63249: result <= 12'b111110111101;
   63250: result <= 12'b111110111101;
   63251: result <= 12'b111110111101;
   63252: result <= 12'b111110111100;
   63253: result <= 12'b111110111100;
   63254: result <= 12'b111110111100;
   63255: result <= 12'b111110111100;
   63256: result <= 12'b111110111100;
   63257: result <= 12'b111110111011;
   63258: result <= 12'b111110111011;
   63259: result <= 12'b111110111011;
   63260: result <= 12'b111110111011;
   63261: result <= 12'b111110111011;
   63262: result <= 12'b111110111010;
   63263: result <= 12'b111110111010;
   63264: result <= 12'b111110111010;
   63265: result <= 12'b111110111010;
   63266: result <= 12'b111110111010;
   63267: result <= 12'b111110111010;
   63268: result <= 12'b111110111001;
   63269: result <= 12'b111110111001;
   63270: result <= 12'b111110111001;
   63271: result <= 12'b111110111001;
   63272: result <= 12'b111110111001;
   63273: result <= 12'b111110111000;
   63274: result <= 12'b111110111000;
   63275: result <= 12'b111110111000;
   63276: result <= 12'b111110111000;
   63277: result <= 12'b111110111000;
   63278: result <= 12'b111110110111;
   63279: result <= 12'b111110110111;
   63280: result <= 12'b111110110111;
   63281: result <= 12'b111110110111;
   63282: result <= 12'b111110110111;
   63283: result <= 12'b111110110110;
   63284: result <= 12'b111110110110;
   63285: result <= 12'b111110110110;
   63286: result <= 12'b111110110110;
   63287: result <= 12'b111110110110;
   63288: result <= 12'b111110110101;
   63289: result <= 12'b111110110101;
   63290: result <= 12'b111110110101;
   63291: result <= 12'b111110110101;
   63292: result <= 12'b111110110101;
   63293: result <= 12'b111110110101;
   63294: result <= 12'b111110110100;
   63295: result <= 12'b111110110100;
   63296: result <= 12'b111110110100;
   63297: result <= 12'b111110110100;
   63298: result <= 12'b111110110100;
   63299: result <= 12'b111110110011;
   63300: result <= 12'b111110110011;
   63301: result <= 12'b111110110011;
   63302: result <= 12'b111110110011;
   63303: result <= 12'b111110110011;
   63304: result <= 12'b111110110010;
   63305: result <= 12'b111110110010;
   63306: result <= 12'b111110110010;
   63307: result <= 12'b111110110010;
   63308: result <= 12'b111110110010;
   63309: result <= 12'b111110110001;
   63310: result <= 12'b111110110001;
   63311: result <= 12'b111110110001;
   63312: result <= 12'b111110110001;
   63313: result <= 12'b111110110001;
   63314: result <= 12'b111110110000;
   63315: result <= 12'b111110110000;
   63316: result <= 12'b111110110000;
   63317: result <= 12'b111110110000;
   63318: result <= 12'b111110110000;
   63319: result <= 12'b111110110000;
   63320: result <= 12'b111110101111;
   63321: result <= 12'b111110101111;
   63322: result <= 12'b111110101111;
   63323: result <= 12'b111110101111;
   63324: result <= 12'b111110101111;
   63325: result <= 12'b111110101110;
   63326: result <= 12'b111110101110;
   63327: result <= 12'b111110101110;
   63328: result <= 12'b111110101110;
   63329: result <= 12'b111110101110;
   63330: result <= 12'b111110101101;
   63331: result <= 12'b111110101101;
   63332: result <= 12'b111110101101;
   63333: result <= 12'b111110101101;
   63334: result <= 12'b111110101101;
   63335: result <= 12'b111110101100;
   63336: result <= 12'b111110101100;
   63337: result <= 12'b111110101100;
   63338: result <= 12'b111110101100;
   63339: result <= 12'b111110101100;
   63340: result <= 12'b111110101100;
   63341: result <= 12'b111110101011;
   63342: result <= 12'b111110101011;
   63343: result <= 12'b111110101011;
   63344: result <= 12'b111110101011;
   63345: result <= 12'b111110101011;
   63346: result <= 12'b111110101010;
   63347: result <= 12'b111110101010;
   63348: result <= 12'b111110101010;
   63349: result <= 12'b111110101010;
   63350: result <= 12'b111110101010;
   63351: result <= 12'b111110101001;
   63352: result <= 12'b111110101001;
   63353: result <= 12'b111110101001;
   63354: result <= 12'b111110101001;
   63355: result <= 12'b111110101001;
   63356: result <= 12'b111110101000;
   63357: result <= 12'b111110101000;
   63358: result <= 12'b111110101000;
   63359: result <= 12'b111110101000;
   63360: result <= 12'b111110101000;
   63361: result <= 12'b111110100111;
   63362: result <= 12'b111110100111;
   63363: result <= 12'b111110100111;
   63364: result <= 12'b111110100111;
   63365: result <= 12'b111110100111;
   63366: result <= 12'b111110100111;
   63367: result <= 12'b111110100110;
   63368: result <= 12'b111110100110;
   63369: result <= 12'b111110100110;
   63370: result <= 12'b111110100110;
   63371: result <= 12'b111110100110;
   63372: result <= 12'b111110100101;
   63373: result <= 12'b111110100101;
   63374: result <= 12'b111110100101;
   63375: result <= 12'b111110100101;
   63376: result <= 12'b111110100101;
   63377: result <= 12'b111110100100;
   63378: result <= 12'b111110100100;
   63379: result <= 12'b111110100100;
   63380: result <= 12'b111110100100;
   63381: result <= 12'b111110100100;
   63382: result <= 12'b111110100011;
   63383: result <= 12'b111110100011;
   63384: result <= 12'b111110100011;
   63385: result <= 12'b111110100011;
   63386: result <= 12'b111110100011;
   63387: result <= 12'b111110100010;
   63388: result <= 12'b111110100010;
   63389: result <= 12'b111110100010;
   63390: result <= 12'b111110100010;
   63391: result <= 12'b111110100010;
   63392: result <= 12'b111110100010;
   63393: result <= 12'b111110100001;
   63394: result <= 12'b111110100001;
   63395: result <= 12'b111110100001;
   63396: result <= 12'b111110100001;
   63397: result <= 12'b111110100001;
   63398: result <= 12'b111110100000;
   63399: result <= 12'b111110100000;
   63400: result <= 12'b111110100000;
   63401: result <= 12'b111110100000;
   63402: result <= 12'b111110100000;
   63403: result <= 12'b111110011111;
   63404: result <= 12'b111110011111;
   63405: result <= 12'b111110011111;
   63406: result <= 12'b111110011111;
   63407: result <= 12'b111110011111;
   63408: result <= 12'b111110011110;
   63409: result <= 12'b111110011110;
   63410: result <= 12'b111110011110;
   63411: result <= 12'b111110011110;
   63412: result <= 12'b111110011110;
   63413: result <= 12'b111110011101;
   63414: result <= 12'b111110011101;
   63415: result <= 12'b111110011101;
   63416: result <= 12'b111110011101;
   63417: result <= 12'b111110011101;
   63418: result <= 12'b111110011101;
   63419: result <= 12'b111110011100;
   63420: result <= 12'b111110011100;
   63421: result <= 12'b111110011100;
   63422: result <= 12'b111110011100;
   63423: result <= 12'b111110011100;
   63424: result <= 12'b111110011011;
   63425: result <= 12'b111110011011;
   63426: result <= 12'b111110011011;
   63427: result <= 12'b111110011011;
   63428: result <= 12'b111110011011;
   63429: result <= 12'b111110011010;
   63430: result <= 12'b111110011010;
   63431: result <= 12'b111110011010;
   63432: result <= 12'b111110011010;
   63433: result <= 12'b111110011010;
   63434: result <= 12'b111110011001;
   63435: result <= 12'b111110011001;
   63436: result <= 12'b111110011001;
   63437: result <= 12'b111110011001;
   63438: result <= 12'b111110011001;
   63439: result <= 12'b111110011000;
   63440: result <= 12'b111110011000;
   63441: result <= 12'b111110011000;
   63442: result <= 12'b111110011000;
   63443: result <= 12'b111110011000;
   63444: result <= 12'b111110011000;
   63445: result <= 12'b111110010111;
   63446: result <= 12'b111110010111;
   63447: result <= 12'b111110010111;
   63448: result <= 12'b111110010111;
   63449: result <= 12'b111110010111;
   63450: result <= 12'b111110010110;
   63451: result <= 12'b111110010110;
   63452: result <= 12'b111110010110;
   63453: result <= 12'b111110010110;
   63454: result <= 12'b111110010110;
   63455: result <= 12'b111110010101;
   63456: result <= 12'b111110010101;
   63457: result <= 12'b111110010101;
   63458: result <= 12'b111110010101;
   63459: result <= 12'b111110010101;
   63460: result <= 12'b111110010100;
   63461: result <= 12'b111110010100;
   63462: result <= 12'b111110010100;
   63463: result <= 12'b111110010100;
   63464: result <= 12'b111110010100;
   63465: result <= 12'b111110010011;
   63466: result <= 12'b111110010011;
   63467: result <= 12'b111110010011;
   63468: result <= 12'b111110010011;
   63469: result <= 12'b111110010011;
   63470: result <= 12'b111110010011;
   63471: result <= 12'b111110010010;
   63472: result <= 12'b111110010010;
   63473: result <= 12'b111110010010;
   63474: result <= 12'b111110010010;
   63475: result <= 12'b111110010010;
   63476: result <= 12'b111110010001;
   63477: result <= 12'b111110010001;
   63478: result <= 12'b111110010001;
   63479: result <= 12'b111110010001;
   63480: result <= 12'b111110010001;
   63481: result <= 12'b111110010000;
   63482: result <= 12'b111110010000;
   63483: result <= 12'b111110010000;
   63484: result <= 12'b111110010000;
   63485: result <= 12'b111110010000;
   63486: result <= 12'b111110001111;
   63487: result <= 12'b111110001111;
   63488: result <= 12'b111110001111;
   63489: result <= 12'b111110001111;
   63490: result <= 12'b111110001111;
   63491: result <= 12'b111110001110;
   63492: result <= 12'b111110001110;
   63493: result <= 12'b111110001110;
   63494: result <= 12'b111110001110;
   63495: result <= 12'b111110001110;
   63496: result <= 12'b111110001110;
   63497: result <= 12'b111110001101;
   63498: result <= 12'b111110001101;
   63499: result <= 12'b111110001101;
   63500: result <= 12'b111110001101;
   63501: result <= 12'b111110001101;
   63502: result <= 12'b111110001100;
   63503: result <= 12'b111110001100;
   63504: result <= 12'b111110001100;
   63505: result <= 12'b111110001100;
   63506: result <= 12'b111110001100;
   63507: result <= 12'b111110001011;
   63508: result <= 12'b111110001011;
   63509: result <= 12'b111110001011;
   63510: result <= 12'b111110001011;
   63511: result <= 12'b111110001011;
   63512: result <= 12'b111110001010;
   63513: result <= 12'b111110001010;
   63514: result <= 12'b111110001010;
   63515: result <= 12'b111110001010;
   63516: result <= 12'b111110001010;
   63517: result <= 12'b111110001001;
   63518: result <= 12'b111110001001;
   63519: result <= 12'b111110001001;
   63520: result <= 12'b111110001001;
   63521: result <= 12'b111110001001;
   63522: result <= 12'b111110001000;
   63523: result <= 12'b111110001000;
   63524: result <= 12'b111110001000;
   63525: result <= 12'b111110001000;
   63526: result <= 12'b111110001000;
   63527: result <= 12'b111110001000;
   63528: result <= 12'b111110000111;
   63529: result <= 12'b111110000111;
   63530: result <= 12'b111110000111;
   63531: result <= 12'b111110000111;
   63532: result <= 12'b111110000111;
   63533: result <= 12'b111110000110;
   63534: result <= 12'b111110000110;
   63535: result <= 12'b111110000110;
   63536: result <= 12'b111110000110;
   63537: result <= 12'b111110000110;
   63538: result <= 12'b111110000101;
   63539: result <= 12'b111110000101;
   63540: result <= 12'b111110000101;
   63541: result <= 12'b111110000101;
   63542: result <= 12'b111110000101;
   63543: result <= 12'b111110000100;
   63544: result <= 12'b111110000100;
   63545: result <= 12'b111110000100;
   63546: result <= 12'b111110000100;
   63547: result <= 12'b111110000100;
   63548: result <= 12'b111110000011;
   63549: result <= 12'b111110000011;
   63550: result <= 12'b111110000011;
   63551: result <= 12'b111110000011;
   63552: result <= 12'b111110000011;
   63553: result <= 12'b111110000011;
   63554: result <= 12'b111110000010;
   63555: result <= 12'b111110000010;
   63556: result <= 12'b111110000010;
   63557: result <= 12'b111110000010;
   63558: result <= 12'b111110000010;
   63559: result <= 12'b111110000001;
   63560: result <= 12'b111110000001;
   63561: result <= 12'b111110000001;
   63562: result <= 12'b111110000001;
   63563: result <= 12'b111110000001;
   63564: result <= 12'b111110000000;
   63565: result <= 12'b111110000000;
   63566: result <= 12'b111110000000;
   63567: result <= 12'b111110000000;
   63568: result <= 12'b111110000000;
   63569: result <= 12'b111101111111;
   63570: result <= 12'b111101111111;
   63571: result <= 12'b111101111111;
   63572: result <= 12'b111101111111;
   63573: result <= 12'b111101111111;
   63574: result <= 12'b111101111110;
   63575: result <= 12'b111101111110;
   63576: result <= 12'b111101111110;
   63577: result <= 12'b111101111110;
   63578: result <= 12'b111101111110;
   63579: result <= 12'b111101111110;
   63580: result <= 12'b111101111101;
   63581: result <= 12'b111101111101;
   63582: result <= 12'b111101111101;
   63583: result <= 12'b111101111101;
   63584: result <= 12'b111101111101;
   63585: result <= 12'b111101111100;
   63586: result <= 12'b111101111100;
   63587: result <= 12'b111101111100;
   63588: result <= 12'b111101111100;
   63589: result <= 12'b111101111100;
   63590: result <= 12'b111101111011;
   63591: result <= 12'b111101111011;
   63592: result <= 12'b111101111011;
   63593: result <= 12'b111101111011;
   63594: result <= 12'b111101111011;
   63595: result <= 12'b111101111010;
   63596: result <= 12'b111101111010;
   63597: result <= 12'b111101111010;
   63598: result <= 12'b111101111010;
   63599: result <= 12'b111101111010;
   63600: result <= 12'b111101111001;
   63601: result <= 12'b111101111001;
   63602: result <= 12'b111101111001;
   63603: result <= 12'b111101111001;
   63604: result <= 12'b111101111001;
   63605: result <= 12'b111101111000;
   63606: result <= 12'b111101111000;
   63607: result <= 12'b111101111000;
   63608: result <= 12'b111101111000;
   63609: result <= 12'b111101111000;
   63610: result <= 12'b111101111000;
   63611: result <= 12'b111101110111;
   63612: result <= 12'b111101110111;
   63613: result <= 12'b111101110111;
   63614: result <= 12'b111101110111;
   63615: result <= 12'b111101110111;
   63616: result <= 12'b111101110110;
   63617: result <= 12'b111101110110;
   63618: result <= 12'b111101110110;
   63619: result <= 12'b111101110110;
   63620: result <= 12'b111101110110;
   63621: result <= 12'b111101110101;
   63622: result <= 12'b111101110101;
   63623: result <= 12'b111101110101;
   63624: result <= 12'b111101110101;
   63625: result <= 12'b111101110101;
   63626: result <= 12'b111101110100;
   63627: result <= 12'b111101110100;
   63628: result <= 12'b111101110100;
   63629: result <= 12'b111101110100;
   63630: result <= 12'b111101110100;
   63631: result <= 12'b111101110011;
   63632: result <= 12'b111101110011;
   63633: result <= 12'b111101110011;
   63634: result <= 12'b111101110011;
   63635: result <= 12'b111101110011;
   63636: result <= 12'b111101110011;
   63637: result <= 12'b111101110010;
   63638: result <= 12'b111101110010;
   63639: result <= 12'b111101110010;
   63640: result <= 12'b111101110010;
   63641: result <= 12'b111101110010;
   63642: result <= 12'b111101110001;
   63643: result <= 12'b111101110001;
   63644: result <= 12'b111101110001;
   63645: result <= 12'b111101110001;
   63646: result <= 12'b111101110001;
   63647: result <= 12'b111101110000;
   63648: result <= 12'b111101110000;
   63649: result <= 12'b111101110000;
   63650: result <= 12'b111101110000;
   63651: result <= 12'b111101110000;
   63652: result <= 12'b111101101111;
   63653: result <= 12'b111101101111;
   63654: result <= 12'b111101101111;
   63655: result <= 12'b111101101111;
   63656: result <= 12'b111101101111;
   63657: result <= 12'b111101101110;
   63658: result <= 12'b111101101110;
   63659: result <= 12'b111101101110;
   63660: result <= 12'b111101101110;
   63661: result <= 12'b111101101110;
   63662: result <= 12'b111101101101;
   63663: result <= 12'b111101101101;
   63664: result <= 12'b111101101101;
   63665: result <= 12'b111101101101;
   63666: result <= 12'b111101101101;
   63667: result <= 12'b111101101101;
   63668: result <= 12'b111101101100;
   63669: result <= 12'b111101101100;
   63670: result <= 12'b111101101100;
   63671: result <= 12'b111101101100;
   63672: result <= 12'b111101101100;
   63673: result <= 12'b111101101011;
   63674: result <= 12'b111101101011;
   63675: result <= 12'b111101101011;
   63676: result <= 12'b111101101011;
   63677: result <= 12'b111101101011;
   63678: result <= 12'b111101101010;
   63679: result <= 12'b111101101010;
   63680: result <= 12'b111101101010;
   63681: result <= 12'b111101101010;
   63682: result <= 12'b111101101010;
   63683: result <= 12'b111101101001;
   63684: result <= 12'b111101101001;
   63685: result <= 12'b111101101001;
   63686: result <= 12'b111101101001;
   63687: result <= 12'b111101101001;
   63688: result <= 12'b111101101000;
   63689: result <= 12'b111101101000;
   63690: result <= 12'b111101101000;
   63691: result <= 12'b111101101000;
   63692: result <= 12'b111101101000;
   63693: result <= 12'b111101100111;
   63694: result <= 12'b111101100111;
   63695: result <= 12'b111101100111;
   63696: result <= 12'b111101100111;
   63697: result <= 12'b111101100111;
   63698: result <= 12'b111101100111;
   63699: result <= 12'b111101100110;
   63700: result <= 12'b111101100110;
   63701: result <= 12'b111101100110;
   63702: result <= 12'b111101100110;
   63703: result <= 12'b111101100110;
   63704: result <= 12'b111101100101;
   63705: result <= 12'b111101100101;
   63706: result <= 12'b111101100101;
   63707: result <= 12'b111101100101;
   63708: result <= 12'b111101100101;
   63709: result <= 12'b111101100100;
   63710: result <= 12'b111101100100;
   63711: result <= 12'b111101100100;
   63712: result <= 12'b111101100100;
   63713: result <= 12'b111101100100;
   63714: result <= 12'b111101100011;
   63715: result <= 12'b111101100011;
   63716: result <= 12'b111101100011;
   63717: result <= 12'b111101100011;
   63718: result <= 12'b111101100011;
   63719: result <= 12'b111101100010;
   63720: result <= 12'b111101100010;
   63721: result <= 12'b111101100010;
   63722: result <= 12'b111101100010;
   63723: result <= 12'b111101100010;
   63724: result <= 12'b111101100001;
   63725: result <= 12'b111101100001;
   63726: result <= 12'b111101100001;
   63727: result <= 12'b111101100001;
   63728: result <= 12'b111101100001;
   63729: result <= 12'b111101100001;
   63730: result <= 12'b111101100000;
   63731: result <= 12'b111101100000;
   63732: result <= 12'b111101100000;
   63733: result <= 12'b111101100000;
   63734: result <= 12'b111101100000;
   63735: result <= 12'b111101011111;
   63736: result <= 12'b111101011111;
   63737: result <= 12'b111101011111;
   63738: result <= 12'b111101011111;
   63739: result <= 12'b111101011111;
   63740: result <= 12'b111101011110;
   63741: result <= 12'b111101011110;
   63742: result <= 12'b111101011110;
   63743: result <= 12'b111101011110;
   63744: result <= 12'b111101011110;
   63745: result <= 12'b111101011101;
   63746: result <= 12'b111101011101;
   63747: result <= 12'b111101011101;
   63748: result <= 12'b111101011101;
   63749: result <= 12'b111101011101;
   63750: result <= 12'b111101011100;
   63751: result <= 12'b111101011100;
   63752: result <= 12'b111101011100;
   63753: result <= 12'b111101011100;
   63754: result <= 12'b111101011100;
   63755: result <= 12'b111101011100;
   63756: result <= 12'b111101011011;
   63757: result <= 12'b111101011011;
   63758: result <= 12'b111101011011;
   63759: result <= 12'b111101011011;
   63760: result <= 12'b111101011011;
   63761: result <= 12'b111101011010;
   63762: result <= 12'b111101011010;
   63763: result <= 12'b111101011010;
   63764: result <= 12'b111101011010;
   63765: result <= 12'b111101011010;
   63766: result <= 12'b111101011001;
   63767: result <= 12'b111101011001;
   63768: result <= 12'b111101011001;
   63769: result <= 12'b111101011001;
   63770: result <= 12'b111101011001;
   63771: result <= 12'b111101011000;
   63772: result <= 12'b111101011000;
   63773: result <= 12'b111101011000;
   63774: result <= 12'b111101011000;
   63775: result <= 12'b111101011000;
   63776: result <= 12'b111101010111;
   63777: result <= 12'b111101010111;
   63778: result <= 12'b111101010111;
   63779: result <= 12'b111101010111;
   63780: result <= 12'b111101010111;
   63781: result <= 12'b111101010110;
   63782: result <= 12'b111101010110;
   63783: result <= 12'b111101010110;
   63784: result <= 12'b111101010110;
   63785: result <= 12'b111101010110;
   63786: result <= 12'b111101010110;
   63787: result <= 12'b111101010101;
   63788: result <= 12'b111101010101;
   63789: result <= 12'b111101010101;
   63790: result <= 12'b111101010101;
   63791: result <= 12'b111101010101;
   63792: result <= 12'b111101010100;
   63793: result <= 12'b111101010100;
   63794: result <= 12'b111101010100;
   63795: result <= 12'b111101010100;
   63796: result <= 12'b111101010100;
   63797: result <= 12'b111101010011;
   63798: result <= 12'b111101010011;
   63799: result <= 12'b111101010011;
   63800: result <= 12'b111101010011;
   63801: result <= 12'b111101010011;
   63802: result <= 12'b111101010010;
   63803: result <= 12'b111101010010;
   63804: result <= 12'b111101010010;
   63805: result <= 12'b111101010010;
   63806: result <= 12'b111101010010;
   63807: result <= 12'b111101010001;
   63808: result <= 12'b111101010001;
   63809: result <= 12'b111101010001;
   63810: result <= 12'b111101010001;
   63811: result <= 12'b111101010001;
   63812: result <= 12'b111101010000;
   63813: result <= 12'b111101010000;
   63814: result <= 12'b111101010000;
   63815: result <= 12'b111101010000;
   63816: result <= 12'b111101010000;
   63817: result <= 12'b111101001111;
   63818: result <= 12'b111101001111;
   63819: result <= 12'b111101001111;
   63820: result <= 12'b111101001111;
   63821: result <= 12'b111101001111;
   63822: result <= 12'b111101001111;
   63823: result <= 12'b111101001110;
   63824: result <= 12'b111101001110;
   63825: result <= 12'b111101001110;
   63826: result <= 12'b111101001110;
   63827: result <= 12'b111101001110;
   63828: result <= 12'b111101001101;
   63829: result <= 12'b111101001101;
   63830: result <= 12'b111101001101;
   63831: result <= 12'b111101001101;
   63832: result <= 12'b111101001101;
   63833: result <= 12'b111101001100;
   63834: result <= 12'b111101001100;
   63835: result <= 12'b111101001100;
   63836: result <= 12'b111101001100;
   63837: result <= 12'b111101001100;
   63838: result <= 12'b111101001011;
   63839: result <= 12'b111101001011;
   63840: result <= 12'b111101001011;
   63841: result <= 12'b111101001011;
   63842: result <= 12'b111101001011;
   63843: result <= 12'b111101001010;
   63844: result <= 12'b111101001010;
   63845: result <= 12'b111101001010;
   63846: result <= 12'b111101001010;
   63847: result <= 12'b111101001010;
   63848: result <= 12'b111101001001;
   63849: result <= 12'b111101001001;
   63850: result <= 12'b111101001001;
   63851: result <= 12'b111101001001;
   63852: result <= 12'b111101001001;
   63853: result <= 12'b111101001001;
   63854: result <= 12'b111101001000;
   63855: result <= 12'b111101001000;
   63856: result <= 12'b111101001000;
   63857: result <= 12'b111101001000;
   63858: result <= 12'b111101001000;
   63859: result <= 12'b111101000111;
   63860: result <= 12'b111101000111;
   63861: result <= 12'b111101000111;
   63862: result <= 12'b111101000111;
   63863: result <= 12'b111101000111;
   63864: result <= 12'b111101000110;
   63865: result <= 12'b111101000110;
   63866: result <= 12'b111101000110;
   63867: result <= 12'b111101000110;
   63868: result <= 12'b111101000110;
   63869: result <= 12'b111101000101;
   63870: result <= 12'b111101000101;
   63871: result <= 12'b111101000101;
   63872: result <= 12'b111101000101;
   63873: result <= 12'b111101000101;
   63874: result <= 12'b111101000100;
   63875: result <= 12'b111101000100;
   63876: result <= 12'b111101000100;
   63877: result <= 12'b111101000100;
   63878: result <= 12'b111101000100;
   63879: result <= 12'b111101000011;
   63880: result <= 12'b111101000011;
   63881: result <= 12'b111101000011;
   63882: result <= 12'b111101000011;
   63883: result <= 12'b111101000011;
   63884: result <= 12'b111101000011;
   63885: result <= 12'b111101000010;
   63886: result <= 12'b111101000010;
   63887: result <= 12'b111101000010;
   63888: result <= 12'b111101000010;
   63889: result <= 12'b111101000010;
   63890: result <= 12'b111101000001;
   63891: result <= 12'b111101000001;
   63892: result <= 12'b111101000001;
   63893: result <= 12'b111101000001;
   63894: result <= 12'b111101000001;
   63895: result <= 12'b111101000000;
   63896: result <= 12'b111101000000;
   63897: result <= 12'b111101000000;
   63898: result <= 12'b111101000000;
   63899: result <= 12'b111101000000;
   63900: result <= 12'b111100111111;
   63901: result <= 12'b111100111111;
   63902: result <= 12'b111100111111;
   63903: result <= 12'b111100111111;
   63904: result <= 12'b111100111111;
   63905: result <= 12'b111100111110;
   63906: result <= 12'b111100111110;
   63907: result <= 12'b111100111110;
   63908: result <= 12'b111100111110;
   63909: result <= 12'b111100111110;
   63910: result <= 12'b111100111101;
   63911: result <= 12'b111100111101;
   63912: result <= 12'b111100111101;
   63913: result <= 12'b111100111101;
   63914: result <= 12'b111100111101;
   63915: result <= 12'b111100111101;
   63916: result <= 12'b111100111100;
   63917: result <= 12'b111100111100;
   63918: result <= 12'b111100111100;
   63919: result <= 12'b111100111100;
   63920: result <= 12'b111100111100;
   63921: result <= 12'b111100111011;
   63922: result <= 12'b111100111011;
   63923: result <= 12'b111100111011;
   63924: result <= 12'b111100111011;
   63925: result <= 12'b111100111011;
   63926: result <= 12'b111100111010;
   63927: result <= 12'b111100111010;
   63928: result <= 12'b111100111010;
   63929: result <= 12'b111100111010;
   63930: result <= 12'b111100111010;
   63931: result <= 12'b111100111001;
   63932: result <= 12'b111100111001;
   63933: result <= 12'b111100111001;
   63934: result <= 12'b111100111001;
   63935: result <= 12'b111100111001;
   63936: result <= 12'b111100111000;
   63937: result <= 12'b111100111000;
   63938: result <= 12'b111100111000;
   63939: result <= 12'b111100111000;
   63940: result <= 12'b111100111000;
   63941: result <= 12'b111100110111;
   63942: result <= 12'b111100110111;
   63943: result <= 12'b111100110111;
   63944: result <= 12'b111100110111;
   63945: result <= 12'b111100110111;
   63946: result <= 12'b111100110110;
   63947: result <= 12'b111100110110;
   63948: result <= 12'b111100110110;
   63949: result <= 12'b111100110110;
   63950: result <= 12'b111100110110;
   63951: result <= 12'b111100110110;
   63952: result <= 12'b111100110101;
   63953: result <= 12'b111100110101;
   63954: result <= 12'b111100110101;
   63955: result <= 12'b111100110101;
   63956: result <= 12'b111100110101;
   63957: result <= 12'b111100110100;
   63958: result <= 12'b111100110100;
   63959: result <= 12'b111100110100;
   63960: result <= 12'b111100110100;
   63961: result <= 12'b111100110100;
   63962: result <= 12'b111100110011;
   63963: result <= 12'b111100110011;
   63964: result <= 12'b111100110011;
   63965: result <= 12'b111100110011;
   63966: result <= 12'b111100110011;
   63967: result <= 12'b111100110010;
   63968: result <= 12'b111100110010;
   63969: result <= 12'b111100110010;
   63970: result <= 12'b111100110010;
   63971: result <= 12'b111100110010;
   63972: result <= 12'b111100110001;
   63973: result <= 12'b111100110001;
   63974: result <= 12'b111100110001;
   63975: result <= 12'b111100110001;
   63976: result <= 12'b111100110001;
   63977: result <= 12'b111100110000;
   63978: result <= 12'b111100110000;
   63979: result <= 12'b111100110000;
   63980: result <= 12'b111100110000;
   63981: result <= 12'b111100110000;
   63982: result <= 12'b111100101111;
   63983: result <= 12'b111100101111;
   63984: result <= 12'b111100101111;
   63985: result <= 12'b111100101111;
   63986: result <= 12'b111100101111;
   63987: result <= 12'b111100101111;
   63988: result <= 12'b111100101110;
   63989: result <= 12'b111100101110;
   63990: result <= 12'b111100101110;
   63991: result <= 12'b111100101110;
   63992: result <= 12'b111100101110;
   63993: result <= 12'b111100101101;
   63994: result <= 12'b111100101101;
   63995: result <= 12'b111100101101;
   63996: result <= 12'b111100101101;
   63997: result <= 12'b111100101101;
   63998: result <= 12'b111100101100;
   63999: result <= 12'b111100101100;
   64000: result <= 12'b111100101100;
   64001: result <= 12'b111100101100;
   64002: result <= 12'b111100101100;
   64003: result <= 12'b111100101011;
   64004: result <= 12'b111100101011;
   64005: result <= 12'b111100101011;
   64006: result <= 12'b111100101011;
   64007: result <= 12'b111100101011;
   64008: result <= 12'b111100101010;
   64009: result <= 12'b111100101010;
   64010: result <= 12'b111100101010;
   64011: result <= 12'b111100101010;
   64012: result <= 12'b111100101010;
   64013: result <= 12'b111100101001;
   64014: result <= 12'b111100101001;
   64015: result <= 12'b111100101001;
   64016: result <= 12'b111100101001;
   64017: result <= 12'b111100101001;
   64018: result <= 12'b111100101001;
   64019: result <= 12'b111100101000;
   64020: result <= 12'b111100101000;
   64021: result <= 12'b111100101000;
   64022: result <= 12'b111100101000;
   64023: result <= 12'b111100101000;
   64024: result <= 12'b111100100111;
   64025: result <= 12'b111100100111;
   64026: result <= 12'b111100100111;
   64027: result <= 12'b111100100111;
   64028: result <= 12'b111100100111;
   64029: result <= 12'b111100100110;
   64030: result <= 12'b111100100110;
   64031: result <= 12'b111100100110;
   64032: result <= 12'b111100100110;
   64033: result <= 12'b111100100110;
   64034: result <= 12'b111100100101;
   64035: result <= 12'b111100100101;
   64036: result <= 12'b111100100101;
   64037: result <= 12'b111100100101;
   64038: result <= 12'b111100100101;
   64039: result <= 12'b111100100100;
   64040: result <= 12'b111100100100;
   64041: result <= 12'b111100100100;
   64042: result <= 12'b111100100100;
   64043: result <= 12'b111100100100;
   64044: result <= 12'b111100100011;
   64045: result <= 12'b111100100011;
   64046: result <= 12'b111100100011;
   64047: result <= 12'b111100100011;
   64048: result <= 12'b111100100011;
   64049: result <= 12'b111100100010;
   64050: result <= 12'b111100100010;
   64051: result <= 12'b111100100010;
   64052: result <= 12'b111100100010;
   64053: result <= 12'b111100100010;
   64054: result <= 12'b111100100010;
   64055: result <= 12'b111100100001;
   64056: result <= 12'b111100100001;
   64057: result <= 12'b111100100001;
   64058: result <= 12'b111100100001;
   64059: result <= 12'b111100100001;
   64060: result <= 12'b111100100000;
   64061: result <= 12'b111100100000;
   64062: result <= 12'b111100100000;
   64063: result <= 12'b111100100000;
   64064: result <= 12'b111100100000;
   64065: result <= 12'b111100011111;
   64066: result <= 12'b111100011111;
   64067: result <= 12'b111100011111;
   64068: result <= 12'b111100011111;
   64069: result <= 12'b111100011111;
   64070: result <= 12'b111100011110;
   64071: result <= 12'b111100011110;
   64072: result <= 12'b111100011110;
   64073: result <= 12'b111100011110;
   64074: result <= 12'b111100011110;
   64075: result <= 12'b111100011101;
   64076: result <= 12'b111100011101;
   64077: result <= 12'b111100011101;
   64078: result <= 12'b111100011101;
   64079: result <= 12'b111100011101;
   64080: result <= 12'b111100011100;
   64081: result <= 12'b111100011100;
   64082: result <= 12'b111100011100;
   64083: result <= 12'b111100011100;
   64084: result <= 12'b111100011100;
   64085: result <= 12'b111100011011;
   64086: result <= 12'b111100011011;
   64087: result <= 12'b111100011011;
   64088: result <= 12'b111100011011;
   64089: result <= 12'b111100011011;
   64090: result <= 12'b111100011011;
   64091: result <= 12'b111100011010;
   64092: result <= 12'b111100011010;
   64093: result <= 12'b111100011010;
   64094: result <= 12'b111100011010;
   64095: result <= 12'b111100011010;
   64096: result <= 12'b111100011001;
   64097: result <= 12'b111100011001;
   64098: result <= 12'b111100011001;
   64099: result <= 12'b111100011001;
   64100: result <= 12'b111100011001;
   64101: result <= 12'b111100011000;
   64102: result <= 12'b111100011000;
   64103: result <= 12'b111100011000;
   64104: result <= 12'b111100011000;
   64105: result <= 12'b111100011000;
   64106: result <= 12'b111100010111;
   64107: result <= 12'b111100010111;
   64108: result <= 12'b111100010111;
   64109: result <= 12'b111100010111;
   64110: result <= 12'b111100010111;
   64111: result <= 12'b111100010110;
   64112: result <= 12'b111100010110;
   64113: result <= 12'b111100010110;
   64114: result <= 12'b111100010110;
   64115: result <= 12'b111100010110;
   64116: result <= 12'b111100010101;
   64117: result <= 12'b111100010101;
   64118: result <= 12'b111100010101;
   64119: result <= 12'b111100010101;
   64120: result <= 12'b111100010101;
   64121: result <= 12'b111100010100;
   64122: result <= 12'b111100010100;
   64123: result <= 12'b111100010100;
   64124: result <= 12'b111100010100;
   64125: result <= 12'b111100010100;
   64126: result <= 12'b111100010100;
   64127: result <= 12'b111100010011;
   64128: result <= 12'b111100010011;
   64129: result <= 12'b111100010011;
   64130: result <= 12'b111100010011;
   64131: result <= 12'b111100010011;
   64132: result <= 12'b111100010010;
   64133: result <= 12'b111100010010;
   64134: result <= 12'b111100010010;
   64135: result <= 12'b111100010010;
   64136: result <= 12'b111100010010;
   64137: result <= 12'b111100010001;
   64138: result <= 12'b111100010001;
   64139: result <= 12'b111100010001;
   64140: result <= 12'b111100010001;
   64141: result <= 12'b111100010001;
   64142: result <= 12'b111100010000;
   64143: result <= 12'b111100010000;
   64144: result <= 12'b111100010000;
   64145: result <= 12'b111100010000;
   64146: result <= 12'b111100010000;
   64147: result <= 12'b111100001111;
   64148: result <= 12'b111100001111;
   64149: result <= 12'b111100001111;
   64150: result <= 12'b111100001111;
   64151: result <= 12'b111100001111;
   64152: result <= 12'b111100001110;
   64153: result <= 12'b111100001110;
   64154: result <= 12'b111100001110;
   64155: result <= 12'b111100001110;
   64156: result <= 12'b111100001110;
   64157: result <= 12'b111100001101;
   64158: result <= 12'b111100001101;
   64159: result <= 12'b111100001101;
   64160: result <= 12'b111100001101;
   64161: result <= 12'b111100001101;
   64162: result <= 12'b111100001101;
   64163: result <= 12'b111100001100;
   64164: result <= 12'b111100001100;
   64165: result <= 12'b111100001100;
   64166: result <= 12'b111100001100;
   64167: result <= 12'b111100001100;
   64168: result <= 12'b111100001011;
   64169: result <= 12'b111100001011;
   64170: result <= 12'b111100001011;
   64171: result <= 12'b111100001011;
   64172: result <= 12'b111100001011;
   64173: result <= 12'b111100001010;
   64174: result <= 12'b111100001010;
   64175: result <= 12'b111100001010;
   64176: result <= 12'b111100001010;
   64177: result <= 12'b111100001010;
   64178: result <= 12'b111100001001;
   64179: result <= 12'b111100001001;
   64180: result <= 12'b111100001001;
   64181: result <= 12'b111100001001;
   64182: result <= 12'b111100001001;
   64183: result <= 12'b111100001000;
   64184: result <= 12'b111100001000;
   64185: result <= 12'b111100001000;
   64186: result <= 12'b111100001000;
   64187: result <= 12'b111100001000;
   64188: result <= 12'b111100000111;
   64189: result <= 12'b111100000111;
   64190: result <= 12'b111100000111;
   64191: result <= 12'b111100000111;
   64192: result <= 12'b111100000111;
   64193: result <= 12'b111100000110;
   64194: result <= 12'b111100000110;
   64195: result <= 12'b111100000110;
   64196: result <= 12'b111100000110;
   64197: result <= 12'b111100000110;
   64198: result <= 12'b111100000101;
   64199: result <= 12'b111100000101;
   64200: result <= 12'b111100000101;
   64201: result <= 12'b111100000101;
   64202: result <= 12'b111100000101;
   64203: result <= 12'b111100000101;
   64204: result <= 12'b111100000100;
   64205: result <= 12'b111100000100;
   64206: result <= 12'b111100000100;
   64207: result <= 12'b111100000100;
   64208: result <= 12'b111100000100;
   64209: result <= 12'b111100000011;
   64210: result <= 12'b111100000011;
   64211: result <= 12'b111100000011;
   64212: result <= 12'b111100000011;
   64213: result <= 12'b111100000011;
   64214: result <= 12'b111100000010;
   64215: result <= 12'b111100000010;
   64216: result <= 12'b111100000010;
   64217: result <= 12'b111100000010;
   64218: result <= 12'b111100000010;
   64219: result <= 12'b111100000001;
   64220: result <= 12'b111100000001;
   64221: result <= 12'b111100000001;
   64222: result <= 12'b111100000001;
   64223: result <= 12'b111100000001;
   64224: result <= 12'b111100000000;
   64225: result <= 12'b111100000000;
   64226: result <= 12'b111100000000;
   64227: result <= 12'b111100000000;
   64228: result <= 12'b111100000000;
   64229: result <= 12'b111111111111;
   64230: result <= 12'b111111111111;
   64231: result <= 12'b111111111111;
   64232: result <= 12'b111111111111;
   64233: result <= 12'b111111111111;
   64234: result <= 12'b111111111110;
   64235: result <= 12'b111111111110;
   64236: result <= 12'b111111111110;
   64237: result <= 12'b111111111110;
   64238: result <= 12'b111111111110;
   64239: result <= 12'b111111111110;
   64240: result <= 12'b111111111101;
   64241: result <= 12'b111111111101;
   64242: result <= 12'b111111111101;
   64243: result <= 12'b111111111101;
   64244: result <= 12'b111111111101;
   64245: result <= 12'b111111111100;
   64246: result <= 12'b111111111100;
   64247: result <= 12'b111111111100;
   64248: result <= 12'b111111111100;
   64249: result <= 12'b111111111100;
   64250: result <= 12'b111111111011;
   64251: result <= 12'b111111111011;
   64252: result <= 12'b111111111011;
   64253: result <= 12'b111111111011;
   64254: result <= 12'b111111111011;
   64255: result <= 12'b111111111010;
   64256: result <= 12'b111111111010;
   64257: result <= 12'b111111111010;
   64258: result <= 12'b111111111010;
   64259: result <= 12'b111111111010;
   64260: result <= 12'b111111111001;
   64261: result <= 12'b111111111001;
   64262: result <= 12'b111111111001;
   64263: result <= 12'b111111111001;
   64264: result <= 12'b111111111001;
   64265: result <= 12'b111111111000;
   64266: result <= 12'b111111111000;
   64267: result <= 12'b111111111000;
   64268: result <= 12'b111111111000;
   64269: result <= 12'b111111111000;
   64270: result <= 12'b111111110111;
   64271: result <= 12'b111111110111;
   64272: result <= 12'b111111110111;
   64273: result <= 12'b111111110111;
   64274: result <= 12'b111111110111;
   64275: result <= 12'b111111110110;
   64276: result <= 12'b111111110110;
   64277: result <= 12'b111111110110;
   64278: result <= 12'b111111110110;
   64279: result <= 12'b111111110110;
   64280: result <= 12'b111111110110;
   64281: result <= 12'b111111110101;
   64282: result <= 12'b111111110101;
   64283: result <= 12'b111111110101;
   64284: result <= 12'b111111110101;
   64285: result <= 12'b111111110101;
   64286: result <= 12'b111111110100;
   64287: result <= 12'b111111110100;
   64288: result <= 12'b111111110100;
   64289: result <= 12'b111111110100;
   64290: result <= 12'b111111110100;
   64291: result <= 12'b111111110011;
   64292: result <= 12'b111111110011;
   64293: result <= 12'b111111110011;
   64294: result <= 12'b111111110011;
   64295: result <= 12'b111111110011;
   64296: result <= 12'b111111110010;
   64297: result <= 12'b111111110010;
   64298: result <= 12'b111111110010;
   64299: result <= 12'b111111110010;
   64300: result <= 12'b111111110010;
   64301: result <= 12'b111111110001;
   64302: result <= 12'b111111110001;
   64303: result <= 12'b111111110001;
   64304: result <= 12'b111111110001;
   64305: result <= 12'b111111110001;
   64306: result <= 12'b111111110000;
   64307: result <= 12'b111111110000;
   64308: result <= 12'b111111110000;
   64309: result <= 12'b111111110000;
   64310: result <= 12'b111111110000;
   64311: result <= 12'b111111101111;
   64312: result <= 12'b111111101111;
   64313: result <= 12'b111111101111;
   64314: result <= 12'b111111101111;
   64315: result <= 12'b111111101111;
   64316: result <= 12'b111111101111;
   64317: result <= 12'b111111101110;
   64318: result <= 12'b111111101110;
   64319: result <= 12'b111111101110;
   64320: result <= 12'b111111101110;
   64321: result <= 12'b111111101110;
   64322: result <= 12'b111111101101;
   64323: result <= 12'b111111101101;
   64324: result <= 12'b111111101101;
   64325: result <= 12'b111111101101;
   64326: result <= 12'b111111101101;
   64327: result <= 12'b111111101100;
   64328: result <= 12'b111111101100;
   64329: result <= 12'b111111101100;
   64330: result <= 12'b111111101100;
   64331: result <= 12'b111111101100;
   64332: result <= 12'b111111101011;
   64333: result <= 12'b111111101011;
   64334: result <= 12'b111111101011;
   64335: result <= 12'b111111101011;
   64336: result <= 12'b111111101011;
   64337: result <= 12'b111111101010;
   64338: result <= 12'b111111101010;
   64339: result <= 12'b111111101010;
   64340: result <= 12'b111111101010;
   64341: result <= 12'b111111101010;
   64342: result <= 12'b111111101001;
   64343: result <= 12'b111111101001;
   64344: result <= 12'b111111101001;
   64345: result <= 12'b111111101001;
   64346: result <= 12'b111111101001;
   64347: result <= 12'b111111101000;
   64348: result <= 12'b111111101000;
   64349: result <= 12'b111111101000;
   64350: result <= 12'b111111101000;
   64351: result <= 12'b111111101000;
   64352: result <= 12'b111111100111;
   64353: result <= 12'b111111100111;
   64354: result <= 12'b111111100111;
   64355: result <= 12'b111111100111;
   64356: result <= 12'b111111100111;
   64357: result <= 12'b111111100111;
   64358: result <= 12'b111111100110;
   64359: result <= 12'b111111100110;
   64360: result <= 12'b111111100110;
   64361: result <= 12'b111111100110;
   64362: result <= 12'b111111100110;
   64363: result <= 12'b111111100101;
   64364: result <= 12'b111111100101;
   64365: result <= 12'b111111100101;
   64366: result <= 12'b111111100101;
   64367: result <= 12'b111111100101;
   64368: result <= 12'b111111100100;
   64369: result <= 12'b111111100100;
   64370: result <= 12'b111111100100;
   64371: result <= 12'b111111100100;
   64372: result <= 12'b111111100100;
   64373: result <= 12'b111111100011;
   64374: result <= 12'b111111100011;
   64375: result <= 12'b111111100011;
   64376: result <= 12'b111111100011;
   64377: result <= 12'b111111100011;
   64378: result <= 12'b111111100010;
   64379: result <= 12'b111111100010;
   64380: result <= 12'b111111100010;
   64381: result <= 12'b111111100010;
   64382: result <= 12'b111111100010;
   64383: result <= 12'b111111100001;
   64384: result <= 12'b111111100001;
   64385: result <= 12'b111111100001;
   64386: result <= 12'b111111100001;
   64387: result <= 12'b111111100001;
   64388: result <= 12'b111111100000;
   64389: result <= 12'b111111100000;
   64390: result <= 12'b111111100000;
   64391: result <= 12'b111111100000;
   64392: result <= 12'b111111100000;
   64393: result <= 12'b111111011111;
   64394: result <= 12'b111111011111;
   64395: result <= 12'b111111011111;
   64396: result <= 12'b111111011111;
   64397: result <= 12'b111111011111;
   64398: result <= 12'b111111011111;
   64399: result <= 12'b111111011110;
   64400: result <= 12'b111111011110;
   64401: result <= 12'b111111011110;
   64402: result <= 12'b111111011110;
   64403: result <= 12'b111111011110;
   64404: result <= 12'b111111011101;
   64405: result <= 12'b111111011101;
   64406: result <= 12'b111111011101;
   64407: result <= 12'b111111011101;
   64408: result <= 12'b111111011101;
   64409: result <= 12'b111111011100;
   64410: result <= 12'b111111011100;
   64411: result <= 12'b111111011100;
   64412: result <= 12'b111111011100;
   64413: result <= 12'b111111011100;
   64414: result <= 12'b111111011011;
   64415: result <= 12'b111111011011;
   64416: result <= 12'b111111011011;
   64417: result <= 12'b111111011011;
   64418: result <= 12'b111111011011;
   64419: result <= 12'b111111011010;
   64420: result <= 12'b111111011010;
   64421: result <= 12'b111111011010;
   64422: result <= 12'b111111011010;
   64423: result <= 12'b111111011010;
   64424: result <= 12'b111111011001;
   64425: result <= 12'b111111011001;
   64426: result <= 12'b111111011001;
   64427: result <= 12'b111111011001;
   64428: result <= 12'b111111011001;
   64429: result <= 12'b111111011000;
   64430: result <= 12'b111111011000;
   64431: result <= 12'b111111011000;
   64432: result <= 12'b111111011000;
   64433: result <= 12'b111111011000;
   64434: result <= 12'b111111010111;
   64435: result <= 12'b111111010111;
   64436: result <= 12'b111111010111;
   64437: result <= 12'b111111010111;
   64438: result <= 12'b111111010111;
   64439: result <= 12'b111111010110;
   64440: result <= 12'b111111010110;
   64441: result <= 12'b111111010110;
   64442: result <= 12'b111111010110;
   64443: result <= 12'b111111010110;
   64444: result <= 12'b111111010110;
   64445: result <= 12'b111111010101;
   64446: result <= 12'b111111010101;
   64447: result <= 12'b111111010101;
   64448: result <= 12'b111111010101;
   64449: result <= 12'b111111010101;
   64450: result <= 12'b111111010100;
   64451: result <= 12'b111111010100;
   64452: result <= 12'b111111010100;
   64453: result <= 12'b111111010100;
   64454: result <= 12'b111111010100;
   64455: result <= 12'b111111010011;
   64456: result <= 12'b111111010011;
   64457: result <= 12'b111111010011;
   64458: result <= 12'b111111010011;
   64459: result <= 12'b111111010011;
   64460: result <= 12'b111111010010;
   64461: result <= 12'b111111010010;
   64462: result <= 12'b111111010010;
   64463: result <= 12'b111111010010;
   64464: result <= 12'b111111010010;
   64465: result <= 12'b111111010001;
   64466: result <= 12'b111111010001;
   64467: result <= 12'b111111010001;
   64468: result <= 12'b111111010001;
   64469: result <= 12'b111111010001;
   64470: result <= 12'b111111010000;
   64471: result <= 12'b111111010000;
   64472: result <= 12'b111111010000;
   64473: result <= 12'b111111010000;
   64474: result <= 12'b111111010000;
   64475: result <= 12'b111111001111;
   64476: result <= 12'b111111001111;
   64477: result <= 12'b111111001111;
   64478: result <= 12'b111111001111;
   64479: result <= 12'b111111001111;
   64480: result <= 12'b111111001110;
   64481: result <= 12'b111111001110;
   64482: result <= 12'b111111001110;
   64483: result <= 12'b111111001110;
   64484: result <= 12'b111111001110;
   64485: result <= 12'b111111001110;
   64486: result <= 12'b111111001101;
   64487: result <= 12'b111111001101;
   64488: result <= 12'b111111001101;
   64489: result <= 12'b111111001101;
   64490: result <= 12'b111111001101;
   64491: result <= 12'b111111001100;
   64492: result <= 12'b111111001100;
   64493: result <= 12'b111111001100;
   64494: result <= 12'b111111001100;
   64495: result <= 12'b111111001100;
   64496: result <= 12'b111111001011;
   64497: result <= 12'b111111001011;
   64498: result <= 12'b111111001011;
   64499: result <= 12'b111111001011;
   64500: result <= 12'b111111001011;
   64501: result <= 12'b111111001010;
   64502: result <= 12'b111111001010;
   64503: result <= 12'b111111001010;
   64504: result <= 12'b111111001010;
   64505: result <= 12'b111111001010;
   64506: result <= 12'b111111001001;
   64507: result <= 12'b111111001001;
   64508: result <= 12'b111111001001;
   64509: result <= 12'b111111001001;
   64510: result <= 12'b111111001001;
   64511: result <= 12'b111111001000;
   64512: result <= 12'b111111001000;
   64513: result <= 12'b111111001000;
   64514: result <= 12'b111111001000;
   64515: result <= 12'b111111001000;
   64516: result <= 12'b111111000111;
   64517: result <= 12'b111111000111;
   64518: result <= 12'b111111000111;
   64519: result <= 12'b111111000111;
   64520: result <= 12'b111111000111;
   64521: result <= 12'b111111000110;
   64522: result <= 12'b111111000110;
   64523: result <= 12'b111111000110;
   64524: result <= 12'b111111000110;
   64525: result <= 12'b111111000110;
   64526: result <= 12'b111111000110;
   64527: result <= 12'b111111000101;
   64528: result <= 12'b111111000101;
   64529: result <= 12'b111111000101;
   64530: result <= 12'b111111000101;
   64531: result <= 12'b111111000101;
   64532: result <= 12'b111111000100;
   64533: result <= 12'b111111000100;
   64534: result <= 12'b111111000100;
   64535: result <= 12'b111111000100;
   64536: result <= 12'b111111000100;
   64537: result <= 12'b111111000011;
   64538: result <= 12'b111111000011;
   64539: result <= 12'b111111000011;
   64540: result <= 12'b111111000011;
   64541: result <= 12'b111111000011;
   64542: result <= 12'b111111000010;
   64543: result <= 12'b111111000010;
   64544: result <= 12'b111111000010;
   64545: result <= 12'b111111000010;
   64546: result <= 12'b111111000010;
   64547: result <= 12'b111111000001;
   64548: result <= 12'b111111000001;
   64549: result <= 12'b111111000001;
   64550: result <= 12'b111111000001;
   64551: result <= 12'b111111000001;
   64552: result <= 12'b111111000000;
   64553: result <= 12'b111111000000;
   64554: result <= 12'b111111000000;
   64555: result <= 12'b111111000000;
   64556: result <= 12'b111111000000;
   64557: result <= 12'b111110111111;
   64558: result <= 12'b111110111111;
   64559: result <= 12'b111110111111;
   64560: result <= 12'b111110111111;
   64561: result <= 12'b111110111111;
   64562: result <= 12'b111110111110;
   64563: result <= 12'b111110111110;
   64564: result <= 12'b111110111110;
   64565: result <= 12'b111110111110;
   64566: result <= 12'b111110111110;
   64567: result <= 12'b111110111101;
   64568: result <= 12'b111110111101;
   64569: result <= 12'b111110111101;
   64570: result <= 12'b111110111101;
   64571: result <= 12'b111110111101;
   64572: result <= 12'b111110111101;
   64573: result <= 12'b111110111100;
   64574: result <= 12'b111110111100;
   64575: result <= 12'b111110111100;
   64576: result <= 12'b111110111100;
   64577: result <= 12'b111110111100;
   64578: result <= 12'b111110111011;
   64579: result <= 12'b111110111011;
   64580: result <= 12'b111110111011;
   64581: result <= 12'b111110111011;
   64582: result <= 12'b111110111011;
   64583: result <= 12'b111110111010;
   64584: result <= 12'b111110111010;
   64585: result <= 12'b111110111010;
   64586: result <= 12'b111110111010;
   64587: result <= 12'b111110111010;
   64588: result <= 12'b111110111001;
   64589: result <= 12'b111110111001;
   64590: result <= 12'b111110111001;
   64591: result <= 12'b111110111001;
   64592: result <= 12'b111110111001;
   64593: result <= 12'b111110111000;
   64594: result <= 12'b111110111000;
   64595: result <= 12'b111110111000;
   64596: result <= 12'b111110111000;
   64597: result <= 12'b111110111000;
   64598: result <= 12'b111110110111;
   64599: result <= 12'b111110110111;
   64600: result <= 12'b111110110111;
   64601: result <= 12'b111110110111;
   64602: result <= 12'b111110110111;
   64603: result <= 12'b111110110110;
   64604: result <= 12'b111110110110;
   64605: result <= 12'b111110110110;
   64606: result <= 12'b111110110110;
   64607: result <= 12'b111110110110;
   64608: result <= 12'b111110110101;
   64609: result <= 12'b111110110101;
   64610: result <= 12'b111110110101;
   64611: result <= 12'b111110110101;
   64612: result <= 12'b111110110101;
   64613: result <= 12'b111110110100;
   64614: result <= 12'b111110110100;
   64615: result <= 12'b111110110100;
   64616: result <= 12'b111110110100;
   64617: result <= 12'b111110110100;
   64618: result <= 12'b111110110100;
   64619: result <= 12'b111110110011;
   64620: result <= 12'b111110110011;
   64621: result <= 12'b111110110011;
   64622: result <= 12'b111110110011;
   64623: result <= 12'b111110110011;
   64624: result <= 12'b111110110010;
   64625: result <= 12'b111110110010;
   64626: result <= 12'b111110110010;
   64627: result <= 12'b111110110010;
   64628: result <= 12'b111110110010;
   64629: result <= 12'b111110110001;
   64630: result <= 12'b111110110001;
   64631: result <= 12'b111110110001;
   64632: result <= 12'b111110110001;
   64633: result <= 12'b111110110001;
   64634: result <= 12'b111110110000;
   64635: result <= 12'b111110110000;
   64636: result <= 12'b111110110000;
   64637: result <= 12'b111110110000;
   64638: result <= 12'b111110110000;
   64639: result <= 12'b111110101111;
   64640: result <= 12'b111110101111;
   64641: result <= 12'b111110101111;
   64642: result <= 12'b111110101111;
   64643: result <= 12'b111110101111;
   64644: result <= 12'b111110101110;
   64645: result <= 12'b111110101110;
   64646: result <= 12'b111110101110;
   64647: result <= 12'b111110101110;
   64648: result <= 12'b111110101110;
   64649: result <= 12'b111110101101;
   64650: result <= 12'b111110101101;
   64651: result <= 12'b111110101101;
   64652: result <= 12'b111110101101;
   64653: result <= 12'b111110101101;
   64654: result <= 12'b111110101100;
   64655: result <= 12'b111110101100;
   64656: result <= 12'b111110101100;
   64657: result <= 12'b111110101100;
   64658: result <= 12'b111110101100;
   64659: result <= 12'b111110101011;
   64660: result <= 12'b111110101011;
   64661: result <= 12'b111110101011;
   64662: result <= 12'b111110101011;
   64663: result <= 12'b111110101011;
   64664: result <= 12'b111110101011;
   64665: result <= 12'b111110101010;
   64666: result <= 12'b111110101010;
   64667: result <= 12'b111110101010;
   64668: result <= 12'b111110101010;
   64669: result <= 12'b111110101010;
   64670: result <= 12'b111110101001;
   64671: result <= 12'b111110101001;
   64672: result <= 12'b111110101001;
   64673: result <= 12'b111110101001;
   64674: result <= 12'b111110101001;
   64675: result <= 12'b111110101000;
   64676: result <= 12'b111110101000;
   64677: result <= 12'b111110101000;
   64678: result <= 12'b111110101000;
   64679: result <= 12'b111110101000;
   64680: result <= 12'b111110100111;
   64681: result <= 12'b111110100111;
   64682: result <= 12'b111110100111;
   64683: result <= 12'b111110100111;
   64684: result <= 12'b111110100111;
   64685: result <= 12'b111110100110;
   64686: result <= 12'b111110100110;
   64687: result <= 12'b111110100110;
   64688: result <= 12'b111110100110;
   64689: result <= 12'b111110100110;
   64690: result <= 12'b111110100101;
   64691: result <= 12'b111110100101;
   64692: result <= 12'b111110100101;
   64693: result <= 12'b111110100101;
   64694: result <= 12'b111110100101;
   64695: result <= 12'b111110100100;
   64696: result <= 12'b111110100100;
   64697: result <= 12'b111110100100;
   64698: result <= 12'b111110100100;
   64699: result <= 12'b111110100100;
   64700: result <= 12'b111110100011;
   64701: result <= 12'b111110100011;
   64702: result <= 12'b111110100011;
   64703: result <= 12'b111110100011;
   64704: result <= 12'b111110100011;
   64705: result <= 12'b111110100010;
   64706: result <= 12'b111110100010;
   64707: result <= 12'b111110100010;
   64708: result <= 12'b111110100010;
   64709: result <= 12'b111110100010;
   64710: result <= 12'b111110100010;
   64711: result <= 12'b111110100001;
   64712: result <= 12'b111110100001;
   64713: result <= 12'b111110100001;
   64714: result <= 12'b111110100001;
   64715: result <= 12'b111110100001;
   64716: result <= 12'b111110100000;
   64717: result <= 12'b111110100000;
   64718: result <= 12'b111110100000;
   64719: result <= 12'b111110100000;
   64720: result <= 12'b111110100000;
   64721: result <= 12'b111110011111;
   64722: result <= 12'b111110011111;
   64723: result <= 12'b111110011111;
   64724: result <= 12'b111110011111;
   64725: result <= 12'b111110011111;
   64726: result <= 12'b111110011110;
   64727: result <= 12'b111110011110;
   64728: result <= 12'b111110011110;
   64729: result <= 12'b111110011110;
   64730: result <= 12'b111110011110;
   64731: result <= 12'b111110011101;
   64732: result <= 12'b111110011101;
   64733: result <= 12'b111110011101;
   64734: result <= 12'b111110011101;
   64735: result <= 12'b111110011101;
   64736: result <= 12'b111110011100;
   64737: result <= 12'b111110011100;
   64738: result <= 12'b111110011100;
   64739: result <= 12'b111110011100;
   64740: result <= 12'b111110011100;
   64741: result <= 12'b111110011011;
   64742: result <= 12'b111110011011;
   64743: result <= 12'b111110011011;
   64744: result <= 12'b111110011011;
   64745: result <= 12'b111110011011;
   64746: result <= 12'b111110011010;
   64747: result <= 12'b111110011010;
   64748: result <= 12'b111110011010;
   64749: result <= 12'b111110011010;
   64750: result <= 12'b111110011010;
   64751: result <= 12'b111110011001;
   64752: result <= 12'b111110011001;
   64753: result <= 12'b111110011001;
   64754: result <= 12'b111110011001;
   64755: result <= 12'b111110011001;
   64756: result <= 12'b111110011001;
   64757: result <= 12'b111110011000;
   64758: result <= 12'b111110011000;
   64759: result <= 12'b111110011000;
   64760: result <= 12'b111110011000;
   64761: result <= 12'b111110011000;
   64762: result <= 12'b111110010111;
   64763: result <= 12'b111110010111;
   64764: result <= 12'b111110010111;
   64765: result <= 12'b111110010111;
   64766: result <= 12'b111110010111;
   64767: result <= 12'b111110010110;
   64768: result <= 12'b111110010110;
   64769: result <= 12'b111110010110;
   64770: result <= 12'b111110010110;
   64771: result <= 12'b111110010110;
   64772: result <= 12'b111110010101;
   64773: result <= 12'b111110010101;
   64774: result <= 12'b111110010101;
   64775: result <= 12'b111110010101;
   64776: result <= 12'b111110010101;
   64777: result <= 12'b111110010100;
   64778: result <= 12'b111110010100;
   64779: result <= 12'b111110010100;
   64780: result <= 12'b111110010100;
   64781: result <= 12'b111110010100;
   64782: result <= 12'b111110010011;
   64783: result <= 12'b111110010011;
   64784: result <= 12'b111110010011;
   64785: result <= 12'b111110010011;
   64786: result <= 12'b111110010011;
   64787: result <= 12'b111110010010;
   64788: result <= 12'b111110010010;
   64789: result <= 12'b111110010010;
   64790: result <= 12'b111110010010;
   64791: result <= 12'b111110010010;
   64792: result <= 12'b111110010001;
   64793: result <= 12'b111110010001;
   64794: result <= 12'b111110010001;
   64795: result <= 12'b111110010001;
   64796: result <= 12'b111110010001;
   64797: result <= 12'b111110010000;
   64798: result <= 12'b111110010000;
   64799: result <= 12'b111110010000;
   64800: result <= 12'b111110010000;
   64801: result <= 12'b111110010000;
   64802: result <= 12'b111110010000;
   64803: result <= 12'b111110001111;
   64804: result <= 12'b111110001111;
   64805: result <= 12'b111110001111;
   64806: result <= 12'b111110001111;
   64807: result <= 12'b111110001111;
   64808: result <= 12'b111110001110;
   64809: result <= 12'b111110001110;
   64810: result <= 12'b111110001110;
   64811: result <= 12'b111110001110;
   64812: result <= 12'b111110001110;
   64813: result <= 12'b111110001101;
   64814: result <= 12'b111110001101;
   64815: result <= 12'b111110001101;
   64816: result <= 12'b111110001101;
   64817: result <= 12'b111110001101;
   64818: result <= 12'b111110001100;
   64819: result <= 12'b111110001100;
   64820: result <= 12'b111110001100;
   64821: result <= 12'b111110001100;
   64822: result <= 12'b111110001100;
   64823: result <= 12'b111110001011;
   64824: result <= 12'b111110001011;
   64825: result <= 12'b111110001011;
   64826: result <= 12'b111110001011;
   64827: result <= 12'b111110001011;
   64828: result <= 12'b111110001010;
   64829: result <= 12'b111110001010;
   64830: result <= 12'b111110001010;
   64831: result <= 12'b111110001010;
   64832: result <= 12'b111110001010;
   64833: result <= 12'b111110001001;
   64834: result <= 12'b111110001001;
   64835: result <= 12'b111110001001;
   64836: result <= 12'b111110001001;
   64837: result <= 12'b111110001001;
   64838: result <= 12'b111110001000;
   64839: result <= 12'b111110001000;
   64840: result <= 12'b111110001000;
   64841: result <= 12'b111110001000;
   64842: result <= 12'b111110001000;
   64843: result <= 12'b111110000111;
   64844: result <= 12'b111110000111;
   64845: result <= 12'b111110000111;
   64846: result <= 12'b111110000111;
   64847: result <= 12'b111110000111;
   64848: result <= 12'b111110000110;
   64849: result <= 12'b111110000110;
   64850: result <= 12'b111110000110;
   64851: result <= 12'b111110000110;
   64852: result <= 12'b111110000110;
   64853: result <= 12'b111110000110;
   64854: result <= 12'b111110000101;
   64855: result <= 12'b111110000101;
   64856: result <= 12'b111110000101;
   64857: result <= 12'b111110000101;
   64858: result <= 12'b111110000101;
   64859: result <= 12'b111110000100;
   64860: result <= 12'b111110000100;
   64861: result <= 12'b111110000100;
   64862: result <= 12'b111110000100;
   64863: result <= 12'b111110000100;
   64864: result <= 12'b111110000011;
   64865: result <= 12'b111110000011;
   64866: result <= 12'b111110000011;
   64867: result <= 12'b111110000011;
   64868: result <= 12'b111110000011;
   64869: result <= 12'b111110000010;
   64870: result <= 12'b111110000010;
   64871: result <= 12'b111110000010;
   64872: result <= 12'b111110000010;
   64873: result <= 12'b111110000010;
   64874: result <= 12'b111110000001;
   64875: result <= 12'b111110000001;
   64876: result <= 12'b111110000001;
   64877: result <= 12'b111110000001;
   64878: result <= 12'b111110000001;
   64879: result <= 12'b111110000000;
   64880: result <= 12'b111110000000;
   64881: result <= 12'b111110000000;
   64882: result <= 12'b111110000000;
   64883: result <= 12'b111110000000;
   64884: result <= 12'b111111111111;
   64885: result <= 12'b111111111111;
   64886: result <= 12'b111111111111;
   64887: result <= 12'b111111111111;
   64888: result <= 12'b111111111111;
   64889: result <= 12'b111111111110;
   64890: result <= 12'b111111111110;
   64891: result <= 12'b111111111110;
   64892: result <= 12'b111111111110;
   64893: result <= 12'b111111111110;
   64894: result <= 12'b111111111101;
   64895: result <= 12'b111111111101;
   64896: result <= 12'b111111111101;
   64897: result <= 12'b111111111101;
   64898: result <= 12'b111111111101;
   64899: result <= 12'b111111111100;
   64900: result <= 12'b111111111100;
   64901: result <= 12'b111111111100;
   64902: result <= 12'b111111111100;
   64903: result <= 12'b111111111100;
   64904: result <= 12'b111111111100;
   64905: result <= 12'b111111111011;
   64906: result <= 12'b111111111011;
   64907: result <= 12'b111111111011;
   64908: result <= 12'b111111111011;
   64909: result <= 12'b111111111011;
   64910: result <= 12'b111111111010;
   64911: result <= 12'b111111111010;
   64912: result <= 12'b111111111010;
   64913: result <= 12'b111111111010;
   64914: result <= 12'b111111111010;
   64915: result <= 12'b111111111001;
   64916: result <= 12'b111111111001;
   64917: result <= 12'b111111111001;
   64918: result <= 12'b111111111001;
   64919: result <= 12'b111111111001;
   64920: result <= 12'b111111111000;
   64921: result <= 12'b111111111000;
   64922: result <= 12'b111111111000;
   64923: result <= 12'b111111111000;
   64924: result <= 12'b111111111000;
   64925: result <= 12'b111111110111;
   64926: result <= 12'b111111110111;
   64927: result <= 12'b111111110111;
   64928: result <= 12'b111111110111;
   64929: result <= 12'b111111110111;
   64930: result <= 12'b111111110110;
   64931: result <= 12'b111111110110;
   64932: result <= 12'b111111110110;
   64933: result <= 12'b111111110110;
   64934: result <= 12'b111111110110;
   64935: result <= 12'b111111110101;
   64936: result <= 12'b111111110101;
   64937: result <= 12'b111111110101;
   64938: result <= 12'b111111110101;
   64939: result <= 12'b111111110101;
   64940: result <= 12'b111111110100;
   64941: result <= 12'b111111110100;
   64942: result <= 12'b111111110100;
   64943: result <= 12'b111111110100;
   64944: result <= 12'b111111110100;
   64945: result <= 12'b111111110011;
   64946: result <= 12'b111111110011;
   64947: result <= 12'b111111110011;
   64948: result <= 12'b111111110011;
   64949: result <= 12'b111111110011;
   64950: result <= 12'b111111110011;
   64951: result <= 12'b111111110010;
   64952: result <= 12'b111111110010;
   64953: result <= 12'b111111110010;
   64954: result <= 12'b111111110010;
   64955: result <= 12'b111111110010;
   64956: result <= 12'b111111110001;
   64957: result <= 12'b111111110001;
   64958: result <= 12'b111111110001;
   64959: result <= 12'b111111110001;
   64960: result <= 12'b111111110001;
   64961: result <= 12'b111111110000;
   64962: result <= 12'b111111110000;
   64963: result <= 12'b111111110000;
   64964: result <= 12'b111111110000;
   64965: result <= 12'b111111110000;
   64966: result <= 12'b111111101111;
   64967: result <= 12'b111111101111;
   64968: result <= 12'b111111101111;
   64969: result <= 12'b111111101111;
   64970: result <= 12'b111111101111;
   64971: result <= 12'b111111101110;
   64972: result <= 12'b111111101110;
   64973: result <= 12'b111111101110;
   64974: result <= 12'b111111101110;
   64975: result <= 12'b111111101110;
   64976: result <= 12'b111111101101;
   64977: result <= 12'b111111101101;
   64978: result <= 12'b111111101101;
   64979: result <= 12'b111111101101;
   64980: result <= 12'b111111101101;
   64981: result <= 12'b111111101100;
   64982: result <= 12'b111111101100;
   64983: result <= 12'b111111101100;
   64984: result <= 12'b111111101100;
   64985: result <= 12'b111111101100;
   64986: result <= 12'b111111101011;
   64987: result <= 12'b111111101011;
   64988: result <= 12'b111111101011;
   64989: result <= 12'b111111101011;
   64990: result <= 12'b111111101011;
   64991: result <= 12'b111111101010;
   64992: result <= 12'b111111101010;
   64993: result <= 12'b111111101010;
   64994: result <= 12'b111111101010;
   64995: result <= 12'b111111101010;
   64996: result <= 12'b111111101001;
   64997: result <= 12'b111111101001;
   64998: result <= 12'b111111101001;
   64999: result <= 12'b111111101001;
   65000: result <= 12'b111111101001;
   65001: result <= 12'b111111101001;
   65002: result <= 12'b111111101000;
   65003: result <= 12'b111111101000;
   65004: result <= 12'b111111101000;
   65005: result <= 12'b111111101000;
   65006: result <= 12'b111111101000;
   65007: result <= 12'b111111100111;
   65008: result <= 12'b111111100111;
   65009: result <= 12'b111111100111;
   65010: result <= 12'b111111100111;
   65011: result <= 12'b111111100111;
   65012: result <= 12'b111111100110;
   65013: result <= 12'b111111100110;
   65014: result <= 12'b111111100110;
   65015: result <= 12'b111111100110;
   65016: result <= 12'b111111100110;
   65017: result <= 12'b111111100101;
   65018: result <= 12'b111111100101;
   65019: result <= 12'b111111100101;
   65020: result <= 12'b111111100101;
   65021: result <= 12'b111111100101;
   65022: result <= 12'b111111100100;
   65023: result <= 12'b111111100100;
   65024: result <= 12'b111111100100;
   65025: result <= 12'b111111100100;
   65026: result <= 12'b111111100100;
   65027: result <= 12'b111111100011;
   65028: result <= 12'b111111100011;
   65029: result <= 12'b111111100011;
   65030: result <= 12'b111111100011;
   65031: result <= 12'b111111100011;
   65032: result <= 12'b111111100010;
   65033: result <= 12'b111111100010;
   65034: result <= 12'b111111100010;
   65035: result <= 12'b111111100010;
   65036: result <= 12'b111111100010;
   65037: result <= 12'b111111100001;
   65038: result <= 12'b111111100001;
   65039: result <= 12'b111111100001;
   65040: result <= 12'b111111100001;
   65041: result <= 12'b111111100001;
   65042: result <= 12'b111111100000;
   65043: result <= 12'b111111100000;
   65044: result <= 12'b111111100000;
   65045: result <= 12'b111111100000;
   65046: result <= 12'b111111100000;
   65047: result <= 12'b111111011111;
   65048: result <= 12'b111111011111;
   65049: result <= 12'b111111011111;
   65050: result <= 12'b111111011111;
   65051: result <= 12'b111111011111;
   65052: result <= 12'b111111011110;
   65053: result <= 12'b111111011110;
   65054: result <= 12'b111111011110;
   65055: result <= 12'b111111011110;
   65056: result <= 12'b111111011110;
   65057: result <= 12'b111111011110;
   65058: result <= 12'b111111011101;
   65059: result <= 12'b111111011101;
   65060: result <= 12'b111111011101;
   65061: result <= 12'b111111011101;
   65062: result <= 12'b111111011101;
   65063: result <= 12'b111111011100;
   65064: result <= 12'b111111011100;
   65065: result <= 12'b111111011100;
   65066: result <= 12'b111111011100;
   65067: result <= 12'b111111011100;
   65068: result <= 12'b111111011011;
   65069: result <= 12'b111111011011;
   65070: result <= 12'b111111011011;
   65071: result <= 12'b111111011011;
   65072: result <= 12'b111111011011;
   65073: result <= 12'b111111011010;
   65074: result <= 12'b111111011010;
   65075: result <= 12'b111111011010;
   65076: result <= 12'b111111011010;
   65077: result <= 12'b111111011010;
   65078: result <= 12'b111111011001;
   65079: result <= 12'b111111011001;
   65080: result <= 12'b111111011001;
   65081: result <= 12'b111111011001;
   65082: result <= 12'b111111011001;
   65083: result <= 12'b111111011000;
   65084: result <= 12'b111111011000;
   65085: result <= 12'b111111011000;
   65086: result <= 12'b111111011000;
   65087: result <= 12'b111111011000;
   65088: result <= 12'b111111010111;
   65089: result <= 12'b111111010111;
   65090: result <= 12'b111111010111;
   65091: result <= 12'b111111010111;
   65092: result <= 12'b111111010111;
   65093: result <= 12'b111111010110;
   65094: result <= 12'b111111010110;
   65095: result <= 12'b111111010110;
   65096: result <= 12'b111111010110;
   65097: result <= 12'b111111010110;
   65098: result <= 12'b111111010101;
   65099: result <= 12'b111111010101;
   65100: result <= 12'b111111010101;
   65101: result <= 12'b111111010101;
   65102: result <= 12'b111111010101;
   65103: result <= 12'b111111010100;
   65104: result <= 12'b111111010100;
   65105: result <= 12'b111111010100;
   65106: result <= 12'b111111010100;
   65107: result <= 12'b111111010100;
   65108: result <= 12'b111111010100;
   65109: result <= 12'b111111010011;
   65110: result <= 12'b111111010011;
   65111: result <= 12'b111111010011;
   65112: result <= 12'b111111010011;
   65113: result <= 12'b111111010011;
   65114: result <= 12'b111111010010;
   65115: result <= 12'b111111010010;
   65116: result <= 12'b111111010010;
   65117: result <= 12'b111111010010;
   65118: result <= 12'b111111010010;
   65119: result <= 12'b111111010001;
   65120: result <= 12'b111111010001;
   65121: result <= 12'b111111010001;
   65122: result <= 12'b111111010001;
   65123: result <= 12'b111111010001;
   65124: result <= 12'b111111010000;
   65125: result <= 12'b111111010000;
   65126: result <= 12'b111111010000;
   65127: result <= 12'b111111010000;
   65128: result <= 12'b111111010000;
   65129: result <= 12'b111111001111;
   65130: result <= 12'b111111001111;
   65131: result <= 12'b111111001111;
   65132: result <= 12'b111111001111;
   65133: result <= 12'b111111001111;
   65134: result <= 12'b111111001110;
   65135: result <= 12'b111111001110;
   65136: result <= 12'b111111001110;
   65137: result <= 12'b111111001110;
   65138: result <= 12'b111111001110;
   65139: result <= 12'b111111001101;
   65140: result <= 12'b111111001101;
   65141: result <= 12'b111111001101;
   65142: result <= 12'b111111001101;
   65143: result <= 12'b111111001101;
   65144: result <= 12'b111111001100;
   65145: result <= 12'b111111001100;
   65146: result <= 12'b111111001100;
   65147: result <= 12'b111111001100;
   65148: result <= 12'b111111001100;
   65149: result <= 12'b111111001011;
   65150: result <= 12'b111111001011;
   65151: result <= 12'b111111001011;
   65152: result <= 12'b111111001011;
   65153: result <= 12'b111111001011;
   65154: result <= 12'b111111001010;
   65155: result <= 12'b111111001010;
   65156: result <= 12'b111111001010;
   65157: result <= 12'b111111001010;
   65158: result <= 12'b111111001010;
   65159: result <= 12'b111111001010;
   65160: result <= 12'b111111001001;
   65161: result <= 12'b111111001001;
   65162: result <= 12'b111111001001;
   65163: result <= 12'b111111001001;
   65164: result <= 12'b111111001001;
   65165: result <= 12'b111111001000;
   65166: result <= 12'b111111001000;
   65167: result <= 12'b111111001000;
   65168: result <= 12'b111111001000;
   65169: result <= 12'b111111001000;
   65170: result <= 12'b111111000111;
   65171: result <= 12'b111111000111;
   65172: result <= 12'b111111000111;
   65173: result <= 12'b111111000111;
   65174: result <= 12'b111111000111;
   65175: result <= 12'b111111000110;
   65176: result <= 12'b111111000110;
   65177: result <= 12'b111111000110;
   65178: result <= 12'b111111000110;
   65179: result <= 12'b111111000110;
   65180: result <= 12'b111111000101;
   65181: result <= 12'b111111000101;
   65182: result <= 12'b111111000101;
   65183: result <= 12'b111111000101;
   65184: result <= 12'b111111000101;
   65185: result <= 12'b111111000100;
   65186: result <= 12'b111111000100;
   65187: result <= 12'b111111000100;
   65188: result <= 12'b111111000100;
   65189: result <= 12'b111111000100;
   65190: result <= 12'b111111000011;
   65191: result <= 12'b111111000011;
   65192: result <= 12'b111111000011;
   65193: result <= 12'b111111000011;
   65194: result <= 12'b111111000011;
   65195: result <= 12'b111111000010;
   65196: result <= 12'b111111000010;
   65197: result <= 12'b111111000010;
   65198: result <= 12'b111111000010;
   65199: result <= 12'b111111000010;
   65200: result <= 12'b111111000001;
   65201: result <= 12'b111111000001;
   65202: result <= 12'b111111000001;
   65203: result <= 12'b111111000001;
   65204: result <= 12'b111111000001;
   65205: result <= 12'b111111000000;
   65206: result <= 12'b111111000000;
   65207: result <= 12'b111111000000;
   65208: result <= 12'b111111000000;
   65209: result <= 12'b111111000000;
   65210: result <= 12'b111111111111;
   65211: result <= 12'b111111111111;
   65212: result <= 12'b111111111111;
   65213: result <= 12'b111111111111;
   65214: result <= 12'b111111111111;
   65215: result <= 12'b111111111111;
   65216: result <= 12'b111111111110;
   65217: result <= 12'b111111111110;
   65218: result <= 12'b111111111110;
   65219: result <= 12'b111111111110;
   65220: result <= 12'b111111111110;
   65221: result <= 12'b111111111101;
   65222: result <= 12'b111111111101;
   65223: result <= 12'b111111111101;
   65224: result <= 12'b111111111101;
   65225: result <= 12'b111111111101;
   65226: result <= 12'b111111111100;
   65227: result <= 12'b111111111100;
   65228: result <= 12'b111111111100;
   65229: result <= 12'b111111111100;
   65230: result <= 12'b111111111100;
   65231: result <= 12'b111111111011;
   65232: result <= 12'b111111111011;
   65233: result <= 12'b111111111011;
   65234: result <= 12'b111111111011;
   65235: result <= 12'b111111111011;
   65236: result <= 12'b111111111010;
   65237: result <= 12'b111111111010;
   65238: result <= 12'b111111111010;
   65239: result <= 12'b111111111010;
   65240: result <= 12'b111111111010;
   65241: result <= 12'b111111111001;
   65242: result <= 12'b111111111001;
   65243: result <= 12'b111111111001;
   65244: result <= 12'b111111111001;
   65245: result <= 12'b111111111001;
   65246: result <= 12'b111111111000;
   65247: result <= 12'b111111111000;
   65248: result <= 12'b111111111000;
   65249: result <= 12'b111111111000;
   65250: result <= 12'b111111111000;
   65251: result <= 12'b111111110111;
   65252: result <= 12'b111111110111;
   65253: result <= 12'b111111110111;
   65254: result <= 12'b111111110111;
   65255: result <= 12'b111111110111;
   65256: result <= 12'b111111110110;
   65257: result <= 12'b111111110110;
   65258: result <= 12'b111111110110;
   65259: result <= 12'b111111110110;
   65260: result <= 12'b111111110110;
   65261: result <= 12'b111111110101;
   65262: result <= 12'b111111110101;
   65263: result <= 12'b111111110101;
   65264: result <= 12'b111111110101;
   65265: result <= 12'b111111110101;
   65266: result <= 12'b111111110101;
   65267: result <= 12'b111111110100;
   65268: result <= 12'b111111110100;
   65269: result <= 12'b111111110100;
   65270: result <= 12'b111111110100;
   65271: result <= 12'b111111110100;
   65272: result <= 12'b111111110011;
   65273: result <= 12'b111111110011;
   65274: result <= 12'b111111110011;
   65275: result <= 12'b111111110011;
   65276: result <= 12'b111111110011;
   65277: result <= 12'b111111110010;
   65278: result <= 12'b111111110010;
   65279: result <= 12'b111111110010;
   65280: result <= 12'b111111110010;
   65281: result <= 12'b111111110010;
   65282: result <= 12'b111111110001;
   65283: result <= 12'b111111110001;
   65284: result <= 12'b111111110001;
   65285: result <= 12'b111111110001;
   65286: result <= 12'b111111110001;
   65287: result <= 12'b111111110000;
   65288: result <= 12'b111111110000;
   65289: result <= 12'b111111110000;
   65290: result <= 12'b111111110000;
   65291: result <= 12'b111111110000;
   65292: result <= 12'b111111101111;
   65293: result <= 12'b111111101111;
   65294: result <= 12'b111111101111;
   65295: result <= 12'b111111101111;
   65296: result <= 12'b111111101111;
   65297: result <= 12'b111111101110;
   65298: result <= 12'b111111101110;
   65299: result <= 12'b111111101110;
   65300: result <= 12'b111111101110;
   65301: result <= 12'b111111101110;
   65302: result <= 12'b111111101101;
   65303: result <= 12'b111111101101;
   65304: result <= 12'b111111101101;
   65305: result <= 12'b111111101101;
   65306: result <= 12'b111111101101;
   65307: result <= 12'b111111101100;
   65308: result <= 12'b111111101100;
   65309: result <= 12'b111111101100;
   65310: result <= 12'b111111101100;
   65311: result <= 12'b111111101100;
   65312: result <= 12'b111111101011;
   65313: result <= 12'b111111101011;
   65314: result <= 12'b111111101011;
   65315: result <= 12'b111111101011;
   65316: result <= 12'b111111101011;
   65317: result <= 12'b111111101010;
   65318: result <= 12'b111111101010;
   65319: result <= 12'b111111101010;
   65320: result <= 12'b111111101010;
   65321: result <= 12'b111111101010;
   65322: result <= 12'b111111101010;
   65323: result <= 12'b111111101001;
   65324: result <= 12'b111111101001;
   65325: result <= 12'b111111101001;
   65326: result <= 12'b111111101001;
   65327: result <= 12'b111111101001;
   65328: result <= 12'b111111101000;
   65329: result <= 12'b111111101000;
   65330: result <= 12'b111111101000;
   65331: result <= 12'b111111101000;
   65332: result <= 12'b111111101000;
   65333: result <= 12'b111111100111;
   65334: result <= 12'b111111100111;
   65335: result <= 12'b111111100111;
   65336: result <= 12'b111111100111;
   65337: result <= 12'b111111100111;
   65338: result <= 12'b111111100110;
   65339: result <= 12'b111111100110;
   65340: result <= 12'b111111100110;
   65341: result <= 12'b111111100110;
   65342: result <= 12'b111111100110;
   65343: result <= 12'b111111100101;
   65344: result <= 12'b111111100101;
   65345: result <= 12'b111111100101;
   65346: result <= 12'b111111100101;
   65347: result <= 12'b111111100101;
   65348: result <= 12'b111111100100;
   65349: result <= 12'b111111100100;
   65350: result <= 12'b111111100100;
   65351: result <= 12'b111111100100;
   65352: result <= 12'b111111100100;
   65353: result <= 12'b111111100011;
   65354: result <= 12'b111111100011;
   65355: result <= 12'b111111100011;
   65356: result <= 12'b111111100011;
   65357: result <= 12'b111111100011;
   65358: result <= 12'b111111100010;
   65359: result <= 12'b111111100010;
   65360: result <= 12'b111111100010;
   65361: result <= 12'b111111100010;
   65362: result <= 12'b111111100010;
   65363: result <= 12'b111111100001;
   65364: result <= 12'b111111100001;
   65365: result <= 12'b111111100001;
   65366: result <= 12'b111111100001;
   65367: result <= 12'b111111100001;
   65368: result <= 12'b111111100000;
   65369: result <= 12'b111111100000;
   65370: result <= 12'b111111100000;
   65371: result <= 12'b111111100000;
   65372: result <= 12'b111111100000;
   65373: result <= 12'b111111100000;
   65374: result <= 12'b111111111111;
   65375: result <= 12'b111111111111;
   65376: result <= 12'b111111111111;
   65377: result <= 12'b111111111111;
   65378: result <= 12'b111111111111;
   65379: result <= 12'b111111111110;
   65380: result <= 12'b111111111110;
   65381: result <= 12'b111111111110;
   65382: result <= 12'b111111111110;
   65383: result <= 12'b111111111110;
   65384: result <= 12'b111111111101;
   65385: result <= 12'b111111111101;
   65386: result <= 12'b111111111101;
   65387: result <= 12'b111111111101;
   65388: result <= 12'b111111111101;
   65389: result <= 12'b111111111100;
   65390: result <= 12'b111111111100;
   65391: result <= 12'b111111111100;
   65392: result <= 12'b111111111100;
   65393: result <= 12'b111111111100;
   65394: result <= 12'b111111111011;
   65395: result <= 12'b111111111011;
   65396: result <= 12'b111111111011;
   65397: result <= 12'b111111111011;
   65398: result <= 12'b111111111011;
   65399: result <= 12'b111111111010;
   65400: result <= 12'b111111111010;
   65401: result <= 12'b111111111010;
   65402: result <= 12'b111111111010;
   65403: result <= 12'b111111111010;
   65404: result <= 12'b111111111001;
   65405: result <= 12'b111111111001;
   65406: result <= 12'b111111111001;
   65407: result <= 12'b111111111001;
   65408: result <= 12'b111111111001;
   65409: result <= 12'b111111111000;
   65410: result <= 12'b111111111000;
   65411: result <= 12'b111111111000;
   65412: result <= 12'b111111111000;
   65413: result <= 12'b111111111000;
   65414: result <= 12'b111111110111;
   65415: result <= 12'b111111110111;
   65416: result <= 12'b111111110111;
   65417: result <= 12'b111111110111;
   65418: result <= 12'b111111110111;
   65419: result <= 12'b111111110110;
   65420: result <= 12'b111111110110;
   65421: result <= 12'b111111110110;
   65422: result <= 12'b111111110110;
   65423: result <= 12'b111111110110;
   65424: result <= 12'b111111110101;
   65425: result <= 12'b111111110101;
   65426: result <= 12'b111111110101;
   65427: result <= 12'b111111110101;
   65428: result <= 12'b111111110101;
   65429: result <= 12'b111111110101;
   65430: result <= 12'b111111110100;
   65431: result <= 12'b111111110100;
   65432: result <= 12'b111111110100;
   65433: result <= 12'b111111110100;
   65434: result <= 12'b111111110100;
   65435: result <= 12'b111111110011;
   65436: result <= 12'b111111110011;
   65437: result <= 12'b111111110011;
   65438: result <= 12'b111111110011;
   65439: result <= 12'b111111110011;
   65440: result <= 12'b111111110010;
   65441: result <= 12'b111111110010;
   65442: result <= 12'b111111110010;
   65443: result <= 12'b111111110010;
   65444: result <= 12'b111111110010;
   65445: result <= 12'b111111110001;
   65446: result <= 12'b111111110001;
   65447: result <= 12'b111111110001;
   65448: result <= 12'b111111110001;
   65449: result <= 12'b111111110001;
   65450: result <= 12'b111111110000;
   65451: result <= 12'b111111110000;
   65452: result <= 12'b111111110000;
   65453: result <= 12'b111111110000;
   65454: result <= 12'b111111110000;
   65455: result <= 12'b111111111111;
   65456: result <= 12'b111111111111;
   65457: result <= 12'b111111111111;
   65458: result <= 12'b111111111111;
   65459: result <= 12'b111111111111;
   65460: result <= 12'b111111111110;
   65461: result <= 12'b111111111110;
   65462: result <= 12'b111111111110;
   65463: result <= 12'b111111111110;
   65464: result <= 12'b111111111110;
   65465: result <= 12'b111111111101;
   65466: result <= 12'b111111111101;
   65467: result <= 12'b111111111101;
   65468: result <= 12'b111111111101;
   65469: result <= 12'b111111111101;
   65470: result <= 12'b111111111100;
   65471: result <= 12'b111111111100;
   65472: result <= 12'b111111111100;
   65473: result <= 12'b111111111100;
   65474: result <= 12'b111111111100;
   65475: result <= 12'b111111111011;
   65476: result <= 12'b111111111011;
   65477: result <= 12'b111111111011;
   65478: result <= 12'b111111111011;
   65479: result <= 12'b111111111011;
   65480: result <= 12'b111111111010;
   65481: result <= 12'b111111111010;
   65482: result <= 12'b111111111010;
   65483: result <= 12'b111111111010;
   65484: result <= 12'b111111111010;
   65485: result <= 12'b111111111010;
   65486: result <= 12'b111111111001;
   65487: result <= 12'b111111111001;
   65488: result <= 12'b111111111001;
   65489: result <= 12'b111111111001;
   65490: result <= 12'b111111111001;
   65491: result <= 12'b111111111000;
   65492: result <= 12'b111111111000;
   65493: result <= 12'b111111111000;
   65494: result <= 12'b111111111000;
   65495: result <= 12'b111111111000;
   65496: result <= 12'b111111111111;
   65497: result <= 12'b111111111111;
   65498: result <= 12'b111111111111;
   65499: result <= 12'b111111111111;
   65500: result <= 12'b111111111111;
   65501: result <= 12'b111111111110;
   65502: result <= 12'b111111111110;
   65503: result <= 12'b111111111110;
   65504: result <= 12'b111111111110;
   65505: result <= 12'b111111111110;
   65506: result <= 12'b111111111101;
   65507: result <= 12'b111111111101;
   65508: result <= 12'b111111111101;
   65509: result <= 12'b111111111101;
   65510: result <= 12'b111111111101;
   65511: result <= 12'b111111111100;
   65512: result <= 12'b111111111100;
   65513: result <= 12'b111111111100;
   65514: result <= 12'b111111111100;
   65515: result <= 12'b111111111100;
   65516: result <= 12'b111111111111;
   65517: result <= 12'b111111111111;
   65518: result <= 12'b111111111111;
   65519: result <= 12'b111111111111;
   65520: result <= 12'b111111111111;
   65521: result <= 12'b111111111110;
   65522: result <= 12'b111111111110;
   65523: result <= 12'b111111111110;
   65524: result <= 12'b111111111110;
   65525: result <= 12'b111111111110;
   65526: result <= 12'b111111111111;
   65527: result <= 12'b111111111111;
   65528: result <= 12'b111111111111;
   65529: result <= 12'b111111111111;
   65530: result <= 12'b111111111111;
   65531: result <= 12'b000000000000;
   65532: result <= 12'b000000000000;
   65533: result <= 12'b000000000000;
   65534: result <= 12'b000000000000;
   65535: result <= 12'b000000000000;
   endcase
endmodule
